magic
tech sky130A
magscale 1 2
timestamp 1712851378
<< metal3 >>
rect -1786 2512 1786 2540
rect -1786 -2512 1702 2512
rect 1766 -2512 1786 2512
rect -1786 -2540 1786 -2512
<< via3 >>
rect 1702 -2512 1766 2512
<< mimcap >>
rect -1746 2460 1454 2500
rect -1746 -2460 -1706 2460
rect 1414 -2460 1454 2460
rect -1746 -2500 1454 -2460
<< mimcapcontact >>
rect -1706 -2460 1414 2460
<< metal4 >>
rect 1686 2512 1782 2528
rect -1707 2460 1415 2461
rect -1707 -2460 -1706 2460
rect 1414 -2460 1415 2460
rect -1707 -2461 1415 -2460
rect 1686 -2512 1702 2512
rect 1766 -2512 1782 2512
rect 1686 -2528 1782 -2512
<< properties >>
string FIXED_BBOX -1786 -2540 1494 2540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 16 l 25 val 815.58 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
