magic
tech sky130A
magscale 1 2
timestamp 1712087189
<< nwell >>
rect -1312 -619 1312 619
<< pmos >>
rect -1116 -400 -716 400
rect -658 -400 -258 400
rect -200 -400 200 400
rect 258 -400 658 400
rect 716 -400 1116 400
<< pdiff >>
rect -1174 388 -1116 400
rect -1174 -388 -1162 388
rect -1128 -388 -1116 388
rect -1174 -400 -1116 -388
rect -716 388 -658 400
rect -716 -388 -704 388
rect -670 -388 -658 388
rect -716 -400 -658 -388
rect -258 388 -200 400
rect -258 -388 -246 388
rect -212 -388 -200 388
rect -258 -400 -200 -388
rect 200 388 258 400
rect 200 -388 212 388
rect 246 -388 258 388
rect 200 -400 258 -388
rect 658 388 716 400
rect 658 -388 670 388
rect 704 -388 716 388
rect 658 -400 716 -388
rect 1116 388 1174 400
rect 1116 -388 1128 388
rect 1162 -388 1174 388
rect 1116 -400 1174 -388
<< pdiffc >>
rect -1162 -388 -1128 388
rect -704 -388 -670 388
rect -246 -388 -212 388
rect 212 -388 246 388
rect 670 -388 704 388
rect 1128 -388 1162 388
<< nsubdiff >>
rect -1276 549 -1180 583
rect 1180 549 1276 583
rect -1276 487 -1242 549
rect 1242 487 1276 549
rect -1276 -549 -1242 -487
rect 1242 -549 1276 -487
rect -1276 -583 -1180 -549
rect 1180 -583 1276 -549
<< nsubdiffcont >>
rect -1180 549 1180 583
rect -1276 -487 -1242 487
rect 1242 -487 1276 487
rect -1180 -583 1180 -549
<< poly >>
rect -1116 481 -716 497
rect -1116 447 -1100 481
rect -732 447 -716 481
rect -1116 400 -716 447
rect -658 481 -258 497
rect -658 447 -642 481
rect -274 447 -258 481
rect -658 400 -258 447
rect -200 481 200 497
rect -200 447 -184 481
rect 184 447 200 481
rect -200 400 200 447
rect 258 481 658 497
rect 258 447 274 481
rect 642 447 658 481
rect 258 400 658 447
rect 716 481 1116 497
rect 716 447 732 481
rect 1100 447 1116 481
rect 716 400 1116 447
rect -1116 -447 -716 -400
rect -1116 -481 -1100 -447
rect -732 -481 -716 -447
rect -1116 -497 -716 -481
rect -658 -447 -258 -400
rect -658 -481 -642 -447
rect -274 -481 -258 -447
rect -658 -497 -258 -481
rect -200 -447 200 -400
rect -200 -481 -184 -447
rect 184 -481 200 -447
rect -200 -497 200 -481
rect 258 -447 658 -400
rect 258 -481 274 -447
rect 642 -481 658 -447
rect 258 -497 658 -481
rect 716 -447 1116 -400
rect 716 -481 732 -447
rect 1100 -481 1116 -447
rect 716 -497 1116 -481
<< polycont >>
rect -1100 447 -732 481
rect -642 447 -274 481
rect -184 447 184 481
rect 274 447 642 481
rect 732 447 1100 481
rect -1100 -481 -732 -447
rect -642 -481 -274 -447
rect -184 -481 184 -447
rect 274 -481 642 -447
rect 732 -481 1100 -447
<< locali >>
rect -1276 549 -1180 583
rect 1180 549 1276 583
rect -1276 487 -1242 549
rect 1242 487 1276 549
rect -1116 447 -1100 481
rect -732 447 -716 481
rect -658 447 -642 481
rect -274 447 -258 481
rect -200 447 -184 481
rect 184 447 200 481
rect 258 447 274 481
rect 642 447 658 481
rect 716 447 732 481
rect 1100 447 1116 481
rect -1162 388 -1128 404
rect -1162 -404 -1128 -388
rect -704 388 -670 404
rect -704 -404 -670 -388
rect -246 388 -212 404
rect -246 -404 -212 -388
rect 212 388 246 404
rect 212 -404 246 -388
rect 670 388 704 404
rect 670 -404 704 -388
rect 1128 388 1162 404
rect 1128 -404 1162 -388
rect -1116 -481 -1100 -447
rect -732 -481 -716 -447
rect -658 -481 -642 -447
rect -274 -481 -258 -447
rect -200 -481 -184 -447
rect 184 -481 200 -447
rect 258 -481 274 -447
rect 642 -481 658 -447
rect 716 -481 732 -447
rect 1100 -481 1116 -447
rect -1276 -549 -1242 -487
rect 1242 -549 1276 -487
rect -1276 -583 -1180 -549
rect 1180 -583 1276 -549
<< viali >>
rect -1100 447 -732 481
rect -642 447 -274 481
rect -184 447 184 481
rect 274 447 642 481
rect 732 447 1100 481
rect -1162 -388 -1128 388
rect -704 -388 -670 388
rect -246 -388 -212 388
rect 212 -388 246 388
rect 670 -388 704 388
rect 1128 -388 1162 388
rect -1100 -481 -732 -447
rect -642 -481 -274 -447
rect -184 -481 184 -447
rect 274 -481 642 -447
rect 732 -481 1100 -447
<< metal1 >>
rect -1112 481 -720 487
rect -1112 447 -1100 481
rect -732 447 -720 481
rect -1112 441 -720 447
rect -654 481 -262 487
rect -654 447 -642 481
rect -274 447 -262 481
rect -654 441 -262 447
rect -196 481 196 487
rect -196 447 -184 481
rect 184 447 196 481
rect -196 441 196 447
rect 262 481 654 487
rect 262 447 274 481
rect 642 447 654 481
rect 262 441 654 447
rect 720 481 1112 487
rect 720 447 732 481
rect 1100 447 1112 481
rect 720 441 1112 447
rect -1168 388 -1122 400
rect -1168 -388 -1162 388
rect -1128 -388 -1122 388
rect -1168 -400 -1122 -388
rect -710 388 -664 400
rect -710 -388 -704 388
rect -670 -388 -664 388
rect -710 -400 -664 -388
rect -252 388 -206 400
rect -252 -388 -246 388
rect -212 -388 -206 388
rect -252 -400 -206 -388
rect 206 388 252 400
rect 206 -388 212 388
rect 246 -388 252 388
rect 206 -400 252 -388
rect 664 388 710 400
rect 664 -388 670 388
rect 704 -388 710 388
rect 664 -400 710 -388
rect 1122 388 1168 400
rect 1122 -388 1128 388
rect 1162 -388 1168 388
rect 1122 -400 1168 -388
rect -1112 -447 -720 -441
rect -1112 -481 -1100 -447
rect -732 -481 -720 -447
rect -1112 -487 -720 -481
rect -654 -447 -262 -441
rect -654 -481 -642 -447
rect -274 -481 -262 -447
rect -654 -487 -262 -481
rect -196 -447 196 -441
rect -196 -481 -184 -447
rect 184 -481 196 -447
rect -196 -487 196 -481
rect 262 -447 654 -441
rect 262 -481 274 -447
rect 642 -481 654 -447
rect 262 -487 654 -481
rect 720 -447 1112 -441
rect 720 -481 732 -447
rect 1100 -481 1112 -447
rect 720 -487 1112 -481
<< properties >>
string FIXED_BBOX -1259 -566 1259 566
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.0 l 2.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
