magic
tech sky130A
timestamp 1712071977
<< pwell >>
rect -139 -1347 139 1347
<< mvnmos >>
rect -25 818 25 1218
rect -25 309 25 709
rect -25 -200 25 200
rect -25 -709 25 -309
rect -25 -1218 25 -818
<< mvndiff >>
rect -54 1212 -25 1218
rect -54 824 -48 1212
rect -31 824 -25 1212
rect -54 818 -25 824
rect 25 1212 54 1218
rect 25 824 31 1212
rect 48 824 54 1212
rect 25 818 54 824
rect -54 703 -25 709
rect -54 315 -48 703
rect -31 315 -25 703
rect -54 309 -25 315
rect 25 703 54 709
rect 25 315 31 703
rect 48 315 54 703
rect 25 309 54 315
rect -54 194 -25 200
rect -54 -194 -48 194
rect -31 -194 -25 194
rect -54 -200 -25 -194
rect 25 194 54 200
rect 25 -194 31 194
rect 48 -194 54 194
rect 25 -200 54 -194
rect -54 -315 -25 -309
rect -54 -703 -48 -315
rect -31 -703 -25 -315
rect -54 -709 -25 -703
rect 25 -315 54 -309
rect 25 -703 31 -315
rect 48 -703 54 -315
rect 25 -709 54 -703
rect -54 -824 -25 -818
rect -54 -1212 -48 -824
rect -31 -1212 -25 -824
rect -54 -1218 -25 -1212
rect 25 -824 54 -818
rect 25 -1212 31 -824
rect 48 -1212 54 -824
rect 25 -1218 54 -1212
<< mvndiffc >>
rect -48 824 -31 1212
rect 31 824 48 1212
rect -48 315 -31 703
rect 31 315 48 703
rect -48 -194 -31 194
rect 31 -194 48 194
rect -48 -703 -31 -315
rect 31 -703 48 -315
rect -48 -1212 -31 -824
rect 31 -1212 48 -824
<< mvpsubdiff >>
rect -121 1323 121 1329
rect -121 1306 -67 1323
rect 67 1306 121 1323
rect -121 1300 121 1306
rect -121 1275 -92 1300
rect -121 -1275 -115 1275
rect -98 -1275 -92 1275
rect 92 1275 121 1300
rect -121 -1300 -92 -1275
rect 92 -1275 98 1275
rect 115 -1275 121 1275
rect 92 -1300 121 -1275
rect -121 -1306 121 -1300
rect -121 -1323 -67 -1306
rect 67 -1323 121 -1306
rect -121 -1329 121 -1323
<< mvpsubdiffcont >>
rect -67 1306 67 1323
rect -115 -1275 -98 1275
rect 98 -1275 115 1275
rect -67 -1323 67 -1306
<< poly >>
rect -25 1254 25 1262
rect -25 1237 -17 1254
rect 17 1237 25 1254
rect -25 1218 25 1237
rect -25 799 25 818
rect -25 782 -17 799
rect 17 782 25 799
rect -25 774 25 782
rect -25 745 25 753
rect -25 728 -17 745
rect 17 728 25 745
rect -25 709 25 728
rect -25 290 25 309
rect -25 273 -17 290
rect 17 273 25 290
rect -25 265 25 273
rect -25 236 25 244
rect -25 219 -17 236
rect 17 219 25 236
rect -25 200 25 219
rect -25 -219 25 -200
rect -25 -236 -17 -219
rect 17 -236 25 -219
rect -25 -244 25 -236
rect -25 -273 25 -265
rect -25 -290 -17 -273
rect 17 -290 25 -273
rect -25 -309 25 -290
rect -25 -728 25 -709
rect -25 -745 -17 -728
rect 17 -745 25 -728
rect -25 -753 25 -745
rect -25 -782 25 -774
rect -25 -799 -17 -782
rect 17 -799 25 -782
rect -25 -818 25 -799
rect -25 -1237 25 -1218
rect -25 -1254 -17 -1237
rect 17 -1254 25 -1237
rect -25 -1262 25 -1254
<< polycont >>
rect -17 1237 17 1254
rect -17 782 17 799
rect -17 728 17 745
rect -17 273 17 290
rect -17 219 17 236
rect -17 -236 17 -219
rect -17 -290 17 -273
rect -17 -745 17 -728
rect -17 -799 17 -782
rect -17 -1254 17 -1237
<< locali >>
rect -115 1306 -67 1323
rect 67 1306 115 1323
rect -115 1275 -98 1306
rect 98 1275 115 1306
rect -25 1237 -17 1254
rect 17 1237 25 1254
rect -48 1212 -31 1220
rect -48 816 -31 824
rect 31 1212 48 1220
rect 31 816 48 824
rect -25 782 -17 799
rect 17 782 25 799
rect -25 728 -17 745
rect 17 728 25 745
rect -48 703 -31 711
rect -48 307 -31 315
rect 31 703 48 711
rect 31 307 48 315
rect -25 273 -17 290
rect 17 273 25 290
rect -25 219 -17 236
rect 17 219 25 236
rect -48 194 -31 202
rect -48 -202 -31 -194
rect 31 194 48 202
rect 31 -202 48 -194
rect -25 -236 -17 -219
rect 17 -236 25 -219
rect -25 -290 -17 -273
rect 17 -290 25 -273
rect -48 -315 -31 -307
rect -48 -711 -31 -703
rect 31 -315 48 -307
rect 31 -711 48 -703
rect -25 -745 -17 -728
rect 17 -745 25 -728
rect -25 -799 -17 -782
rect 17 -799 25 -782
rect -48 -824 -31 -816
rect -48 -1220 -31 -1212
rect 31 -824 48 -816
rect 31 -1220 48 -1212
rect -25 -1254 -17 -1237
rect 17 -1254 25 -1237
rect -115 -1306 -98 -1275
rect 98 -1306 115 -1275
rect -115 -1323 -67 -1306
rect 67 -1323 115 -1306
<< viali >>
rect -17 1237 17 1254
rect -48 824 -31 1212
rect 31 824 48 1212
rect -17 782 17 799
rect -17 728 17 745
rect -48 315 -31 703
rect 31 315 48 703
rect -17 273 17 290
rect -17 219 17 236
rect -48 -194 -31 194
rect 31 -194 48 194
rect -17 -236 17 -219
rect -17 -290 17 -273
rect -48 -703 -31 -315
rect 31 -703 48 -315
rect -17 -745 17 -728
rect -17 -799 17 -782
rect -48 -1212 -31 -824
rect 31 -1212 48 -824
rect -17 -1254 17 -1237
<< metal1 >>
rect -23 1254 23 1257
rect -23 1237 -17 1254
rect 17 1237 23 1254
rect -23 1234 23 1237
rect -51 1212 -28 1218
rect -51 824 -48 1212
rect -31 824 -28 1212
rect -51 818 -28 824
rect 28 1212 51 1218
rect 28 824 31 1212
rect 48 824 51 1212
rect 28 818 51 824
rect -23 799 23 802
rect -23 782 -17 799
rect 17 782 23 799
rect -23 779 23 782
rect -23 745 23 748
rect -23 728 -17 745
rect 17 728 23 745
rect -23 725 23 728
rect -51 703 -28 709
rect -51 315 -48 703
rect -31 315 -28 703
rect -51 309 -28 315
rect 28 703 51 709
rect 28 315 31 703
rect 48 315 51 703
rect 28 309 51 315
rect -23 290 23 293
rect -23 273 -17 290
rect 17 273 23 290
rect -23 270 23 273
rect -23 236 23 239
rect -23 219 -17 236
rect 17 219 23 236
rect -23 216 23 219
rect -51 194 -28 200
rect -51 -194 -48 194
rect -31 -194 -28 194
rect -51 -200 -28 -194
rect 28 194 51 200
rect 28 -194 31 194
rect 48 -194 51 194
rect 28 -200 51 -194
rect -23 -219 23 -216
rect -23 -236 -17 -219
rect 17 -236 23 -219
rect -23 -239 23 -236
rect -23 -273 23 -270
rect -23 -290 -17 -273
rect 17 -290 23 -273
rect -23 -293 23 -290
rect -51 -315 -28 -309
rect -51 -703 -48 -315
rect -31 -703 -28 -315
rect -51 -709 -28 -703
rect 28 -315 51 -309
rect 28 -703 31 -315
rect 48 -703 51 -315
rect 28 -709 51 -703
rect -23 -728 23 -725
rect -23 -745 -17 -728
rect 17 -745 23 -728
rect -23 -748 23 -745
rect -23 -782 23 -779
rect -23 -799 -17 -782
rect 17 -799 23 -782
rect -23 -802 23 -799
rect -51 -824 -28 -818
rect -51 -1212 -48 -824
rect -31 -1212 -28 -824
rect -51 -1218 -28 -1212
rect 28 -824 51 -818
rect 28 -1212 31 -824
rect 48 -1212 51 -824
rect 28 -1218 51 -1212
rect -23 -1237 23 -1234
rect -23 -1254 -17 -1237
rect 17 -1254 23 -1237
rect -23 -1257 23 -1254
<< properties >>
string FIXED_BBOX -106 -1314 106 1314
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 0.5 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
