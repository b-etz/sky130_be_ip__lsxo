magic
tech sky130A
magscale 1 2
timestamp 1712875330
<< error_s >>
rect 803 -1832 1124 -652
rect 1332 -1517 8216 -951
<< psubdiff >>
rect 1548 -682 1572 -622
rect 1632 -682 1656 -622
rect 4234 -682 4258 -622
rect 4318 -682 4342 -622
rect 7920 -682 7944 -622
rect 8004 -682 8028 -622
rect 472 -1694 532 -1670
rect 472 -1778 532 -1754
rect 1548 -1846 1572 -1786
rect 1632 -1846 1656 -1786
rect 4232 -1846 4256 -1786
rect 4316 -1846 4340 -1786
rect 7920 -1846 7944 -1786
rect 8004 -1846 8028 -1786
<< psubdiffcont >>
rect 1572 -682 1632 -622
rect 4258 -682 4318 -622
rect 7944 -682 8004 -622
rect 472 -1754 532 -1694
rect 1572 -1846 1632 -1786
rect 4256 -1846 4316 -1786
rect 7944 -1846 8004 -1786
<< locali >>
rect 216 -598 798 -584
rect 216 -770 230 -598
rect 402 -644 798 -598
rect 402 -770 416 -644
rect 216 -784 416 -770
rect 758 -776 798 -644
rect 1556 -682 1572 -622
rect 1632 -682 1648 -622
rect 4242 -682 4258 -622
rect 4318 -682 4334 -622
rect 7928 -682 7944 -622
rect 8004 -682 8020 -622
rect 742 -1412 886 -1390
rect 742 -1460 762 -1412
rect 862 -1460 886 -1412
rect 472 -1694 532 -1678
rect 472 -1770 532 -1754
rect 594 -1822 660 -1660
rect 594 -1842 694 -1822
rect 766 -1956 866 -1728
rect 968 -1822 1034 -1660
rect 968 -1842 1068 -1822
rect 1214 -1956 1314 -928
rect 1556 -1846 1572 -1786
rect 1632 -1846 1648 -1786
rect 4240 -1846 4256 -1786
rect 4316 -1846 4332 -1786
rect 7928 -1846 7944 -1786
rect 8004 -1846 8020 -1786
rect 490 -2056 1314 -1956
rect 490 -2068 690 -2056
rect 490 -2400 504 -2068
rect 676 -2400 690 -2068
rect 490 -2416 690 -2400
<< viali >>
rect 230 -770 402 -598
rect 758 -900 798 -812
rect 692 -1014 784 -980
rect 690 -1130 782 -1096
rect 758 -1268 798 -1190
rect 762 -1512 862 -1412
rect 594 -1922 694 -1842
rect 968 -1922 1068 -1842
rect 504 -2400 676 -2068
<< metal1 >>
rect 988 -304 1188 -290
rect 988 -478 1002 -304
rect 1174 -478 1188 -304
rect 988 -490 1188 -478
rect 216 -594 416 -584
rect 216 -774 226 -594
rect 406 -774 416 -594
rect 1038 -690 1134 -490
rect 8176 -742 8478 -642
rect 216 -784 416 -774
rect 742 -812 990 -798
rect 742 -904 756 -812
rect 976 -904 990 -812
rect 742 -918 990 -904
rect 678 -964 798 -958
rect 678 -1016 686 -964
rect 792 -1016 798 -964
rect 678 -1022 798 -1016
rect 678 -1090 798 -1084
rect 678 -1142 686 -1090
rect 792 -1142 798 -1090
rect 678 -1148 798 -1142
rect 740 -1190 988 -1184
rect 740 -1198 758 -1190
rect 798 -1198 988 -1190
rect 740 -1290 754 -1198
rect 974 -1290 988 -1198
rect 1086 -1282 1434 -1186
rect 740 -1304 988 -1290
rect 740 -1412 886 -1390
rect 740 -1512 762 -1412
rect 862 -1512 886 -1412
rect 740 -1556 886 -1512
rect 740 -1688 820 -1556
rect 740 -1756 746 -1688
rect 814 -1756 820 -1688
rect 8378 -1726 8478 -742
rect 740 -1762 820 -1756
rect 576 -1842 1086 -1826
rect 576 -1922 594 -1842
rect 694 -1922 968 -1842
rect 1068 -1922 1086 -1842
rect 576 -1938 1086 -1922
rect 490 -2068 690 -2056
rect 490 -2400 504 -2068
rect 676 -2400 690 -2068
rect 490 -2416 690 -2400
rect 886 -2106 1086 -1938
rect 1714 -1988 2504 -1976
rect 1714 -2066 1726 -1988
rect 2492 -2066 2504 -1988
rect 1714 -2074 2504 -2066
rect 2606 -2106 2706 -1792
rect 8176 -1826 8478 -1726
rect 886 -2206 1704 -2106
rect 2516 -2206 2706 -2106
rect 886 -2416 1086 -2206
<< via1 >>
rect 1002 -478 1174 -304
rect 226 -598 406 -594
rect 226 -770 230 -598
rect 230 -770 402 -598
rect 402 -770 406 -598
rect 226 -774 406 -770
rect 756 -900 758 -812
rect 758 -900 798 -812
rect 798 -900 976 -812
rect 756 -904 976 -900
rect 686 -980 792 -964
rect 686 -1014 692 -980
rect 692 -1014 784 -980
rect 784 -1014 792 -980
rect 686 -1016 792 -1014
rect 686 -1096 792 -1090
rect 686 -1130 690 -1096
rect 690 -1130 782 -1096
rect 782 -1130 792 -1096
rect 686 -1142 792 -1130
rect 754 -1268 758 -1198
rect 758 -1268 798 -1198
rect 798 -1268 974 -1198
rect 754 -1290 974 -1268
rect 746 -1756 814 -1688
rect 1726 -2066 2492 -1988
<< metal2 >>
rect 988 -304 1188 -290
rect 988 -478 1002 -304
rect 1174 -478 1188 -304
rect 988 -490 1188 -478
rect 1370 -542 8252 -442
rect 216 -594 416 -584
rect 216 -774 226 -594
rect 406 -774 416 -594
rect 216 -784 416 -774
rect 910 -642 1470 -542
rect 910 -798 990 -642
rect 742 -812 990 -798
rect 216 -950 416 -830
rect 742 -904 756 -812
rect 976 -904 990 -812
rect 742 -918 990 -904
rect 1256 -950 1336 -868
rect 8152 -930 8252 -542
rect 216 -964 1336 -950
rect 216 -1016 686 -964
rect 792 -1016 1336 -964
rect 216 -1030 1336 -1016
rect 216 -1090 1336 -1076
rect 216 -1142 686 -1090
rect 792 -1142 1336 -1090
rect 216 -1156 1336 -1142
rect 216 -1276 416 -1156
rect 740 -1198 988 -1184
rect 740 -1290 754 -1198
rect 974 -1290 988 -1198
rect 740 -1304 988 -1290
rect 740 -1688 820 -1682
rect 740 -1756 746 -1688
rect 814 -1756 820 -1688
rect 740 -1978 820 -1756
rect 908 -1826 988 -1304
rect 1256 -1608 1336 -1156
rect 908 -1926 2902 -1826
rect 8150 -1926 8250 -1538
rect 740 -1988 2504 -1978
rect 740 -2038 1726 -1988
rect 1714 -2066 1726 -2038
rect 2492 -2066 2504 -1988
rect 2802 -2026 8250 -1926
rect 1714 -2074 2504 -2066
use ripple_dly_4  x1
timestamp 1712867472
transform 1 0 1024 0 -1 -1868
box 232 -1226 7274 -586
use ripple_dly_4  x2
timestamp 1712867472
transform 1 0 1024 0 1 -600
box 232 -1226 7274 -586
use sky130_fd_sc_hd__a221o_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712867472
transform 0 1 542 -1 0 -690
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_0  x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712867472
transform 0 1 542 -1 0 -1426
box -38 -48 406 592
use sky130_fd_pr__nfet_01v8_AHZR5K  XM3
timestamp 1712867472
transform 1 0 2110 0 1 -2156
box -596 -260 596 260
<< labels >>
flabel space 1370 -673 8178 -642 0 FreeSans 800 0 0 0 dvss
flabel metal1 886 -2416 1086 -1922 0 FreeSans 800 0 0 0 clkout
port 4 nsew
flabel metal1 490 -2416 690 -2056 0 FreeSans 800 0 0 0 clkin
port 3 nsew
flabel metal2 216 -1030 416 -830 0 FreeSans 800 0 0 0 ena
port 5 nsew
flabel metal2 216 -1276 416 -1076 0 FreeSans 800 0 0 0 stby_b
port 8 nsew
flabel metal2 216 -784 416 -584 0 FreeSans 800 0 0 0 stby
port 6 nsew
flabel metal2 988 -490 1188 -290 0 FreeSans 800 0 0 0 dvdd
port 1 nsew
<< end >>
