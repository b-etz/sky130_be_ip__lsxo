magic
tech sky130A
magscale 1 2
timestamp 1712849042
<< metal3 >>
rect -4892 6932 -120 6960
rect -4892 2508 -204 6932
rect -140 2508 -120 6932
rect -4892 2480 -120 2508
rect 120 6932 4892 6960
rect 120 2508 4808 6932
rect 4872 2508 4892 6932
rect 120 2480 4892 2508
rect -4892 2212 -120 2240
rect -4892 -2212 -204 2212
rect -140 -2212 -120 2212
rect -4892 -2240 -120 -2212
rect 120 2212 4892 2240
rect 120 -2212 4808 2212
rect 4872 -2212 4892 2212
rect 120 -2240 4892 -2212
rect -4892 -2508 -120 -2480
rect -4892 -6932 -204 -2508
rect -140 -6932 -120 -2508
rect -4892 -6960 -120 -6932
rect 120 -2508 4892 -2480
rect 120 -6932 4808 -2508
rect 4872 -6932 4892 -2508
rect 120 -6960 4892 -6932
<< via3 >>
rect -204 2508 -140 6932
rect 4808 2508 4872 6932
rect -204 -2212 -140 2212
rect 4808 -2212 4872 2212
rect -204 -6932 -140 -2508
rect 4808 -6932 4872 -2508
<< mimcap >>
rect -4852 6880 -452 6920
rect -4852 2560 -4812 6880
rect -492 2560 -452 6880
rect -4852 2520 -452 2560
rect 160 6880 4560 6920
rect 160 2560 200 6880
rect 4520 2560 4560 6880
rect 160 2520 4560 2560
rect -4852 2160 -452 2200
rect -4852 -2160 -4812 2160
rect -492 -2160 -452 2160
rect -4852 -2200 -452 -2160
rect 160 2160 4560 2200
rect 160 -2160 200 2160
rect 4520 -2160 4560 2160
rect 160 -2200 4560 -2160
rect -4852 -2560 -452 -2520
rect -4852 -6880 -4812 -2560
rect -492 -6880 -452 -2560
rect -4852 -6920 -452 -6880
rect 160 -2560 4560 -2520
rect 160 -6880 200 -2560
rect 4520 -6880 4560 -2560
rect 160 -6920 4560 -6880
<< mimcapcontact >>
rect -4812 2560 -492 6880
rect 200 2560 4520 6880
rect -4812 -2160 -492 2160
rect 200 -2160 4520 2160
rect -4812 -6880 -492 -2560
rect 200 -6880 4520 -2560
<< metal4 >>
rect -2704 6881 -2600 7080
rect -224 6932 -120 7080
rect -4813 6880 -491 6881
rect -4813 2560 -4812 6880
rect -492 2560 -491 6880
rect -4813 2559 -491 2560
rect -2704 2161 -2600 2559
rect -224 2508 -204 6932
rect -140 2508 -120 6932
rect 2308 6881 2412 7080
rect 4788 6932 4892 7080
rect 199 6880 4521 6881
rect 199 2560 200 6880
rect 4520 2560 4521 6880
rect 199 2559 4521 2560
rect -224 2212 -120 2508
rect -4813 2160 -491 2161
rect -4813 -2160 -4812 2160
rect -492 -2160 -491 2160
rect -4813 -2161 -491 -2160
rect -2704 -2559 -2600 -2161
rect -224 -2212 -204 2212
rect -140 -2212 -120 2212
rect 2308 2161 2412 2559
rect 4788 2508 4808 6932
rect 4872 2508 4892 6932
rect 4788 2212 4892 2508
rect 199 2160 4521 2161
rect 199 -2160 200 2160
rect 4520 -2160 4521 2160
rect 199 -2161 4521 -2160
rect -224 -2508 -120 -2212
rect -4813 -2560 -491 -2559
rect -4813 -6880 -4812 -2560
rect -492 -6880 -491 -2560
rect -4813 -6881 -491 -6880
rect -2704 -7080 -2600 -6881
rect -224 -6932 -204 -2508
rect -140 -6932 -120 -2508
rect 2308 -2559 2412 -2161
rect 4788 -2212 4808 2212
rect 4872 -2212 4892 2212
rect 4788 -2508 4892 -2212
rect 199 -2560 4521 -2559
rect 199 -6880 200 -2560
rect 4520 -6880 4521 -2560
rect 199 -6881 4521 -6880
rect -224 -7080 -120 -6932
rect 2308 -7080 2412 -6881
rect 4788 -6932 4808 -2508
rect 4872 -6932 4892 -2508
rect 4788 -7080 4892 -6932
<< properties >>
string FIXED_BBOX 120 2480 4600 6960
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 22 l 22 val 984.72 carea 2.00 cperi 0.19 nx 2 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
