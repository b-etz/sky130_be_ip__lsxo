magic
tech sky130A
magscale 1 2
timestamp 1713142410
<< nwell >>
rect -2770 -1161 2770 1161
<< mvpmos >>
rect -2512 64 -2112 864
rect -1934 64 -1534 864
rect -1356 64 -956 864
rect -778 64 -378 864
rect -200 64 200 864
rect 378 64 778 864
rect 956 64 1356 864
rect 1534 64 1934 864
rect 2112 64 2512 864
rect -2512 -864 -2112 -64
rect -1934 -864 -1534 -64
rect -1356 -864 -956 -64
rect -778 -864 -378 -64
rect -200 -864 200 -64
rect 378 -864 778 -64
rect 956 -864 1356 -64
rect 1534 -864 1934 -64
rect 2112 -864 2512 -64
<< mvpdiff >>
rect -2570 852 -2512 864
rect -2570 76 -2558 852
rect -2524 76 -2512 852
rect -2570 64 -2512 76
rect -2112 852 -2054 864
rect -2112 76 -2100 852
rect -2066 76 -2054 852
rect -2112 64 -2054 76
rect -1992 852 -1934 864
rect -1992 76 -1980 852
rect -1946 76 -1934 852
rect -1992 64 -1934 76
rect -1534 852 -1476 864
rect -1534 76 -1522 852
rect -1488 76 -1476 852
rect -1534 64 -1476 76
rect -1414 852 -1356 864
rect -1414 76 -1402 852
rect -1368 76 -1356 852
rect -1414 64 -1356 76
rect -956 852 -898 864
rect -956 76 -944 852
rect -910 76 -898 852
rect -956 64 -898 76
rect -836 852 -778 864
rect -836 76 -824 852
rect -790 76 -778 852
rect -836 64 -778 76
rect -378 852 -320 864
rect -378 76 -366 852
rect -332 76 -320 852
rect -378 64 -320 76
rect -258 852 -200 864
rect -258 76 -246 852
rect -212 76 -200 852
rect -258 64 -200 76
rect 200 852 258 864
rect 200 76 212 852
rect 246 76 258 852
rect 200 64 258 76
rect 320 852 378 864
rect 320 76 332 852
rect 366 76 378 852
rect 320 64 378 76
rect 778 852 836 864
rect 778 76 790 852
rect 824 76 836 852
rect 778 64 836 76
rect 898 852 956 864
rect 898 76 910 852
rect 944 76 956 852
rect 898 64 956 76
rect 1356 852 1414 864
rect 1356 76 1368 852
rect 1402 76 1414 852
rect 1356 64 1414 76
rect 1476 852 1534 864
rect 1476 76 1488 852
rect 1522 76 1534 852
rect 1476 64 1534 76
rect 1934 852 1992 864
rect 1934 76 1946 852
rect 1980 76 1992 852
rect 1934 64 1992 76
rect 2054 852 2112 864
rect 2054 76 2066 852
rect 2100 76 2112 852
rect 2054 64 2112 76
rect 2512 852 2570 864
rect 2512 76 2524 852
rect 2558 76 2570 852
rect 2512 64 2570 76
rect -2570 -76 -2512 -64
rect -2570 -852 -2558 -76
rect -2524 -852 -2512 -76
rect -2570 -864 -2512 -852
rect -2112 -76 -2054 -64
rect -2112 -852 -2100 -76
rect -2066 -852 -2054 -76
rect -2112 -864 -2054 -852
rect -1992 -76 -1934 -64
rect -1992 -852 -1980 -76
rect -1946 -852 -1934 -76
rect -1992 -864 -1934 -852
rect -1534 -76 -1476 -64
rect -1534 -852 -1522 -76
rect -1488 -852 -1476 -76
rect -1534 -864 -1476 -852
rect -1414 -76 -1356 -64
rect -1414 -852 -1402 -76
rect -1368 -852 -1356 -76
rect -1414 -864 -1356 -852
rect -956 -76 -898 -64
rect -956 -852 -944 -76
rect -910 -852 -898 -76
rect -956 -864 -898 -852
rect -836 -76 -778 -64
rect -836 -852 -824 -76
rect -790 -852 -778 -76
rect -836 -864 -778 -852
rect -378 -76 -320 -64
rect -378 -852 -366 -76
rect -332 -852 -320 -76
rect -378 -864 -320 -852
rect -258 -76 -200 -64
rect -258 -852 -246 -76
rect -212 -852 -200 -76
rect -258 -864 -200 -852
rect 200 -76 258 -64
rect 200 -852 212 -76
rect 246 -852 258 -76
rect 200 -864 258 -852
rect 320 -76 378 -64
rect 320 -852 332 -76
rect 366 -852 378 -76
rect 320 -864 378 -852
rect 778 -76 836 -64
rect 778 -852 790 -76
rect 824 -852 836 -76
rect 778 -864 836 -852
rect 898 -76 956 -64
rect 898 -852 910 -76
rect 944 -852 956 -76
rect 898 -864 956 -852
rect 1356 -76 1414 -64
rect 1356 -852 1368 -76
rect 1402 -852 1414 -76
rect 1356 -864 1414 -852
rect 1476 -76 1534 -64
rect 1476 -852 1488 -76
rect 1522 -852 1534 -76
rect 1476 -864 1534 -852
rect 1934 -76 1992 -64
rect 1934 -852 1946 -76
rect 1980 -852 1992 -76
rect 1934 -864 1992 -852
rect 2054 -76 2112 -64
rect 2054 -852 2066 -76
rect 2100 -852 2112 -76
rect 2054 -864 2112 -852
rect 2512 -76 2570 -64
rect 2512 -852 2524 -76
rect 2558 -852 2570 -76
rect 2512 -864 2570 -852
<< mvpdiffc >>
rect -2558 76 -2524 852
rect -2100 76 -2066 852
rect -1980 76 -1946 852
rect -1522 76 -1488 852
rect -1402 76 -1368 852
rect -944 76 -910 852
rect -824 76 -790 852
rect -366 76 -332 852
rect -246 76 -212 852
rect 212 76 246 852
rect 332 76 366 852
rect 790 76 824 852
rect 910 76 944 852
rect 1368 76 1402 852
rect 1488 76 1522 852
rect 1946 76 1980 852
rect 2066 76 2100 852
rect 2524 76 2558 852
rect -2558 -852 -2524 -76
rect -2100 -852 -2066 -76
rect -1980 -852 -1946 -76
rect -1522 -852 -1488 -76
rect -1402 -852 -1368 -76
rect -944 -852 -910 -76
rect -824 -852 -790 -76
rect -366 -852 -332 -76
rect -246 -852 -212 -76
rect 212 -852 246 -76
rect 332 -852 366 -76
rect 790 -852 824 -76
rect 910 -852 944 -76
rect 1368 -852 1402 -76
rect 1488 -852 1522 -76
rect 1946 -852 1980 -76
rect 2066 -852 2100 -76
rect 2524 -852 2558 -76
<< mvnsubdiff >>
rect -2704 1083 2704 1095
rect -2704 1049 -2596 1083
rect 2596 1049 2704 1083
rect -2704 1037 2704 1049
rect -2704 987 -2646 1037
rect -2704 -987 -2692 987
rect -2658 -987 -2646 987
rect 2646 987 2704 1037
rect -2704 -1037 -2646 -987
rect 2646 -987 2658 987
rect 2692 -987 2704 987
rect 2646 -1037 2704 -987
rect -2704 -1049 2704 -1037
rect -2704 -1083 -2596 -1049
rect 2596 -1083 2704 -1049
rect -2704 -1095 2704 -1083
<< mvnsubdiffcont >>
rect -2596 1049 2596 1083
rect -2692 -987 -2658 987
rect 2658 -987 2692 987
rect -2596 -1083 2596 -1049
<< poly >>
rect -2512 945 -2112 961
rect -2512 911 -2496 945
rect -2128 911 -2112 945
rect -2512 864 -2112 911
rect -1934 945 -1534 961
rect -1934 911 -1918 945
rect -1550 911 -1534 945
rect -1934 864 -1534 911
rect -1356 945 -956 961
rect -1356 911 -1340 945
rect -972 911 -956 945
rect -1356 864 -956 911
rect -778 945 -378 961
rect -778 911 -762 945
rect -394 911 -378 945
rect -778 864 -378 911
rect -200 945 200 961
rect -200 911 -184 945
rect 184 911 200 945
rect -200 864 200 911
rect 378 945 778 961
rect 378 911 394 945
rect 762 911 778 945
rect 378 864 778 911
rect 956 945 1356 961
rect 956 911 972 945
rect 1340 911 1356 945
rect 956 864 1356 911
rect 1534 945 1934 961
rect 1534 911 1550 945
rect 1918 911 1934 945
rect 1534 864 1934 911
rect 2112 945 2512 961
rect 2112 911 2128 945
rect 2496 911 2512 945
rect 2112 864 2512 911
rect -2512 17 -2112 64
rect -2512 -17 -2496 17
rect -2128 -17 -2112 17
rect -2512 -64 -2112 -17
rect -1934 17 -1534 64
rect -1934 -17 -1918 17
rect -1550 -17 -1534 17
rect -1934 -64 -1534 -17
rect -1356 17 -956 64
rect -1356 -17 -1340 17
rect -972 -17 -956 17
rect -1356 -64 -956 -17
rect -778 17 -378 64
rect -778 -17 -762 17
rect -394 -17 -378 17
rect -778 -64 -378 -17
rect -200 17 200 64
rect -200 -17 -184 17
rect 184 -17 200 17
rect -200 -64 200 -17
rect 378 17 778 64
rect 378 -17 394 17
rect 762 -17 778 17
rect 378 -64 778 -17
rect 956 17 1356 64
rect 956 -17 972 17
rect 1340 -17 1356 17
rect 956 -64 1356 -17
rect 1534 17 1934 64
rect 1534 -17 1550 17
rect 1918 -17 1934 17
rect 1534 -64 1934 -17
rect 2112 17 2512 64
rect 2112 -17 2128 17
rect 2496 -17 2512 17
rect 2112 -64 2512 -17
rect -2512 -911 -2112 -864
rect -2512 -945 -2496 -911
rect -2128 -945 -2112 -911
rect -2512 -961 -2112 -945
rect -1934 -911 -1534 -864
rect -1934 -945 -1918 -911
rect -1550 -945 -1534 -911
rect -1934 -961 -1534 -945
rect -1356 -911 -956 -864
rect -1356 -945 -1340 -911
rect -972 -945 -956 -911
rect -1356 -961 -956 -945
rect -778 -911 -378 -864
rect -778 -945 -762 -911
rect -394 -945 -378 -911
rect -778 -961 -378 -945
rect -200 -911 200 -864
rect -200 -945 -184 -911
rect 184 -945 200 -911
rect -200 -961 200 -945
rect 378 -911 778 -864
rect 378 -945 394 -911
rect 762 -945 778 -911
rect 378 -961 778 -945
rect 956 -911 1356 -864
rect 956 -945 972 -911
rect 1340 -945 1356 -911
rect 956 -961 1356 -945
rect 1534 -911 1934 -864
rect 1534 -945 1550 -911
rect 1918 -945 1934 -911
rect 1534 -961 1934 -945
rect 2112 -911 2512 -864
rect 2112 -945 2128 -911
rect 2496 -945 2512 -911
rect 2112 -961 2512 -945
<< polycont >>
rect -2496 911 -2128 945
rect -1918 911 -1550 945
rect -1340 911 -972 945
rect -762 911 -394 945
rect -184 911 184 945
rect 394 911 762 945
rect 972 911 1340 945
rect 1550 911 1918 945
rect 2128 911 2496 945
rect -2496 -17 -2128 17
rect -1918 -17 -1550 17
rect -1340 -17 -972 17
rect -762 -17 -394 17
rect -184 -17 184 17
rect 394 -17 762 17
rect 972 -17 1340 17
rect 1550 -17 1918 17
rect 2128 -17 2496 17
rect -2496 -945 -2128 -911
rect -1918 -945 -1550 -911
rect -1340 -945 -972 -911
rect -762 -945 -394 -911
rect -184 -945 184 -911
rect 394 -945 762 -911
rect 972 -945 1340 -911
rect 1550 -945 1918 -911
rect 2128 -945 2496 -911
<< locali >>
rect -2692 1049 -2596 1083
rect 2596 1049 2692 1083
rect -2692 987 -2658 1049
rect 2658 987 2692 1049
rect -2512 911 -2496 945
rect -2128 911 -2112 945
rect -1934 911 -1918 945
rect -1550 911 -1534 945
rect -1356 911 -1340 945
rect -972 911 -956 945
rect -778 911 -762 945
rect -394 911 -378 945
rect -200 911 -184 945
rect 184 911 200 945
rect 378 911 394 945
rect 762 911 778 945
rect 956 911 972 945
rect 1340 911 1356 945
rect 1534 911 1550 945
rect 1918 911 1934 945
rect 2112 911 2128 945
rect 2496 911 2512 945
rect -2558 852 -2524 868
rect -2558 60 -2524 76
rect -2100 852 -2066 868
rect -2100 60 -2066 76
rect -1980 852 -1946 868
rect -1980 60 -1946 76
rect -1522 852 -1488 868
rect -1522 60 -1488 76
rect -1402 852 -1368 868
rect -1402 60 -1368 76
rect -944 852 -910 868
rect -944 60 -910 76
rect -824 852 -790 868
rect -824 60 -790 76
rect -366 852 -332 868
rect -366 60 -332 76
rect -246 852 -212 868
rect -246 60 -212 76
rect 212 852 246 868
rect 212 60 246 76
rect 332 852 366 868
rect 332 60 366 76
rect 790 852 824 868
rect 790 60 824 76
rect 910 852 944 868
rect 910 60 944 76
rect 1368 852 1402 868
rect 1368 60 1402 76
rect 1488 852 1522 868
rect 1488 60 1522 76
rect 1946 852 1980 868
rect 1946 60 1980 76
rect 2066 852 2100 868
rect 2066 60 2100 76
rect 2524 852 2558 868
rect 2524 60 2558 76
rect -2512 -17 -2496 17
rect -2128 -17 -2112 17
rect -1934 -17 -1918 17
rect -1550 -17 -1534 17
rect -1356 -17 -1340 17
rect -972 -17 -956 17
rect -778 -17 -762 17
rect -394 -17 -378 17
rect -200 -17 -184 17
rect 184 -17 200 17
rect 378 -17 394 17
rect 762 -17 778 17
rect 956 -17 972 17
rect 1340 -17 1356 17
rect 1534 -17 1550 17
rect 1918 -17 1934 17
rect 2112 -17 2128 17
rect 2496 -17 2512 17
rect -2558 -76 -2524 -60
rect -2558 -868 -2524 -852
rect -2100 -76 -2066 -60
rect -2100 -868 -2066 -852
rect -1980 -76 -1946 -60
rect -1980 -868 -1946 -852
rect -1522 -76 -1488 -60
rect -1522 -868 -1488 -852
rect -1402 -76 -1368 -60
rect -1402 -868 -1368 -852
rect -944 -76 -910 -60
rect -944 -868 -910 -852
rect -824 -76 -790 -60
rect -824 -868 -790 -852
rect -366 -76 -332 -60
rect -366 -868 -332 -852
rect -246 -76 -212 -60
rect -246 -868 -212 -852
rect 212 -76 246 -60
rect 212 -868 246 -852
rect 332 -76 366 -60
rect 332 -868 366 -852
rect 790 -76 824 -60
rect 790 -868 824 -852
rect 910 -76 944 -60
rect 910 -868 944 -852
rect 1368 -76 1402 -60
rect 1368 -868 1402 -852
rect 1488 -76 1522 -60
rect 1488 -868 1522 -852
rect 1946 -76 1980 -60
rect 1946 -868 1980 -852
rect 2066 -76 2100 -60
rect 2066 -868 2100 -852
rect 2524 -76 2558 -60
rect 2524 -868 2558 -852
rect -2512 -945 -2496 -911
rect -2128 -945 -2112 -911
rect -1934 -945 -1918 -911
rect -1550 -945 -1534 -911
rect -1356 -945 -1340 -911
rect -972 -945 -956 -911
rect -778 -945 -762 -911
rect -394 -945 -378 -911
rect -200 -945 -184 -911
rect 184 -945 200 -911
rect 378 -945 394 -911
rect 762 -945 778 -911
rect 956 -945 972 -911
rect 1340 -945 1356 -911
rect 1534 -945 1550 -911
rect 1918 -945 1934 -911
rect 2112 -945 2128 -911
rect 2496 -945 2512 -911
rect -2692 -1049 -2658 -987
rect 2658 -1049 2692 -987
rect -2692 -1083 -2596 -1049
rect 2596 -1083 2692 -1049
<< viali >>
rect -2459 911 -2165 945
rect -1881 911 -1587 945
rect -1303 911 -1009 945
rect -725 911 -431 945
rect -147 911 147 945
rect 431 911 725 945
rect 1009 911 1303 945
rect 1587 911 1881 945
rect 2165 911 2459 945
rect -2558 76 -2524 852
rect -2100 76 -2066 852
rect -1980 76 -1946 852
rect -1522 76 -1488 852
rect -1402 76 -1368 852
rect -944 76 -910 852
rect -824 76 -790 852
rect -366 76 -332 852
rect -246 76 -212 852
rect 212 76 246 852
rect 332 76 366 852
rect 790 76 824 852
rect 910 76 944 852
rect 1368 76 1402 852
rect 1488 76 1522 852
rect 1946 76 1980 852
rect 2066 76 2100 852
rect 2524 76 2558 852
rect -2459 -17 -2165 17
rect -1881 -17 -1587 17
rect -1303 -17 -1009 17
rect -725 -17 -431 17
rect -147 -17 147 17
rect 431 -17 725 17
rect 1009 -17 1303 17
rect 1587 -17 1881 17
rect 2165 -17 2459 17
rect -2558 -852 -2524 -76
rect -2100 -852 -2066 -76
rect -1980 -852 -1946 -76
rect -1522 -852 -1488 -76
rect -1402 -852 -1368 -76
rect -944 -852 -910 -76
rect -824 -852 -790 -76
rect -366 -852 -332 -76
rect -246 -852 -212 -76
rect 212 -852 246 -76
rect 332 -852 366 -76
rect 790 -852 824 -76
rect 910 -852 944 -76
rect 1368 -852 1402 -76
rect 1488 -852 1522 -76
rect 1946 -852 1980 -76
rect 2066 -852 2100 -76
rect 2524 -852 2558 -76
rect -2459 -945 -2165 -911
rect -1881 -945 -1587 -911
rect -1303 -945 -1009 -911
rect -725 -945 -431 -911
rect -147 -945 147 -911
rect 431 -945 725 -911
rect 1009 -945 1303 -911
rect 1587 -945 1881 -911
rect 2165 -945 2459 -911
<< metal1 >>
rect -2471 945 -2153 951
rect -2471 911 -2459 945
rect -2165 911 -2153 945
rect -2471 905 -2153 911
rect -1893 945 -1575 951
rect -1893 911 -1881 945
rect -1587 911 -1575 945
rect -1893 905 -1575 911
rect -1315 945 -997 951
rect -1315 911 -1303 945
rect -1009 911 -997 945
rect -1315 905 -997 911
rect -737 945 -419 951
rect -737 911 -725 945
rect -431 911 -419 945
rect -737 905 -419 911
rect -159 945 159 951
rect -159 911 -147 945
rect 147 911 159 945
rect -159 905 159 911
rect 419 945 737 951
rect 419 911 431 945
rect 725 911 737 945
rect 419 905 737 911
rect 997 945 1315 951
rect 997 911 1009 945
rect 1303 911 1315 945
rect 997 905 1315 911
rect 1575 945 1893 951
rect 1575 911 1587 945
rect 1881 911 1893 945
rect 1575 905 1893 911
rect 2153 945 2471 951
rect 2153 911 2165 945
rect 2459 911 2471 945
rect 2153 905 2471 911
rect -2564 852 -2518 864
rect -2564 76 -2558 852
rect -2524 76 -2518 852
rect -2564 64 -2518 76
rect -2106 852 -2060 864
rect -2106 76 -2100 852
rect -2066 76 -2060 852
rect -2106 64 -2060 76
rect -1986 852 -1940 864
rect -1986 76 -1980 852
rect -1946 76 -1940 852
rect -1986 64 -1940 76
rect -1528 852 -1482 864
rect -1528 76 -1522 852
rect -1488 76 -1482 852
rect -1528 64 -1482 76
rect -1408 852 -1362 864
rect -1408 76 -1402 852
rect -1368 76 -1362 852
rect -1408 64 -1362 76
rect -950 852 -904 864
rect -950 76 -944 852
rect -910 76 -904 852
rect -950 64 -904 76
rect -830 852 -784 864
rect -830 76 -824 852
rect -790 76 -784 852
rect -830 64 -784 76
rect -372 852 -326 864
rect -372 76 -366 852
rect -332 76 -326 852
rect -372 64 -326 76
rect -252 852 -206 864
rect -252 76 -246 852
rect -212 76 -206 852
rect -252 64 -206 76
rect 206 852 252 864
rect 206 76 212 852
rect 246 76 252 852
rect 206 64 252 76
rect 326 852 372 864
rect 326 76 332 852
rect 366 76 372 852
rect 326 64 372 76
rect 784 852 830 864
rect 784 76 790 852
rect 824 76 830 852
rect 784 64 830 76
rect 904 852 950 864
rect 904 76 910 852
rect 944 76 950 852
rect 904 64 950 76
rect 1362 852 1408 864
rect 1362 76 1368 852
rect 1402 76 1408 852
rect 1362 64 1408 76
rect 1482 852 1528 864
rect 1482 76 1488 852
rect 1522 76 1528 852
rect 1482 64 1528 76
rect 1940 852 1986 864
rect 1940 76 1946 852
rect 1980 76 1986 852
rect 1940 64 1986 76
rect 2060 852 2106 864
rect 2060 76 2066 852
rect 2100 76 2106 852
rect 2060 64 2106 76
rect 2518 852 2564 864
rect 2518 76 2524 852
rect 2558 76 2564 852
rect 2518 64 2564 76
rect -2471 17 -2153 23
rect -2471 -17 -2459 17
rect -2165 -17 -2153 17
rect -2471 -23 -2153 -17
rect -1893 17 -1575 23
rect -1893 -17 -1881 17
rect -1587 -17 -1575 17
rect -1893 -23 -1575 -17
rect -1315 17 -997 23
rect -1315 -17 -1303 17
rect -1009 -17 -997 17
rect -1315 -23 -997 -17
rect -737 17 -419 23
rect -737 -17 -725 17
rect -431 -17 -419 17
rect -737 -23 -419 -17
rect -159 17 159 23
rect -159 -17 -147 17
rect 147 -17 159 17
rect -159 -23 159 -17
rect 419 17 737 23
rect 419 -17 431 17
rect 725 -17 737 17
rect 419 -23 737 -17
rect 997 17 1315 23
rect 997 -17 1009 17
rect 1303 -17 1315 17
rect 997 -23 1315 -17
rect 1575 17 1893 23
rect 1575 -17 1587 17
rect 1881 -17 1893 17
rect 1575 -23 1893 -17
rect 2153 17 2471 23
rect 2153 -17 2165 17
rect 2459 -17 2471 17
rect 2153 -23 2471 -17
rect -2564 -76 -2518 -64
rect -2564 -852 -2558 -76
rect -2524 -852 -2518 -76
rect -2564 -864 -2518 -852
rect -2106 -76 -2060 -64
rect -2106 -852 -2100 -76
rect -2066 -852 -2060 -76
rect -2106 -864 -2060 -852
rect -1986 -76 -1940 -64
rect -1986 -852 -1980 -76
rect -1946 -852 -1940 -76
rect -1986 -864 -1940 -852
rect -1528 -76 -1482 -64
rect -1528 -852 -1522 -76
rect -1488 -852 -1482 -76
rect -1528 -864 -1482 -852
rect -1408 -76 -1362 -64
rect -1408 -852 -1402 -76
rect -1368 -852 -1362 -76
rect -1408 -864 -1362 -852
rect -950 -76 -904 -64
rect -950 -852 -944 -76
rect -910 -852 -904 -76
rect -950 -864 -904 -852
rect -830 -76 -784 -64
rect -830 -852 -824 -76
rect -790 -852 -784 -76
rect -830 -864 -784 -852
rect -372 -76 -326 -64
rect -372 -852 -366 -76
rect -332 -852 -326 -76
rect -372 -864 -326 -852
rect -252 -76 -206 -64
rect -252 -852 -246 -76
rect -212 -852 -206 -76
rect -252 -864 -206 -852
rect 206 -76 252 -64
rect 206 -852 212 -76
rect 246 -852 252 -76
rect 206 -864 252 -852
rect 326 -76 372 -64
rect 326 -852 332 -76
rect 366 -852 372 -76
rect 326 -864 372 -852
rect 784 -76 830 -64
rect 784 -852 790 -76
rect 824 -852 830 -76
rect 784 -864 830 -852
rect 904 -76 950 -64
rect 904 -852 910 -76
rect 944 -852 950 -76
rect 904 -864 950 -852
rect 1362 -76 1408 -64
rect 1362 -852 1368 -76
rect 1402 -852 1408 -76
rect 1362 -864 1408 -852
rect 1482 -76 1528 -64
rect 1482 -852 1488 -76
rect 1522 -852 1528 -76
rect 1482 -864 1528 -852
rect 1940 -76 1986 -64
rect 1940 -852 1946 -76
rect 1980 -852 1986 -76
rect 1940 -864 1986 -852
rect 2060 -76 2106 -64
rect 2060 -852 2066 -76
rect 2100 -852 2106 -76
rect 2060 -864 2106 -852
rect 2518 -76 2564 -64
rect 2518 -852 2524 -76
rect 2558 -852 2564 -76
rect 2518 -864 2564 -852
rect -2471 -911 -2153 -905
rect -2471 -945 -2459 -911
rect -2165 -945 -2153 -911
rect -2471 -951 -2153 -945
rect -1893 -911 -1575 -905
rect -1893 -945 -1881 -911
rect -1587 -945 -1575 -911
rect -1893 -951 -1575 -945
rect -1315 -911 -997 -905
rect -1315 -945 -1303 -911
rect -1009 -945 -997 -911
rect -1315 -951 -997 -945
rect -737 -911 -419 -905
rect -737 -945 -725 -911
rect -431 -945 -419 -911
rect -737 -951 -419 -945
rect -159 -911 159 -905
rect -159 -945 -147 -911
rect 147 -945 159 -911
rect -159 -951 159 -945
rect 419 -911 737 -905
rect 419 -945 431 -911
rect 725 -945 737 -911
rect 419 -951 737 -945
rect 997 -911 1315 -905
rect 997 -945 1009 -911
rect 1303 -945 1315 -911
rect 997 -951 1315 -945
rect 1575 -911 1893 -905
rect 1575 -945 1587 -911
rect 1881 -945 1893 -911
rect 1575 -951 1893 -945
rect 2153 -911 2471 -905
rect 2153 -945 2165 -911
rect 2459 -945 2471 -911
rect 2153 -951 2471 -945
<< properties >>
string FIXED_BBOX -2675 -1066 2675 1066
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 2.0 m 2 nf 9 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
