magic
tech sky130A
timestamp 1712848480
<< pwell >>
rect -901 -329 901 329
<< mvnmos >>
rect -787 -200 -587 200
rect -558 -200 -358 200
rect -329 -200 -129 200
rect -100 -200 100 200
rect 129 -200 329 200
rect 358 -200 558 200
rect 587 -200 787 200
<< mvndiff >>
rect -816 194 -787 200
rect -816 -194 -810 194
rect -793 -194 -787 194
rect -816 -200 -787 -194
rect -587 194 -558 200
rect -587 -194 -581 194
rect -564 -194 -558 194
rect -587 -200 -558 -194
rect -358 194 -329 200
rect -358 -194 -352 194
rect -335 -194 -329 194
rect -358 -200 -329 -194
rect -129 194 -100 200
rect -129 -194 -123 194
rect -106 -194 -100 194
rect -129 -200 -100 -194
rect 100 194 129 200
rect 100 -194 106 194
rect 123 -194 129 194
rect 100 -200 129 -194
rect 329 194 358 200
rect 329 -194 335 194
rect 352 -194 358 194
rect 329 -200 358 -194
rect 558 194 587 200
rect 558 -194 564 194
rect 581 -194 587 194
rect 558 -200 587 -194
rect 787 194 816 200
rect 787 -194 793 194
rect 810 -194 816 194
rect 787 -200 816 -194
<< mvndiffc >>
rect -810 -194 -793 194
rect -581 -194 -564 194
rect -352 -194 -335 194
rect -123 -194 -106 194
rect 106 -194 123 194
rect 335 -194 352 194
rect 564 -194 581 194
rect 793 -194 810 194
<< mvpsubdiff >>
rect -883 305 883 311
rect -883 288 -829 305
rect 829 288 883 305
rect -883 282 883 288
rect -883 257 -854 282
rect -883 -257 -877 257
rect -860 -257 -854 257
rect 854 257 883 282
rect -883 -282 -854 -257
rect 854 -257 860 257
rect 877 -257 883 257
rect 854 -282 883 -257
rect -883 -288 883 -282
rect -883 -305 -829 -288
rect 829 -305 883 -288
rect -883 -311 883 -305
<< mvpsubdiffcont >>
rect -829 288 829 305
rect -877 -257 -860 257
rect 860 -257 877 257
rect -829 -305 829 -288
<< poly >>
rect -787 236 -587 244
rect -787 219 -779 236
rect -595 219 -587 236
rect -787 200 -587 219
rect -558 236 -358 244
rect -558 219 -550 236
rect -366 219 -358 236
rect -558 200 -358 219
rect -329 236 -129 244
rect -329 219 -321 236
rect -137 219 -129 236
rect -329 200 -129 219
rect -100 236 100 244
rect -100 219 -92 236
rect 92 219 100 236
rect -100 200 100 219
rect 129 236 329 244
rect 129 219 137 236
rect 321 219 329 236
rect 129 200 329 219
rect 358 236 558 244
rect 358 219 366 236
rect 550 219 558 236
rect 358 200 558 219
rect 587 236 787 244
rect 587 219 595 236
rect 779 219 787 236
rect 587 200 787 219
rect -787 -219 -587 -200
rect -787 -236 -779 -219
rect -595 -236 -587 -219
rect -787 -244 -587 -236
rect -558 -219 -358 -200
rect -558 -236 -550 -219
rect -366 -236 -358 -219
rect -558 -244 -358 -236
rect -329 -219 -129 -200
rect -329 -236 -321 -219
rect -137 -236 -129 -219
rect -329 -244 -129 -236
rect -100 -219 100 -200
rect -100 -236 -92 -219
rect 92 -236 100 -219
rect -100 -244 100 -236
rect 129 -219 329 -200
rect 129 -236 137 -219
rect 321 -236 329 -219
rect 129 -244 329 -236
rect 358 -219 558 -200
rect 358 -236 366 -219
rect 550 -236 558 -219
rect 358 -244 558 -236
rect 587 -219 787 -200
rect 587 -236 595 -219
rect 779 -236 787 -219
rect 587 -244 787 -236
<< polycont >>
rect -779 219 -595 236
rect -550 219 -366 236
rect -321 219 -137 236
rect -92 219 92 236
rect 137 219 321 236
rect 366 219 550 236
rect 595 219 779 236
rect -779 -236 -595 -219
rect -550 -236 -366 -219
rect -321 -236 -137 -219
rect -92 -236 92 -219
rect 137 -236 321 -219
rect 366 -236 550 -219
rect 595 -236 779 -219
<< locali >>
rect -877 288 -829 305
rect 829 288 877 305
rect -877 257 -860 288
rect 860 257 877 288
rect -787 219 -779 236
rect -595 219 -587 236
rect -558 219 -550 236
rect -366 219 -358 236
rect -329 219 -321 236
rect -137 219 -129 236
rect -100 219 -92 236
rect 92 219 100 236
rect 129 219 137 236
rect 321 219 329 236
rect 358 219 366 236
rect 550 219 558 236
rect 587 219 595 236
rect 779 219 787 236
rect -810 194 -793 202
rect -810 -202 -793 -194
rect -581 194 -564 202
rect -581 -202 -564 -194
rect -352 194 -335 202
rect -352 -202 -335 -194
rect -123 194 -106 202
rect -123 -202 -106 -194
rect 106 194 123 202
rect 106 -202 123 -194
rect 335 194 352 202
rect 335 -202 352 -194
rect 564 194 581 202
rect 564 -202 581 -194
rect 793 194 810 202
rect 793 -202 810 -194
rect -787 -236 -779 -219
rect -595 -236 -587 -219
rect -558 -236 -550 -219
rect -366 -236 -358 -219
rect -329 -236 -321 -219
rect -137 -236 -129 -219
rect -100 -236 -92 -219
rect 92 -236 100 -219
rect 129 -236 137 -219
rect 321 -236 329 -219
rect 358 -236 366 -219
rect 550 -236 558 -219
rect 587 -236 595 -219
rect 779 -236 787 -219
rect -877 -288 -860 -257
rect 860 -288 877 -257
rect -877 -305 -829 -288
rect 829 -305 877 -288
<< viali >>
rect -779 219 -595 236
rect -550 219 -366 236
rect -321 219 -137 236
rect -92 219 92 236
rect 137 219 321 236
rect 366 219 550 236
rect 595 219 779 236
rect -810 -194 -793 194
rect -581 -194 -564 194
rect -352 -194 -335 194
rect -123 -194 -106 194
rect 106 -194 123 194
rect 335 -194 352 194
rect 564 -194 581 194
rect 793 -194 810 194
rect -779 -236 -595 -219
rect -550 -236 -366 -219
rect -321 -236 -137 -219
rect -92 -236 92 -219
rect 137 -236 321 -219
rect 366 -236 550 -219
rect 595 -236 779 -219
<< metal1 >>
rect -785 236 -589 239
rect -785 219 -779 236
rect -595 219 -589 236
rect -785 216 -589 219
rect -556 236 -360 239
rect -556 219 -550 236
rect -366 219 -360 236
rect -556 216 -360 219
rect -327 236 -131 239
rect -327 219 -321 236
rect -137 219 -131 236
rect -327 216 -131 219
rect -98 236 98 239
rect -98 219 -92 236
rect 92 219 98 236
rect -98 216 98 219
rect 131 236 327 239
rect 131 219 137 236
rect 321 219 327 236
rect 131 216 327 219
rect 360 236 556 239
rect 360 219 366 236
rect 550 219 556 236
rect 360 216 556 219
rect 589 236 785 239
rect 589 219 595 236
rect 779 219 785 236
rect 589 216 785 219
rect -813 194 -790 200
rect -813 -194 -810 194
rect -793 -194 -790 194
rect -813 -200 -790 -194
rect -584 194 -561 200
rect -584 -194 -581 194
rect -564 -194 -561 194
rect -584 -200 -561 -194
rect -355 194 -332 200
rect -355 -194 -352 194
rect -335 -194 -332 194
rect -355 -200 -332 -194
rect -126 194 -103 200
rect -126 -194 -123 194
rect -106 -194 -103 194
rect -126 -200 -103 -194
rect 103 194 126 200
rect 103 -194 106 194
rect 123 -194 126 194
rect 103 -200 126 -194
rect 332 194 355 200
rect 332 -194 335 194
rect 352 -194 355 194
rect 332 -200 355 -194
rect 561 194 584 200
rect 561 -194 564 194
rect 581 -194 584 194
rect 561 -200 584 -194
rect 790 194 813 200
rect 790 -194 793 194
rect 810 -194 813 194
rect 790 -200 813 -194
rect -785 -219 -589 -216
rect -785 -236 -779 -219
rect -595 -236 -589 -219
rect -785 -239 -589 -236
rect -556 -219 -360 -216
rect -556 -236 -550 -219
rect -366 -236 -360 -219
rect -556 -239 -360 -236
rect -327 -219 -131 -216
rect -327 -236 -321 -219
rect -137 -236 -131 -219
rect -327 -239 -131 -236
rect -98 -219 98 -216
rect -98 -236 -92 -219
rect 92 -236 98 -219
rect -98 -239 98 -236
rect 131 -219 327 -216
rect 131 -236 137 -219
rect 321 -236 327 -219
rect 131 -239 327 -236
rect 360 -219 556 -216
rect 360 -236 366 -219
rect 550 -236 556 -219
rect 360 -239 556 -236
rect 589 -219 785 -216
rect 589 -236 595 -219
rect 779 -236 785 -219
rect 589 -239 785 -236
<< properties >>
string FIXED_BBOX -868 -296 868 296
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4 l 2 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
