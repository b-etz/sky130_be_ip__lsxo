magic
tech sky130A
magscale 1 2
timestamp 1713142410
<< pwell >>
rect -957 -610 957 610
<< nmos >>
rect -761 -400 -661 400
rect -603 -400 -503 400
rect -445 -400 -345 400
rect -287 -400 -187 400
rect -129 -400 -29 400
rect 29 -400 129 400
rect 187 -400 287 400
rect 345 -400 445 400
rect 503 -400 603 400
rect 661 -400 761 400
<< ndiff >>
rect -819 388 -761 400
rect -819 -388 -807 388
rect -773 -388 -761 388
rect -819 -400 -761 -388
rect -661 388 -603 400
rect -661 -388 -649 388
rect -615 -388 -603 388
rect -661 -400 -603 -388
rect -503 388 -445 400
rect -503 -388 -491 388
rect -457 -388 -445 388
rect -503 -400 -445 -388
rect -345 388 -287 400
rect -345 -388 -333 388
rect -299 -388 -287 388
rect -345 -400 -287 -388
rect -187 388 -129 400
rect -187 -388 -175 388
rect -141 -388 -129 388
rect -187 -400 -129 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 129 388 187 400
rect 129 -388 141 388
rect 175 -388 187 388
rect 129 -400 187 -388
rect 287 388 345 400
rect 287 -388 299 388
rect 333 -388 345 388
rect 287 -400 345 -388
rect 445 388 503 400
rect 445 -388 457 388
rect 491 -388 503 388
rect 445 -400 503 -388
rect 603 388 661 400
rect 603 -388 615 388
rect 649 -388 661 388
rect 603 -400 661 -388
rect 761 388 819 400
rect 761 -388 773 388
rect 807 -388 819 388
rect 761 -400 819 -388
<< ndiffc >>
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
<< psubdiff >>
rect -921 540 -825 574
rect 825 540 921 574
rect -921 478 -887 540
rect 887 478 921 540
rect -921 -540 -887 -478
rect 887 -540 921 -478
rect -921 -574 -825 -540
rect 825 -574 921 -540
<< psubdiffcont >>
rect -825 540 825 574
rect -921 -478 -887 478
rect 887 -478 921 478
rect -825 -574 825 -540
<< poly >>
rect -761 472 -661 488
rect -761 438 -745 472
rect -677 438 -661 472
rect -761 400 -661 438
rect -603 472 -503 488
rect -603 438 -587 472
rect -519 438 -503 472
rect -603 400 -503 438
rect -445 472 -345 488
rect -445 438 -429 472
rect -361 438 -345 472
rect -445 400 -345 438
rect -287 472 -187 488
rect -287 438 -271 472
rect -203 438 -187 472
rect -287 400 -187 438
rect -129 472 -29 488
rect -129 438 -113 472
rect -45 438 -29 472
rect -129 400 -29 438
rect 29 472 129 488
rect 29 438 45 472
rect 113 438 129 472
rect 29 400 129 438
rect 187 472 287 488
rect 187 438 203 472
rect 271 438 287 472
rect 187 400 287 438
rect 345 472 445 488
rect 345 438 361 472
rect 429 438 445 472
rect 345 400 445 438
rect 503 472 603 488
rect 503 438 519 472
rect 587 438 603 472
rect 503 400 603 438
rect 661 472 761 488
rect 661 438 677 472
rect 745 438 761 472
rect 661 400 761 438
rect -761 -438 -661 -400
rect -761 -472 -745 -438
rect -677 -472 -661 -438
rect -761 -488 -661 -472
rect -603 -438 -503 -400
rect -603 -472 -587 -438
rect -519 -472 -503 -438
rect -603 -488 -503 -472
rect -445 -438 -345 -400
rect -445 -472 -429 -438
rect -361 -472 -345 -438
rect -445 -488 -345 -472
rect -287 -438 -187 -400
rect -287 -472 -271 -438
rect -203 -472 -187 -438
rect -287 -488 -187 -472
rect -129 -438 -29 -400
rect -129 -472 -113 -438
rect -45 -472 -29 -438
rect -129 -488 -29 -472
rect 29 -438 129 -400
rect 29 -472 45 -438
rect 113 -472 129 -438
rect 29 -488 129 -472
rect 187 -438 287 -400
rect 187 -472 203 -438
rect 271 -472 287 -438
rect 187 -488 287 -472
rect 345 -438 445 -400
rect 345 -472 361 -438
rect 429 -472 445 -438
rect 345 -488 445 -472
rect 503 -438 603 -400
rect 503 -472 519 -438
rect 587 -472 603 -438
rect 503 -488 603 -472
rect 661 -438 761 -400
rect 661 -472 677 -438
rect 745 -472 761 -438
rect 661 -488 761 -472
<< polycont >>
rect -745 438 -677 472
rect -587 438 -519 472
rect -429 438 -361 472
rect -271 438 -203 472
rect -113 438 -45 472
rect 45 438 113 472
rect 203 438 271 472
rect 361 438 429 472
rect 519 438 587 472
rect 677 438 745 472
rect -745 -472 -677 -438
rect -587 -472 -519 -438
rect -429 -472 -361 -438
rect -271 -472 -203 -438
rect -113 -472 -45 -438
rect 45 -472 113 -438
rect 203 -472 271 -438
rect 361 -472 429 -438
rect 519 -472 587 -438
rect 677 -472 745 -438
<< locali >>
rect -921 540 -825 574
rect 825 540 921 574
rect -921 478 -887 540
rect 887 478 921 540
rect -761 438 -745 472
rect -677 438 -661 472
rect -603 438 -587 472
rect -519 438 -503 472
rect -445 438 -429 472
rect -361 438 -345 472
rect -287 438 -271 472
rect -203 438 -187 472
rect -129 438 -113 472
rect -45 438 -29 472
rect 29 438 45 472
rect 113 438 129 472
rect 187 438 203 472
rect 271 438 287 472
rect 345 438 361 472
rect 429 438 445 472
rect 503 438 519 472
rect 587 438 603 472
rect 661 438 677 472
rect 745 438 761 472
rect -807 388 -773 404
rect -807 -404 -773 -388
rect -649 388 -615 404
rect -649 -404 -615 -388
rect -491 388 -457 404
rect -491 -404 -457 -388
rect -333 388 -299 404
rect -333 -404 -299 -388
rect -175 388 -141 404
rect -175 -404 -141 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 141 388 175 404
rect 141 -404 175 -388
rect 299 388 333 404
rect 299 -404 333 -388
rect 457 388 491 404
rect 457 -404 491 -388
rect 615 388 649 404
rect 615 -404 649 -388
rect 773 388 807 404
rect 773 -404 807 -388
rect -761 -472 -745 -438
rect -677 -472 -661 -438
rect -603 -472 -587 -438
rect -519 -472 -503 -438
rect -445 -472 -429 -438
rect -361 -472 -345 -438
rect -287 -472 -271 -438
rect -203 -472 -187 -438
rect -129 -472 -113 -438
rect -45 -472 -29 -438
rect 29 -472 45 -438
rect 113 -472 129 -438
rect 187 -472 203 -438
rect 271 -472 287 -438
rect 345 -472 361 -438
rect 429 -472 445 -438
rect 503 -472 519 -438
rect 587 -472 603 -438
rect 661 -472 677 -438
rect 745 -472 761 -438
rect -921 -540 -887 -478
rect 887 -540 921 -478
rect -921 -574 -825 -540
rect 825 -574 921 -540
<< viali >>
rect -745 438 -677 472
rect -587 438 -519 472
rect -429 438 -361 472
rect -271 438 -203 472
rect -113 438 -45 472
rect 45 438 113 472
rect 203 438 271 472
rect 361 438 429 472
rect 519 438 587 472
rect 677 438 745 472
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
rect -745 -472 -677 -438
rect -587 -472 -519 -438
rect -429 -472 -361 -438
rect -271 -472 -203 -438
rect -113 -472 -45 -438
rect 45 -472 113 -438
rect 203 -472 271 -438
rect 361 -472 429 -438
rect 519 -472 587 -438
rect 677 -472 745 -438
<< metal1 >>
rect -757 472 -665 478
rect -757 438 -745 472
rect -677 438 -665 472
rect -757 432 -665 438
rect -599 472 -507 478
rect -599 438 -587 472
rect -519 438 -507 472
rect -599 432 -507 438
rect -441 472 -349 478
rect -441 438 -429 472
rect -361 438 -349 472
rect -441 432 -349 438
rect -283 472 -191 478
rect -283 438 -271 472
rect -203 438 -191 472
rect -283 432 -191 438
rect -125 472 -33 478
rect -125 438 -113 472
rect -45 438 -33 472
rect -125 432 -33 438
rect 33 472 125 478
rect 33 438 45 472
rect 113 438 125 472
rect 33 432 125 438
rect 191 472 283 478
rect 191 438 203 472
rect 271 438 283 472
rect 191 432 283 438
rect 349 472 441 478
rect 349 438 361 472
rect 429 438 441 472
rect 349 432 441 438
rect 507 472 599 478
rect 507 438 519 472
rect 587 438 599 472
rect 507 432 599 438
rect 665 472 757 478
rect 665 438 677 472
rect 745 438 757 472
rect 665 432 757 438
rect -813 388 -767 400
rect -813 -388 -807 388
rect -773 -388 -767 388
rect -813 -400 -767 -388
rect -655 388 -609 400
rect -655 -388 -649 388
rect -615 -388 -609 388
rect -655 -400 -609 -388
rect -497 388 -451 400
rect -497 -388 -491 388
rect -457 -388 -451 388
rect -497 -400 -451 -388
rect -339 388 -293 400
rect -339 -388 -333 388
rect -299 -388 -293 388
rect -339 -400 -293 -388
rect -181 388 -135 400
rect -181 -388 -175 388
rect -141 -388 -135 388
rect -181 -400 -135 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 135 388 181 400
rect 135 -388 141 388
rect 175 -388 181 388
rect 135 -400 181 -388
rect 293 388 339 400
rect 293 -388 299 388
rect 333 -388 339 388
rect 293 -400 339 -388
rect 451 388 497 400
rect 451 -388 457 388
rect 491 -388 497 388
rect 451 -400 497 -388
rect 609 388 655 400
rect 609 -388 615 388
rect 649 -388 655 388
rect 609 -400 655 -388
rect 767 388 813 400
rect 767 -388 773 388
rect 807 -388 813 388
rect 767 -400 813 -388
rect -757 -438 -665 -432
rect -757 -472 -745 -438
rect -677 -472 -665 -438
rect -757 -478 -665 -472
rect -599 -438 -507 -432
rect -599 -472 -587 -438
rect -519 -472 -507 -438
rect -599 -478 -507 -472
rect -441 -438 -349 -432
rect -441 -472 -429 -438
rect -361 -472 -349 -438
rect -441 -478 -349 -472
rect -283 -438 -191 -432
rect -283 -472 -271 -438
rect -203 -472 -191 -438
rect -283 -478 -191 -472
rect -125 -438 -33 -432
rect -125 -472 -113 -438
rect -45 -472 -33 -438
rect -125 -478 -33 -472
rect 33 -438 125 -432
rect 33 -472 45 -438
rect 113 -472 125 -438
rect 33 -478 125 -472
rect 191 -438 283 -432
rect 191 -472 203 -438
rect 271 -472 283 -438
rect 191 -478 283 -472
rect 349 -438 441 -432
rect 349 -472 361 -438
rect 429 -472 441 -438
rect 349 -478 441 -472
rect 507 -438 599 -432
rect 507 -472 519 -438
rect 587 -472 599 -438
rect 507 -478 599 -472
rect 665 -438 757 -432
rect 665 -472 677 -438
rect 745 -472 757 -438
rect 665 -478 757 -472
<< properties >>
string FIXED_BBOX -904 -557 904 557
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.0 l 0.5 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
