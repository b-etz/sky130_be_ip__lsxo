magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< pwell >>
rect -948 -26582 948 26582
<< psubdiff >>
rect -912 26512 -816 26546
rect 816 26512 912 26546
rect -912 26450 -878 26512
rect 878 26450 912 26512
rect -912 -26512 -878 -26450
rect 878 -26512 912 -26450
rect -912 -26546 -816 -26512
rect 816 -26546 912 -26512
<< psubdiffcont >>
rect -816 26512 816 26546
rect -912 -26450 -878 26450
rect 878 -26450 912 26450
rect -816 -26546 816 -26512
<< xpolycontact >>
rect -782 25984 -712 26416
rect -782 -26416 -712 -25984
rect -616 25984 -546 26416
rect -616 -26416 -546 -25984
rect -450 25984 -380 26416
rect -450 -26416 -380 -25984
rect -284 25984 -214 26416
rect -284 -26416 -214 -25984
rect -118 25984 -48 26416
rect -118 -26416 -48 -25984
rect 48 25984 118 26416
rect 48 -26416 118 -25984
rect 214 25984 284 26416
rect 214 -26416 284 -25984
rect 380 25984 450 26416
rect 380 -26416 450 -25984
rect 546 25984 616 26416
rect 546 -26416 616 -25984
rect 712 25984 782 26416
rect 712 -26416 782 -25984
<< xpolyres >>
rect -782 -25984 -712 25984
rect -616 -25984 -546 25984
rect -450 -25984 -380 25984
rect -284 -25984 -214 25984
rect -118 -25984 -48 25984
rect 48 -25984 118 25984
rect 214 -25984 284 25984
rect 380 -25984 450 25984
rect 546 -25984 616 25984
rect 712 -25984 782 25984
<< locali >>
rect -912 26512 -816 26546
rect 816 26512 912 26546
rect -912 26450 -878 26512
rect 878 26450 912 26512
rect -912 -26512 -878 -26450
rect 878 -26512 912 -26450
rect -912 -26546 -816 -26512
rect 816 -26546 912 -26512
<< viali >>
rect -766 26001 -728 26398
rect -600 26001 -562 26398
rect -434 26001 -396 26398
rect -268 26001 -230 26398
rect -102 26001 -64 26398
rect 64 26001 102 26398
rect 230 26001 268 26398
rect 396 26001 434 26398
rect 562 26001 600 26398
rect 728 26001 766 26398
rect -766 -26398 -728 -26001
rect -600 -26398 -562 -26001
rect -434 -26398 -396 -26001
rect -268 -26398 -230 -26001
rect -102 -26398 -64 -26001
rect 64 -26398 102 -26001
rect 230 -26398 268 -26001
rect 396 -26398 434 -26001
rect 562 -26398 600 -26001
rect 728 -26398 766 -26001
<< metal1 >>
rect -772 26398 -722 26410
rect -772 26001 -766 26398
rect -728 26001 -722 26398
rect -772 25989 -722 26001
rect -606 26398 -556 26410
rect -606 26001 -600 26398
rect -562 26001 -556 26398
rect -606 25989 -556 26001
rect -440 26398 -390 26410
rect -440 26001 -434 26398
rect -396 26001 -390 26398
rect -440 25989 -390 26001
rect -274 26398 -224 26410
rect -274 26001 -268 26398
rect -230 26001 -224 26398
rect -274 25989 -224 26001
rect -108 26398 -58 26410
rect -108 26001 -102 26398
rect -64 26001 -58 26398
rect -108 25989 -58 26001
rect 58 26398 108 26410
rect 58 26001 64 26398
rect 102 26001 108 26398
rect 58 25989 108 26001
rect 224 26398 274 26410
rect 224 26001 230 26398
rect 268 26001 274 26398
rect 224 25989 274 26001
rect 390 26398 440 26410
rect 390 26001 396 26398
rect 434 26001 440 26398
rect 390 25989 440 26001
rect 556 26398 606 26410
rect 556 26001 562 26398
rect 600 26001 606 26398
rect 556 25989 606 26001
rect 722 26398 772 26410
rect 722 26001 728 26398
rect 766 26001 772 26398
rect 722 25989 772 26001
rect -772 -26001 -722 -25989
rect -772 -26398 -766 -26001
rect -728 -26398 -722 -26001
rect -772 -26410 -722 -26398
rect -606 -26001 -556 -25989
rect -606 -26398 -600 -26001
rect -562 -26398 -556 -26001
rect -606 -26410 -556 -26398
rect -440 -26001 -390 -25989
rect -440 -26398 -434 -26001
rect -396 -26398 -390 -26001
rect -440 -26410 -390 -26398
rect -274 -26001 -224 -25989
rect -274 -26398 -268 -26001
rect -230 -26398 -224 -26001
rect -274 -26410 -224 -26398
rect -108 -26001 -58 -25989
rect -108 -26398 -102 -26001
rect -64 -26398 -58 -26001
rect -108 -26410 -58 -26398
rect 58 -26001 108 -25989
rect 58 -26398 64 -26001
rect 102 -26398 108 -26001
rect 58 -26410 108 -26398
rect 224 -26001 274 -25989
rect 224 -26398 230 -26001
rect 268 -26398 274 -26001
rect 224 -26410 274 -26398
rect 390 -26001 440 -25989
rect 390 -26398 396 -26001
rect 434 -26398 440 -26001
rect 390 -26410 440 -26398
rect 556 -26001 606 -25989
rect 556 -26398 562 -26001
rect 600 -26398 606 -26001
rect 556 -26410 606 -26398
rect 722 -26001 772 -25989
rect 722 -26398 728 -26001
rect 766 -26398 772 -26001
rect 722 -26410 772 -26398
<< properties >>
string FIXED_BBOX -895 -26529 895 26529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 260.0 m 1 nx 10 wmin 0.350 lmin 0.50 rho 2000 val 1.486meg dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
