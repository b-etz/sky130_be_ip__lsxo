magic
tech sky130A
magscale 1 2
timestamp 1713224303
<< dnwell >>
rect 1926 -9006 6422 -3446
rect 8780 -10312 25248 -4220
rect 1706 -23624 25490 -11618
<< nwell >>
rect 3211 -1638 3532 -1194
rect 4798 -1638 5119 -1194
rect 3216 -2542 3808 -1904
rect 4528 -2542 5120 -1904
rect 7326 -3206 9240 -1968
rect 11222 -3266 11838 -1872
rect 14249 -2892 14570 -1620
rect 14830 -2577 22174 -2011
rect 1846 -3652 6502 -3366
rect 1846 -8800 2132 -3652
rect 2552 -6530 3868 -5132
rect 4468 -6530 5784 -5132
rect 3614 -8352 4862 -6958
rect 6216 -8800 6502 -3652
rect 1846 -9086 6502 -8800
rect 8700 -4426 25328 -4140
rect 8700 -10106 8986 -4426
rect 10486 -7136 15282 -5770
rect 16002 -7194 18292 -5800
rect 18732 -6866 20724 -6328
rect 21216 -6958 22066 -6192
rect 22912 -6846 24150 -6254
rect 9578 -9276 10116 -7284
rect 25042 -10106 25328 -4426
rect 8700 -10392 25328 -10106
rect 1626 -11824 25570 -11538
rect 1626 -23418 1912 -11824
rect 22304 -18036 24626 -12496
rect 21178 -23158 21544 -22792
rect 22604 -23160 22970 -22794
rect 25284 -23418 25570 -11824
rect 1626 -23704 25570 -23418
<< pwell >>
rect 2750 -1180 3116 -814
rect 5220 -1180 5586 -814
rect 2988 -1321 3145 -1235
rect 2971 -1355 3127 -1325
rect 2933 -1389 3127 -1355
rect 2971 -1599 3127 -1389
rect 5185 -1321 5342 -1235
rect 5203 -1355 5359 -1325
rect 5203 -1389 5397 -1355
rect 5203 -1599 5359 -1389
rect 14026 -1747 14183 -1661
rect 14009 -1780 14191 -1751
rect 13971 -1814 14191 -1780
rect 2616 -2532 3208 -1912
rect 5128 -2532 5720 -1912
rect 9252 -3202 11166 -1982
rect 12564 -3248 13084 -2056
rect 14009 -2482 14191 -1814
rect 14009 -2515 14145 -2490
rect 13971 -2549 14145 -2515
rect 14009 -2851 14145 -2549
rect 14989 -1771 15023 -1733
rect 15541 -1771 15575 -1733
rect 17749 -1771 17783 -1733
rect 19957 -1771 19991 -1733
rect 14871 -1945 14957 -1788
rect 14974 -1907 15356 -1771
rect 15423 -1945 15509 -1788
rect 15513 -1907 17616 -1771
rect 16415 -1951 16601 -1907
rect 17145 -1953 17616 -1907
rect 17631 -1945 17717 -1788
rect 17721 -1907 19824 -1771
rect 18623 -1951 18809 -1907
rect 19353 -1953 19824 -1907
rect 19839 -1945 19925 -1788
rect 19929 -1907 22032 -1771
rect 20831 -1951 21017 -1907
rect 21561 -1953 22032 -1907
rect 22047 -1945 22133 -1788
rect 14871 -2800 14957 -2643
rect 14974 -2817 15356 -2681
rect 15423 -2800 15509 -2643
rect 16415 -2681 16601 -2637
rect 17145 -2681 17616 -2635
rect 15513 -2817 17616 -2681
rect 17631 -2800 17717 -2643
rect 18623 -2681 18809 -2637
rect 19353 -2681 19824 -2635
rect 17721 -2817 19824 -2681
rect 19839 -2800 19925 -2643
rect 20831 -2681 21017 -2637
rect 21561 -2681 22032 -2635
rect 19929 -2817 22032 -2681
rect 22047 -2800 22133 -2643
rect 14989 -2855 15023 -2817
rect 15541 -2855 15575 -2817
rect 17749 -2855 17783 -2817
rect 19957 -2855 19991 -2817
rect 14960 -3476 16152 -2956
rect 2500 -4984 3920 -3868
rect 4416 -4984 5836 -3868
rect 2269 -8311 3457 -6995
rect 10430 -5616 15332 -4700
rect 16064 -5748 18230 -4528
rect 18752 -5844 20744 -5324
rect 21216 -5926 22066 -5196
rect 23224 -5844 23794 -5252
rect 8998 -9542 9518 -7550
rect 10454 -9998 24818 -7272
rect 7098 -12708 7754 -11992
rect 8040 -12652 13412 -12052
rect 2968 -13656 19132 -12756
rect 1966 -18246 19530 -13694
rect 19740 -15686 21966 -12518
rect 20206 -18156 21522 -15862
rect 1964 -22670 25128 -18284
rect 21040 -22792 21682 -22670
rect 20322 -23168 20688 -22802
rect 21040 -23158 21178 -22792
rect 21544 -23158 21682 -22792
rect 21040 -23296 21682 -23158
rect 22466 -22794 23108 -22670
rect 22466 -23160 22604 -22794
rect 22970 -23160 23108 -22794
rect 22466 -23298 23108 -23160
rect 23430 -23170 23796 -22804
<< nmos >>
rect 2812 -2322 3012 -2122
rect 5324 -2322 5524 -2122
rect 9448 -2992 9548 -2192
rect 9606 -2992 9706 -2192
rect 9764 -2992 9864 -2192
rect 9922 -2992 10022 -2192
rect 10080 -2992 10180 -2192
rect 10238 -2992 10338 -2192
rect 10396 -2992 10496 -2192
rect 10554 -2992 10654 -2192
rect 10712 -2992 10812 -2192
rect 10870 -2992 10970 -2192
rect 12774 -3052 12874 -2252
rect 15156 -3266 15956 -3166
rect 16260 -5538 16660 -4738
rect 16718 -5538 17118 -4738
rect 17176 -5538 17576 -4738
rect 17634 -5538 18034 -4738
rect 18948 -5634 20548 -5534
rect 21412 -5506 21612 -5406
rect 21670 -5506 21870 -5406
rect 21412 -5716 21612 -5616
rect 21670 -5716 21870 -5616
rect 23434 -5648 23584 -5448
rect 9208 -9346 9308 -7746
<< scnmos >>
rect 2997 -1433 3101 -1403
rect 5229 -1433 5333 -1403
rect 2997 -1521 3101 -1491
rect 5229 -1521 5333 -1491
rect 14035 -1859 14165 -1829
rect 14035 -1955 14165 -1925
rect 15053 -1881 15083 -1797
rect 15125 -1881 15155 -1797
rect 15247 -1881 15277 -1797
rect 14035 -2027 14165 -1997
rect 14035 -2215 14165 -2185
rect 15591 -1881 15621 -1797
rect 15675 -1881 15705 -1797
rect 15930 -1881 15960 -1797
rect 16025 -1869 16055 -1797
rect 16121 -1869 16151 -1797
rect 16287 -1881 16317 -1797
rect 16359 -1881 16389 -1797
rect 14035 -2311 14165 -2281
rect 16491 -1925 16521 -1797
rect 16590 -1869 16620 -1797
rect 16699 -1869 16729 -1797
rect 16795 -1881 16825 -1797
rect 16944 -1881 16974 -1797
rect 17035 -1881 17065 -1797
rect 17223 -1927 17253 -1797
rect 17411 -1881 17441 -1797
rect 17508 -1927 17538 -1797
rect 17799 -1881 17829 -1797
rect 17883 -1881 17913 -1797
rect 18138 -1881 18168 -1797
rect 18233 -1869 18263 -1797
rect 18329 -1869 18359 -1797
rect 18495 -1881 18525 -1797
rect 18567 -1881 18597 -1797
rect 18699 -1925 18729 -1797
rect 18798 -1869 18828 -1797
rect 18907 -1869 18937 -1797
rect 19003 -1881 19033 -1797
rect 19152 -1881 19182 -1797
rect 19243 -1881 19273 -1797
rect 19431 -1927 19461 -1797
rect 19619 -1881 19649 -1797
rect 19716 -1927 19746 -1797
rect 20007 -1881 20037 -1797
rect 20091 -1881 20121 -1797
rect 20346 -1881 20376 -1797
rect 20441 -1869 20471 -1797
rect 20537 -1869 20567 -1797
rect 20703 -1881 20733 -1797
rect 20775 -1881 20805 -1797
rect 20907 -1925 20937 -1797
rect 21006 -1869 21036 -1797
rect 21115 -1869 21145 -1797
rect 21211 -1881 21241 -1797
rect 21360 -1881 21390 -1797
rect 21451 -1881 21481 -1797
rect 21639 -1927 21669 -1797
rect 21827 -1881 21857 -1797
rect 21924 -1927 21954 -1797
rect 14035 -2404 14165 -2374
rect 14035 -2598 14119 -2568
rect 14035 -2701 14119 -2671
rect 14035 -2773 14119 -2743
rect 15053 -2791 15083 -2707
rect 15125 -2791 15155 -2707
rect 15247 -2791 15277 -2707
rect 15591 -2791 15621 -2707
rect 15675 -2791 15705 -2707
rect 15930 -2791 15960 -2707
rect 16025 -2791 16055 -2719
rect 16121 -2791 16151 -2719
rect 16287 -2791 16317 -2707
rect 16359 -2791 16389 -2707
rect 16491 -2791 16521 -2663
rect 16590 -2791 16620 -2719
rect 16699 -2791 16729 -2719
rect 16795 -2791 16825 -2707
rect 16944 -2791 16974 -2707
rect 17035 -2791 17065 -2707
rect 17223 -2791 17253 -2661
rect 17411 -2791 17441 -2707
rect 17508 -2791 17538 -2661
rect 17799 -2791 17829 -2707
rect 17883 -2791 17913 -2707
rect 18138 -2791 18168 -2707
rect 18233 -2791 18263 -2719
rect 18329 -2791 18359 -2719
rect 18495 -2791 18525 -2707
rect 18567 -2791 18597 -2707
rect 18699 -2791 18729 -2663
rect 18798 -2791 18828 -2719
rect 18907 -2791 18937 -2719
rect 19003 -2791 19033 -2707
rect 19152 -2791 19182 -2707
rect 19243 -2791 19273 -2707
rect 19431 -2791 19461 -2661
rect 19619 -2791 19649 -2707
rect 19716 -2791 19746 -2661
rect 20007 -2791 20037 -2707
rect 20091 -2791 20121 -2707
rect 20346 -2791 20376 -2707
rect 20441 -2791 20471 -2719
rect 20537 -2791 20567 -2719
rect 20703 -2791 20733 -2707
rect 20775 -2791 20805 -2707
rect 20907 -2791 20937 -2663
rect 21006 -2791 21036 -2719
rect 21115 -2791 21145 -2719
rect 21211 -2791 21241 -2707
rect 21360 -2791 21390 -2707
rect 21451 -2791 21481 -2707
rect 21639 -2791 21669 -2661
rect 21827 -2791 21857 -2707
rect 21924 -2791 21954 -2661
<< pmos >>
rect 3412 -2323 3612 -2123
rect 4724 -2323 4924 -2123
rect 7522 -2987 7622 -2187
rect 7680 -2987 7780 -2187
rect 7838 -2987 7938 -2187
rect 7996 -2987 8096 -2187
rect 8154 -2987 8254 -2187
rect 8312 -2987 8412 -2187
rect 8470 -2987 8570 -2187
rect 8628 -2987 8728 -2187
rect 8786 -2987 8886 -2187
rect 8944 -2987 9044 -2187
rect 10682 -6389 11082 -5989
rect 11254 -6389 11654 -5989
rect 11826 -6389 12226 -5989
rect 12398 -6389 12798 -5989
rect 12970 -6389 13370 -5989
rect 13542 -6389 13942 -5989
rect 14114 -6389 14514 -5989
rect 14686 -6389 15086 -5989
rect 10682 -6917 11082 -6517
rect 11254 -6917 11654 -6517
rect 11826 -6917 12226 -6517
rect 12398 -6917 12798 -6517
rect 12970 -6917 13370 -6517
rect 13542 -6917 13942 -6517
rect 14114 -6917 14514 -6517
rect 14686 -6917 15086 -6517
rect 18928 -6647 20528 -6547
rect 21412 -6511 21612 -6411
rect 21670 -6511 21870 -6411
rect 21412 -6739 21612 -6639
rect 21670 -6739 21870 -6639
rect 23131 -6650 23931 -6450
rect 9797 -9080 9897 -7480
<< scpmoshvt >>
rect 3289 -1433 3447 -1403
rect 4883 -1433 5041 -1403
rect 3289 -1521 3447 -1491
rect 4883 -1521 5041 -1491
rect 14285 -1859 14485 -1829
rect 14285 -1943 14485 -1913
rect 14285 -2027 14485 -1997
rect 14285 -2215 14485 -2185
rect 15053 -2247 15083 -2163
rect 15141 -2247 15171 -2163
rect 15295 -2247 15325 -2119
rect 15591 -2241 15621 -2113
rect 15675 -2241 15705 -2113
rect 15942 -2247 15972 -2163
rect 16034 -2247 16064 -2163
rect 16133 -2247 16163 -2163
rect 16273 -2247 16303 -2163
rect 16370 -2247 16400 -2163
rect 16567 -2247 16597 -2079
rect 16666 -2247 16696 -2163
rect 16752 -2247 16782 -2163
rect 16836 -2247 16866 -2163
rect 16944 -2247 16974 -2163
rect 17028 -2247 17058 -2163
rect 17192 -2247 17222 -2047
rect 17411 -2247 17441 -2119
rect 17508 -2247 17538 -2047
rect 17799 -2241 17829 -2113
rect 17883 -2241 17913 -2113
rect 18150 -2247 18180 -2163
rect 18242 -2247 18272 -2163
rect 18341 -2247 18371 -2163
rect 18481 -2247 18511 -2163
rect 18578 -2247 18608 -2163
rect 18775 -2247 18805 -2079
rect 18874 -2247 18904 -2163
rect 18960 -2247 18990 -2163
rect 19044 -2247 19074 -2163
rect 19152 -2247 19182 -2163
rect 19236 -2247 19266 -2163
rect 19400 -2247 19430 -2047
rect 19619 -2247 19649 -2119
rect 19716 -2247 19746 -2047
rect 20007 -2241 20037 -2113
rect 20091 -2241 20121 -2113
rect 20358 -2247 20388 -2163
rect 20450 -2247 20480 -2163
rect 20549 -2247 20579 -2163
rect 20689 -2247 20719 -2163
rect 20786 -2247 20816 -2163
rect 20983 -2247 21013 -2079
rect 21082 -2247 21112 -2163
rect 21168 -2247 21198 -2163
rect 21252 -2247 21282 -2163
rect 21360 -2247 21390 -2163
rect 21444 -2247 21474 -2163
rect 21608 -2247 21638 -2047
rect 21827 -2247 21857 -2119
rect 21924 -2247 21954 -2047
rect 14285 -2311 14485 -2281
rect 14285 -2404 14485 -2374
rect 15053 -2425 15083 -2341
rect 15141 -2425 15171 -2341
rect 15295 -2469 15325 -2341
rect 14401 -2598 14485 -2568
rect 14357 -2701 14485 -2671
rect 15591 -2475 15621 -2347
rect 15675 -2475 15705 -2347
rect 15942 -2425 15972 -2341
rect 16034 -2425 16064 -2341
rect 16133 -2425 16163 -2341
rect 16273 -2425 16303 -2341
rect 16370 -2425 16400 -2341
rect 14357 -2773 14485 -2743
rect 16567 -2509 16597 -2341
rect 16666 -2425 16696 -2341
rect 16752 -2425 16782 -2341
rect 16836 -2425 16866 -2341
rect 16944 -2425 16974 -2341
rect 17028 -2425 17058 -2341
rect 17192 -2541 17222 -2341
rect 17411 -2469 17441 -2341
rect 17508 -2541 17538 -2341
rect 17799 -2475 17829 -2347
rect 17883 -2475 17913 -2347
rect 18150 -2425 18180 -2341
rect 18242 -2425 18272 -2341
rect 18341 -2425 18371 -2341
rect 18481 -2425 18511 -2341
rect 18578 -2425 18608 -2341
rect 18775 -2509 18805 -2341
rect 18874 -2425 18904 -2341
rect 18960 -2425 18990 -2341
rect 19044 -2425 19074 -2341
rect 19152 -2425 19182 -2341
rect 19236 -2425 19266 -2341
rect 19400 -2541 19430 -2341
rect 19619 -2469 19649 -2341
rect 19716 -2541 19746 -2341
rect 20007 -2475 20037 -2347
rect 20091 -2475 20121 -2347
rect 20358 -2425 20388 -2341
rect 20450 -2425 20480 -2341
rect 20549 -2425 20579 -2341
rect 20689 -2425 20719 -2341
rect 20786 -2425 20816 -2341
rect 20983 -2509 21013 -2341
rect 21082 -2425 21112 -2341
rect 21168 -2425 21198 -2341
rect 21252 -2425 21282 -2341
rect 21360 -2425 21390 -2341
rect 21444 -2425 21474 -2341
rect 21608 -2541 21638 -2341
rect 21827 -2469 21857 -2341
rect 21924 -2541 21954 -2341
<< mvnmos >>
rect 2728 -4726 2828 -4126
rect 2886 -4726 2986 -4126
rect 3434 -4726 3534 -4126
rect 3592 -4726 3692 -4126
rect 4644 -4726 4744 -4126
rect 4802 -4726 4902 -4126
rect 5350 -4726 5450 -4126
rect 5508 -4726 5608 -4126
rect 2497 -8053 2597 -7253
rect 2655 -8053 2755 -7253
rect 2813 -8053 2913 -7253
rect 2971 -8053 3071 -7253
rect 3129 -8053 3229 -7253
rect 10658 -5358 11058 -4958
rect 11236 -5358 11636 -4958
rect 11814 -5358 12214 -4958
rect 12392 -5358 12792 -4958
rect 12970 -5358 13370 -4958
rect 13548 -5358 13948 -4958
rect 14126 -5358 14526 -4958
rect 14704 -5358 15104 -4958
rect 7326 -12450 7526 -12250
rect 8268 -12394 9868 -12310
rect 9926 -12394 11526 -12310
rect 11584 -12394 13184 -12310
rect 19998 -13146 20798 -12746
rect 20908 -13146 21708 -12746
rect 19998 -13724 20798 -13324
rect 20908 -13724 21708 -13324
rect 19998 -14302 20798 -13902
rect 20908 -14302 21708 -13902
rect 19998 -14880 20798 -14480
rect 20908 -14880 21708 -14480
rect 19998 -15458 20798 -15058
rect 20908 -15458 21708 -15058
rect 20464 -16190 21264 -16090
rect 20464 -16348 21264 -16248
rect 20464 -16506 21264 -16406
rect 20464 -16664 21264 -16564
rect 20464 -16822 21264 -16722
rect 20464 -16980 21264 -16880
rect 20464 -17138 21264 -17038
rect 20464 -17296 21264 -17196
rect 20464 -17454 21264 -17354
rect 20464 -17612 21264 -17512
rect 20464 -17770 21264 -17670
rect 20464 -17928 21264 -17828
<< mvpmos >>
rect 11480 -2969 11580 -2169
rect 2810 -5629 3610 -5429
rect 2810 -6233 3610 -6033
rect 4726 -5629 5526 -5429
rect 4726 -6233 5526 -6033
rect 3872 -8055 3972 -7255
rect 4030 -8055 4130 -7255
rect 4188 -8055 4288 -7255
rect 4346 -8055 4446 -7255
rect 4504 -8055 4604 -7255
rect 16260 -6897 16660 -6097
rect 16718 -6897 17118 -6097
rect 17176 -6897 17576 -6097
rect 17634 -6897 18034 -6097
rect 22601 -13154 23401 -12754
rect 23529 -13154 24329 -12754
rect 22601 -13732 23401 -13332
rect 23529 -13732 24329 -13332
rect 22601 -14310 23401 -13910
rect 23529 -14310 24329 -13910
rect 22601 -14888 23401 -14488
rect 23529 -14888 24329 -14488
rect 22601 -15466 23401 -15066
rect 23529 -15466 24329 -15066
rect 22601 -16044 23401 -15644
rect 23529 -16044 24329 -15644
rect 22601 -16622 23401 -16222
rect 23529 -16622 24329 -16222
rect 22601 -17200 23401 -16800
rect 23529 -17200 24329 -16800
rect 22601 -17778 23401 -17378
rect 23529 -17778 24329 -17378
<< ndiff >>
rect 2997 -1359 3101 -1351
rect 2997 -1393 3022 -1359
rect 3056 -1393 3101 -1359
rect 2997 -1403 3101 -1393
rect 5229 -1359 5333 -1351
rect 5229 -1393 5274 -1359
rect 5308 -1393 5333 -1359
rect 5229 -1403 5333 -1393
rect 2997 -1445 3101 -1433
rect 2997 -1479 3009 -1445
rect 3043 -1479 3101 -1445
rect 2997 -1491 3101 -1479
rect 5229 -1445 5333 -1433
rect 5229 -1479 5287 -1445
rect 5321 -1479 5333 -1445
rect 5229 -1491 5333 -1479
rect 2997 -1531 3101 -1521
rect 2997 -1565 3039 -1531
rect 3073 -1565 3101 -1531
rect 2997 -1573 3101 -1565
rect 5229 -1531 5333 -1521
rect 5229 -1565 5257 -1531
rect 5291 -1565 5333 -1531
rect 5229 -1573 5333 -1565
rect 14035 -1785 14165 -1777
rect 14035 -1819 14083 -1785
rect 14117 -1819 14165 -1785
rect 14035 -1829 14165 -1819
rect 14035 -1869 14165 -1859
rect 14035 -1903 14059 -1869
rect 14093 -1903 14165 -1869
rect 14035 -1925 14165 -1903
rect 2754 -2134 2812 -2122
rect 2754 -2310 2766 -2134
rect 2800 -2310 2812 -2134
rect 2754 -2322 2812 -2310
rect 3012 -2134 3070 -2122
rect 3012 -2310 3024 -2134
rect 3058 -2310 3070 -2134
rect 3012 -2322 3070 -2310
rect 15000 -1822 15053 -1797
rect 15000 -1856 15008 -1822
rect 15042 -1856 15053 -1822
rect 15000 -1881 15053 -1856
rect 15083 -1881 15125 -1797
rect 15155 -1805 15247 -1797
rect 15155 -1839 15179 -1805
rect 15213 -1839 15247 -1805
rect 15155 -1881 15247 -1839
rect 15277 -1809 15330 -1797
rect 15277 -1843 15288 -1809
rect 15322 -1843 15330 -1809
rect 15277 -1881 15330 -1843
rect 5266 -2134 5324 -2122
rect 5266 -2310 5278 -2134
rect 5312 -2310 5324 -2134
rect 5266 -2322 5324 -2310
rect 5524 -2134 5582 -2122
rect 5524 -2310 5536 -2134
rect 5570 -2310 5582 -2134
rect 5524 -2322 5582 -2310
rect 9390 -2204 9448 -2192
rect 9390 -2980 9402 -2204
rect 9436 -2980 9448 -2204
rect 9390 -2992 9448 -2980
rect 9548 -2204 9606 -2192
rect 9548 -2980 9560 -2204
rect 9594 -2980 9606 -2204
rect 9548 -2992 9606 -2980
rect 9706 -2204 9764 -2192
rect 9706 -2980 9718 -2204
rect 9752 -2980 9764 -2204
rect 9706 -2992 9764 -2980
rect 9864 -2204 9922 -2192
rect 9864 -2980 9876 -2204
rect 9910 -2980 9922 -2204
rect 9864 -2992 9922 -2980
rect 10022 -2204 10080 -2192
rect 10022 -2980 10034 -2204
rect 10068 -2980 10080 -2204
rect 10022 -2992 10080 -2980
rect 10180 -2204 10238 -2192
rect 10180 -2980 10192 -2204
rect 10226 -2980 10238 -2204
rect 10180 -2992 10238 -2980
rect 10338 -2204 10396 -2192
rect 10338 -2980 10350 -2204
rect 10384 -2980 10396 -2204
rect 10338 -2992 10396 -2980
rect 10496 -2204 10554 -2192
rect 10496 -2980 10508 -2204
rect 10542 -2980 10554 -2204
rect 10496 -2992 10554 -2980
rect 10654 -2204 10712 -2192
rect 10654 -2980 10666 -2204
rect 10700 -2980 10712 -2204
rect 10654 -2992 10712 -2980
rect 10812 -2204 10870 -2192
rect 10812 -2980 10824 -2204
rect 10858 -2980 10870 -2204
rect 10812 -2992 10870 -2980
rect 10970 -2204 11028 -2192
rect 10970 -2980 10982 -2204
rect 11016 -2980 11028 -2204
rect 10970 -2992 11028 -2980
rect 14035 -1997 14165 -1955
rect 14035 -2037 14165 -2027
rect 14035 -2071 14055 -2037
rect 14089 -2071 14165 -2037
rect 14035 -2079 14165 -2071
rect 14035 -2141 14165 -2133
rect 14035 -2175 14055 -2141
rect 14089 -2175 14165 -2141
rect 14035 -2185 14165 -2175
rect 12774 -2206 12874 -2194
rect 12774 -2240 12786 -2206
rect 12862 -2240 12874 -2206
rect 12774 -2252 12874 -2240
rect 12774 -3064 12874 -3052
rect 12774 -3098 12786 -3064
rect 12862 -3098 12874 -3064
rect 12774 -3110 12874 -3098
rect 15539 -1835 15591 -1797
rect 15539 -1869 15547 -1835
rect 15581 -1869 15591 -1835
rect 15539 -1881 15591 -1869
rect 15621 -1809 15675 -1797
rect 15621 -1843 15631 -1809
rect 15665 -1843 15675 -1809
rect 15621 -1881 15675 -1843
rect 15705 -1835 15757 -1797
rect 15705 -1869 15715 -1835
rect 15749 -1869 15757 -1835
rect 15705 -1881 15757 -1869
rect 15825 -1805 15930 -1797
rect 15825 -1839 15837 -1805
rect 15871 -1839 15930 -1805
rect 15825 -1881 15930 -1839
rect 15960 -1811 16025 -1797
rect 15960 -1845 15970 -1811
rect 16004 -1845 16025 -1811
rect 15960 -1869 16025 -1845
rect 16055 -1811 16121 -1797
rect 16055 -1845 16077 -1811
rect 16111 -1845 16121 -1811
rect 16055 -1869 16121 -1845
rect 16151 -1869 16287 -1797
rect 15960 -1881 16010 -1869
rect 16169 -1881 16287 -1869
rect 16317 -1881 16359 -1797
rect 16389 -1809 16491 -1797
rect 16389 -1843 16423 -1809
rect 16457 -1843 16491 -1809
rect 16389 -1881 16491 -1843
rect 14035 -2281 14165 -2215
rect 16441 -1925 16491 -1881
rect 16521 -1805 16590 -1797
rect 16521 -1839 16535 -1805
rect 16569 -1839 16590 -1805
rect 16521 -1869 16590 -1839
rect 16620 -1809 16699 -1797
rect 16620 -1843 16645 -1809
rect 16679 -1843 16699 -1809
rect 16620 -1869 16699 -1843
rect 16729 -1869 16795 -1797
rect 16521 -1925 16575 -1869
rect 16745 -1881 16795 -1869
rect 16825 -1805 16944 -1797
rect 16825 -1839 16857 -1805
rect 16891 -1839 16944 -1805
rect 16825 -1881 16944 -1839
rect 16974 -1881 17035 -1797
rect 17065 -1825 17117 -1797
rect 17065 -1859 17075 -1825
rect 17109 -1859 17117 -1825
rect 17065 -1881 17117 -1859
rect 17171 -1848 17223 -1797
rect 17171 -1882 17179 -1848
rect 17213 -1882 17223 -1848
rect 17171 -1927 17223 -1882
rect 17253 -1813 17305 -1797
rect 17253 -1847 17263 -1813
rect 17297 -1847 17305 -1813
rect 17253 -1881 17305 -1847
rect 17359 -1835 17411 -1797
rect 17359 -1869 17367 -1835
rect 17401 -1869 17411 -1835
rect 17359 -1881 17411 -1869
rect 17441 -1829 17508 -1797
rect 17441 -1863 17464 -1829
rect 17498 -1863 17508 -1829
rect 17441 -1881 17508 -1863
rect 17253 -1915 17263 -1881
rect 17297 -1915 17305 -1881
rect 17253 -1927 17305 -1915
rect 17456 -1927 17508 -1881
rect 17538 -1859 17590 -1797
rect 17538 -1893 17548 -1859
rect 17582 -1893 17590 -1859
rect 17538 -1927 17590 -1893
rect 17747 -1835 17799 -1797
rect 17747 -1869 17755 -1835
rect 17789 -1869 17799 -1835
rect 17747 -1881 17799 -1869
rect 17829 -1809 17883 -1797
rect 17829 -1843 17839 -1809
rect 17873 -1843 17883 -1809
rect 17829 -1881 17883 -1843
rect 17913 -1835 17965 -1797
rect 17913 -1869 17923 -1835
rect 17957 -1869 17965 -1835
rect 17913 -1881 17965 -1869
rect 18033 -1805 18138 -1797
rect 18033 -1839 18045 -1805
rect 18079 -1839 18138 -1805
rect 18033 -1881 18138 -1839
rect 18168 -1811 18233 -1797
rect 18168 -1845 18178 -1811
rect 18212 -1845 18233 -1811
rect 18168 -1869 18233 -1845
rect 18263 -1811 18329 -1797
rect 18263 -1845 18285 -1811
rect 18319 -1845 18329 -1811
rect 18263 -1869 18329 -1845
rect 18359 -1869 18495 -1797
rect 18168 -1881 18218 -1869
rect 18377 -1881 18495 -1869
rect 18525 -1881 18567 -1797
rect 18597 -1809 18699 -1797
rect 18597 -1843 18631 -1809
rect 18665 -1843 18699 -1809
rect 18597 -1881 18699 -1843
rect 18649 -1925 18699 -1881
rect 18729 -1805 18798 -1797
rect 18729 -1839 18743 -1805
rect 18777 -1839 18798 -1805
rect 18729 -1869 18798 -1839
rect 18828 -1809 18907 -1797
rect 18828 -1843 18853 -1809
rect 18887 -1843 18907 -1809
rect 18828 -1869 18907 -1843
rect 18937 -1869 19003 -1797
rect 18729 -1925 18783 -1869
rect 18953 -1881 19003 -1869
rect 19033 -1805 19152 -1797
rect 19033 -1839 19065 -1805
rect 19099 -1839 19152 -1805
rect 19033 -1881 19152 -1839
rect 19182 -1881 19243 -1797
rect 19273 -1825 19325 -1797
rect 19273 -1859 19283 -1825
rect 19317 -1859 19325 -1825
rect 19273 -1881 19325 -1859
rect 19379 -1848 19431 -1797
rect 19379 -1882 19387 -1848
rect 19421 -1882 19431 -1848
rect 19379 -1927 19431 -1882
rect 19461 -1813 19513 -1797
rect 19461 -1847 19471 -1813
rect 19505 -1847 19513 -1813
rect 19461 -1881 19513 -1847
rect 19567 -1835 19619 -1797
rect 19567 -1869 19575 -1835
rect 19609 -1869 19619 -1835
rect 19567 -1881 19619 -1869
rect 19649 -1829 19716 -1797
rect 19649 -1863 19672 -1829
rect 19706 -1863 19716 -1829
rect 19649 -1881 19716 -1863
rect 19461 -1915 19471 -1881
rect 19505 -1915 19513 -1881
rect 19461 -1927 19513 -1915
rect 19664 -1927 19716 -1881
rect 19746 -1859 19798 -1797
rect 19746 -1893 19756 -1859
rect 19790 -1893 19798 -1859
rect 19746 -1927 19798 -1893
rect 19955 -1835 20007 -1797
rect 19955 -1869 19963 -1835
rect 19997 -1869 20007 -1835
rect 19955 -1881 20007 -1869
rect 20037 -1809 20091 -1797
rect 20037 -1843 20047 -1809
rect 20081 -1843 20091 -1809
rect 20037 -1881 20091 -1843
rect 20121 -1835 20173 -1797
rect 20121 -1869 20131 -1835
rect 20165 -1869 20173 -1835
rect 20121 -1881 20173 -1869
rect 20241 -1805 20346 -1797
rect 20241 -1839 20253 -1805
rect 20287 -1839 20346 -1805
rect 20241 -1881 20346 -1839
rect 20376 -1811 20441 -1797
rect 20376 -1845 20386 -1811
rect 20420 -1845 20441 -1811
rect 20376 -1869 20441 -1845
rect 20471 -1811 20537 -1797
rect 20471 -1845 20493 -1811
rect 20527 -1845 20537 -1811
rect 20471 -1869 20537 -1845
rect 20567 -1869 20703 -1797
rect 20376 -1881 20426 -1869
rect 20585 -1881 20703 -1869
rect 20733 -1881 20775 -1797
rect 20805 -1809 20907 -1797
rect 20805 -1843 20839 -1809
rect 20873 -1843 20907 -1809
rect 20805 -1881 20907 -1843
rect 20857 -1925 20907 -1881
rect 20937 -1805 21006 -1797
rect 20937 -1839 20951 -1805
rect 20985 -1839 21006 -1805
rect 20937 -1869 21006 -1839
rect 21036 -1809 21115 -1797
rect 21036 -1843 21061 -1809
rect 21095 -1843 21115 -1809
rect 21036 -1869 21115 -1843
rect 21145 -1869 21211 -1797
rect 20937 -1925 20991 -1869
rect 21161 -1881 21211 -1869
rect 21241 -1805 21360 -1797
rect 21241 -1839 21273 -1805
rect 21307 -1839 21360 -1805
rect 21241 -1881 21360 -1839
rect 21390 -1881 21451 -1797
rect 21481 -1825 21533 -1797
rect 21481 -1859 21491 -1825
rect 21525 -1859 21533 -1825
rect 21481 -1881 21533 -1859
rect 21587 -1848 21639 -1797
rect 21587 -1882 21595 -1848
rect 21629 -1882 21639 -1848
rect 21587 -1927 21639 -1882
rect 21669 -1813 21721 -1797
rect 21669 -1847 21679 -1813
rect 21713 -1847 21721 -1813
rect 21669 -1881 21721 -1847
rect 21775 -1835 21827 -1797
rect 21775 -1869 21783 -1835
rect 21817 -1869 21827 -1835
rect 21775 -1881 21827 -1869
rect 21857 -1829 21924 -1797
rect 21857 -1863 21880 -1829
rect 21914 -1863 21924 -1829
rect 21857 -1881 21924 -1863
rect 21669 -1915 21679 -1881
rect 21713 -1915 21721 -1881
rect 21669 -1927 21721 -1915
rect 21872 -1927 21924 -1881
rect 21954 -1859 22006 -1797
rect 21954 -1893 21964 -1859
rect 21998 -1893 22006 -1859
rect 21954 -1927 22006 -1893
rect 14035 -2321 14165 -2311
rect 14035 -2355 14051 -2321
rect 14085 -2355 14165 -2321
rect 14035 -2374 14165 -2355
rect 14035 -2414 14165 -2404
rect 14035 -2448 14055 -2414
rect 14089 -2448 14165 -2414
rect 14035 -2456 14165 -2448
rect 14035 -2524 14119 -2516
rect 14035 -2558 14060 -2524
rect 14094 -2558 14119 -2524
rect 14035 -2568 14119 -2558
rect 14035 -2617 14119 -2598
rect 14035 -2651 14043 -2617
rect 14077 -2651 14119 -2617
rect 14035 -2671 14119 -2651
rect 14035 -2743 14119 -2701
rect 14035 -2783 14119 -2773
rect 14035 -2817 14055 -2783
rect 14089 -2817 14119 -2783
rect 14035 -2825 14119 -2817
rect 15000 -2732 15053 -2707
rect 15000 -2766 15008 -2732
rect 15042 -2766 15053 -2732
rect 15000 -2791 15053 -2766
rect 15083 -2791 15125 -2707
rect 15155 -2749 15247 -2707
rect 15155 -2783 15179 -2749
rect 15213 -2783 15247 -2749
rect 15155 -2791 15247 -2783
rect 15277 -2745 15330 -2707
rect 15277 -2779 15288 -2745
rect 15322 -2779 15330 -2745
rect 15539 -2719 15591 -2707
rect 15539 -2753 15547 -2719
rect 15581 -2753 15591 -2719
rect 15277 -2791 15330 -2779
rect 15539 -2791 15591 -2753
rect 15621 -2745 15675 -2707
rect 15621 -2779 15631 -2745
rect 15665 -2779 15675 -2745
rect 15621 -2791 15675 -2779
rect 15705 -2719 15757 -2707
rect 15705 -2753 15715 -2719
rect 15749 -2753 15757 -2719
rect 15705 -2791 15757 -2753
rect 15825 -2749 15930 -2707
rect 15825 -2783 15837 -2749
rect 15871 -2783 15930 -2749
rect 15825 -2791 15930 -2783
rect 15960 -2719 16010 -2707
rect 16441 -2707 16491 -2663
rect 16169 -2719 16287 -2707
rect 15960 -2743 16025 -2719
rect 15960 -2777 15970 -2743
rect 16004 -2777 16025 -2743
rect 15960 -2791 16025 -2777
rect 16055 -2743 16121 -2719
rect 16055 -2777 16077 -2743
rect 16111 -2777 16121 -2743
rect 16055 -2791 16121 -2777
rect 16151 -2791 16287 -2719
rect 16317 -2791 16359 -2707
rect 16389 -2745 16491 -2707
rect 16389 -2779 16423 -2745
rect 16457 -2779 16491 -2745
rect 16389 -2791 16491 -2779
rect 16521 -2719 16575 -2663
rect 17171 -2706 17223 -2661
rect 16745 -2719 16795 -2707
rect 16521 -2749 16590 -2719
rect 16521 -2783 16535 -2749
rect 16569 -2783 16590 -2749
rect 16521 -2791 16590 -2783
rect 16620 -2745 16699 -2719
rect 16620 -2779 16645 -2745
rect 16679 -2779 16699 -2745
rect 16620 -2791 16699 -2779
rect 16729 -2791 16795 -2719
rect 16825 -2749 16944 -2707
rect 16825 -2783 16857 -2749
rect 16891 -2783 16944 -2749
rect 16825 -2791 16944 -2783
rect 16974 -2791 17035 -2707
rect 17065 -2729 17117 -2707
rect 17065 -2763 17075 -2729
rect 17109 -2763 17117 -2729
rect 17065 -2791 17117 -2763
rect 17171 -2740 17179 -2706
rect 17213 -2740 17223 -2706
rect 17171 -2791 17223 -2740
rect 17253 -2673 17305 -2661
rect 17253 -2707 17263 -2673
rect 17297 -2707 17305 -2673
rect 17456 -2707 17508 -2661
rect 17253 -2741 17305 -2707
rect 17253 -2775 17263 -2741
rect 17297 -2775 17305 -2741
rect 17253 -2791 17305 -2775
rect 17359 -2719 17411 -2707
rect 17359 -2753 17367 -2719
rect 17401 -2753 17411 -2719
rect 17359 -2791 17411 -2753
rect 17441 -2725 17508 -2707
rect 17441 -2759 17464 -2725
rect 17498 -2759 17508 -2725
rect 17441 -2791 17508 -2759
rect 17538 -2695 17590 -2661
rect 17538 -2729 17548 -2695
rect 17582 -2729 17590 -2695
rect 17538 -2791 17590 -2729
rect 17747 -2719 17799 -2707
rect 17747 -2753 17755 -2719
rect 17789 -2753 17799 -2719
rect 17747 -2791 17799 -2753
rect 17829 -2745 17883 -2707
rect 17829 -2779 17839 -2745
rect 17873 -2779 17883 -2745
rect 17829 -2791 17883 -2779
rect 17913 -2719 17965 -2707
rect 17913 -2753 17923 -2719
rect 17957 -2753 17965 -2719
rect 17913 -2791 17965 -2753
rect 18033 -2749 18138 -2707
rect 18033 -2783 18045 -2749
rect 18079 -2783 18138 -2749
rect 18033 -2791 18138 -2783
rect 18168 -2719 18218 -2707
rect 18649 -2707 18699 -2663
rect 18377 -2719 18495 -2707
rect 18168 -2743 18233 -2719
rect 18168 -2777 18178 -2743
rect 18212 -2777 18233 -2743
rect 18168 -2791 18233 -2777
rect 18263 -2743 18329 -2719
rect 18263 -2777 18285 -2743
rect 18319 -2777 18329 -2743
rect 18263 -2791 18329 -2777
rect 18359 -2791 18495 -2719
rect 18525 -2791 18567 -2707
rect 18597 -2745 18699 -2707
rect 18597 -2779 18631 -2745
rect 18665 -2779 18699 -2745
rect 18597 -2791 18699 -2779
rect 18729 -2719 18783 -2663
rect 19379 -2706 19431 -2661
rect 18953 -2719 19003 -2707
rect 18729 -2749 18798 -2719
rect 18729 -2783 18743 -2749
rect 18777 -2783 18798 -2749
rect 18729 -2791 18798 -2783
rect 18828 -2745 18907 -2719
rect 18828 -2779 18853 -2745
rect 18887 -2779 18907 -2745
rect 18828 -2791 18907 -2779
rect 18937 -2791 19003 -2719
rect 19033 -2749 19152 -2707
rect 19033 -2783 19065 -2749
rect 19099 -2783 19152 -2749
rect 19033 -2791 19152 -2783
rect 19182 -2791 19243 -2707
rect 19273 -2729 19325 -2707
rect 19273 -2763 19283 -2729
rect 19317 -2763 19325 -2729
rect 19273 -2791 19325 -2763
rect 19379 -2740 19387 -2706
rect 19421 -2740 19431 -2706
rect 19379 -2791 19431 -2740
rect 19461 -2673 19513 -2661
rect 19461 -2707 19471 -2673
rect 19505 -2707 19513 -2673
rect 19664 -2707 19716 -2661
rect 19461 -2741 19513 -2707
rect 19461 -2775 19471 -2741
rect 19505 -2775 19513 -2741
rect 19461 -2791 19513 -2775
rect 19567 -2719 19619 -2707
rect 19567 -2753 19575 -2719
rect 19609 -2753 19619 -2719
rect 19567 -2791 19619 -2753
rect 19649 -2725 19716 -2707
rect 19649 -2759 19672 -2725
rect 19706 -2759 19716 -2725
rect 19649 -2791 19716 -2759
rect 19746 -2695 19798 -2661
rect 19746 -2729 19756 -2695
rect 19790 -2729 19798 -2695
rect 19746 -2791 19798 -2729
rect 19955 -2719 20007 -2707
rect 19955 -2753 19963 -2719
rect 19997 -2753 20007 -2719
rect 19955 -2791 20007 -2753
rect 20037 -2745 20091 -2707
rect 20037 -2779 20047 -2745
rect 20081 -2779 20091 -2745
rect 20037 -2791 20091 -2779
rect 20121 -2719 20173 -2707
rect 20121 -2753 20131 -2719
rect 20165 -2753 20173 -2719
rect 20121 -2791 20173 -2753
rect 20241 -2749 20346 -2707
rect 20241 -2783 20253 -2749
rect 20287 -2783 20346 -2749
rect 20241 -2791 20346 -2783
rect 20376 -2719 20426 -2707
rect 20857 -2707 20907 -2663
rect 20585 -2719 20703 -2707
rect 20376 -2743 20441 -2719
rect 20376 -2777 20386 -2743
rect 20420 -2777 20441 -2743
rect 20376 -2791 20441 -2777
rect 20471 -2743 20537 -2719
rect 20471 -2777 20493 -2743
rect 20527 -2777 20537 -2743
rect 20471 -2791 20537 -2777
rect 20567 -2791 20703 -2719
rect 20733 -2791 20775 -2707
rect 20805 -2745 20907 -2707
rect 20805 -2779 20839 -2745
rect 20873 -2779 20907 -2745
rect 20805 -2791 20907 -2779
rect 20937 -2719 20991 -2663
rect 21587 -2706 21639 -2661
rect 21161 -2719 21211 -2707
rect 20937 -2749 21006 -2719
rect 20937 -2783 20951 -2749
rect 20985 -2783 21006 -2749
rect 20937 -2791 21006 -2783
rect 21036 -2745 21115 -2719
rect 21036 -2779 21061 -2745
rect 21095 -2779 21115 -2745
rect 21036 -2791 21115 -2779
rect 21145 -2791 21211 -2719
rect 21241 -2749 21360 -2707
rect 21241 -2783 21273 -2749
rect 21307 -2783 21360 -2749
rect 21241 -2791 21360 -2783
rect 21390 -2791 21451 -2707
rect 21481 -2729 21533 -2707
rect 21481 -2763 21491 -2729
rect 21525 -2763 21533 -2729
rect 21481 -2791 21533 -2763
rect 21587 -2740 21595 -2706
rect 21629 -2740 21639 -2706
rect 21587 -2791 21639 -2740
rect 21669 -2673 21721 -2661
rect 21669 -2707 21679 -2673
rect 21713 -2707 21721 -2673
rect 21872 -2707 21924 -2661
rect 21669 -2741 21721 -2707
rect 21669 -2775 21679 -2741
rect 21713 -2775 21721 -2741
rect 21669 -2791 21721 -2775
rect 21775 -2719 21827 -2707
rect 21775 -2753 21783 -2719
rect 21817 -2753 21827 -2719
rect 21775 -2791 21827 -2753
rect 21857 -2725 21924 -2707
rect 21857 -2759 21880 -2725
rect 21914 -2759 21924 -2725
rect 21857 -2791 21924 -2759
rect 21954 -2695 22006 -2661
rect 21954 -2729 21964 -2695
rect 21998 -2729 22006 -2695
rect 21954 -2791 22006 -2729
rect 15098 -3178 15156 -3166
rect 15098 -3254 15110 -3178
rect 15144 -3254 15156 -3178
rect 15098 -3266 15156 -3254
rect 15956 -3178 16014 -3166
rect 15956 -3254 15968 -3178
rect 16002 -3254 16014 -3178
rect 15956 -3266 16014 -3254
rect 16202 -4750 16260 -4738
rect 16202 -5526 16214 -4750
rect 16248 -5526 16260 -4750
rect 16202 -5538 16260 -5526
rect 16660 -4750 16718 -4738
rect 16660 -5526 16672 -4750
rect 16706 -5526 16718 -4750
rect 16660 -5538 16718 -5526
rect 17118 -4750 17176 -4738
rect 17118 -5526 17130 -4750
rect 17164 -5526 17176 -4750
rect 17118 -5538 17176 -5526
rect 17576 -4750 17634 -4738
rect 17576 -5526 17588 -4750
rect 17622 -5526 17634 -4750
rect 17576 -5538 17634 -5526
rect 18034 -4750 18092 -4738
rect 18034 -5526 18046 -4750
rect 18080 -5526 18092 -4750
rect 18034 -5538 18092 -5526
rect 18890 -5546 18948 -5534
rect 18890 -5622 18902 -5546
rect 18936 -5622 18948 -5546
rect 18890 -5634 18948 -5622
rect 20548 -5546 20606 -5534
rect 20548 -5622 20560 -5546
rect 20594 -5622 20606 -5546
rect 20548 -5634 20606 -5622
rect 21354 -5418 21412 -5406
rect 21354 -5494 21366 -5418
rect 21400 -5494 21412 -5418
rect 21354 -5506 21412 -5494
rect 21612 -5418 21670 -5406
rect 21612 -5494 21624 -5418
rect 21658 -5494 21670 -5418
rect 21612 -5506 21670 -5494
rect 21870 -5418 21928 -5406
rect 21870 -5494 21882 -5418
rect 21916 -5494 21928 -5418
rect 21870 -5506 21928 -5494
rect 21354 -5628 21412 -5616
rect 21354 -5704 21366 -5628
rect 21400 -5704 21412 -5628
rect 21354 -5716 21412 -5704
rect 21612 -5628 21670 -5616
rect 21612 -5704 21624 -5628
rect 21658 -5704 21670 -5628
rect 21612 -5716 21670 -5704
rect 21870 -5628 21928 -5616
rect 21870 -5704 21882 -5628
rect 21916 -5704 21928 -5628
rect 21870 -5716 21928 -5704
rect 23434 -5402 23584 -5390
rect 23434 -5436 23446 -5402
rect 23572 -5436 23584 -5402
rect 23434 -5448 23584 -5436
rect 23434 -5660 23584 -5648
rect 23434 -5694 23446 -5660
rect 23572 -5694 23584 -5660
rect 23434 -5706 23584 -5694
rect 9208 -7700 9308 -7688
rect 9208 -7734 9220 -7700
rect 9296 -7734 9308 -7700
rect 9208 -7746 9308 -7734
rect 9208 -9358 9308 -9346
rect 9208 -9392 9220 -9358
rect 9296 -9392 9308 -9358
rect 9208 -9404 9308 -9392
<< pdiff >>
rect 3289 -1359 3447 -1351
rect 3289 -1393 3325 -1359
rect 3359 -1393 3393 -1359
rect 3427 -1393 3447 -1359
rect 3289 -1403 3447 -1393
rect 4883 -1359 5041 -1351
rect 4883 -1393 4903 -1359
rect 4937 -1393 4971 -1359
rect 5005 -1393 5041 -1359
rect 4883 -1403 5041 -1393
rect 3289 -1445 3447 -1433
rect 3289 -1479 3325 -1445
rect 3359 -1479 3393 -1445
rect 3427 -1479 3447 -1445
rect 3289 -1491 3447 -1479
rect 4883 -1445 5041 -1433
rect 4883 -1479 4903 -1445
rect 4937 -1479 4971 -1445
rect 5005 -1479 5041 -1445
rect 4883 -1491 5041 -1479
rect 3289 -1531 3447 -1521
rect 3289 -1565 3312 -1531
rect 3346 -1565 3393 -1531
rect 3427 -1565 3447 -1531
rect 3289 -1573 3447 -1565
rect 4883 -1531 5041 -1521
rect 4883 -1565 4903 -1531
rect 4937 -1565 4984 -1531
rect 5018 -1565 5041 -1531
rect 4883 -1573 5041 -1565
rect 14285 -1785 14485 -1777
rect 14285 -1819 14301 -1785
rect 14335 -1819 14431 -1785
rect 14465 -1819 14485 -1785
rect 14285 -1829 14485 -1819
rect 14285 -1869 14485 -1859
rect 3354 -2135 3412 -2123
rect 3354 -2311 3366 -2135
rect 3400 -2311 3412 -2135
rect 3354 -2323 3412 -2311
rect 3612 -2135 3670 -2123
rect 3612 -2311 3624 -2135
rect 3658 -2311 3670 -2135
rect 3612 -2323 3670 -2311
rect 4666 -2135 4724 -2123
rect 4666 -2311 4678 -2135
rect 4712 -2311 4724 -2135
rect 4666 -2323 4724 -2311
rect 4924 -2135 4982 -2123
rect 4924 -2311 4936 -2135
rect 4970 -2311 4982 -2135
rect 4924 -2323 4982 -2311
rect 14285 -1903 14363 -1869
rect 14397 -1903 14431 -1869
rect 14465 -1903 14485 -1869
rect 14285 -1913 14485 -1903
rect 14285 -1953 14485 -1943
rect 7464 -2199 7522 -2187
rect 7464 -2975 7476 -2199
rect 7510 -2975 7522 -2199
rect 7464 -2987 7522 -2975
rect 7622 -2199 7680 -2187
rect 7622 -2975 7634 -2199
rect 7668 -2975 7680 -2199
rect 7622 -2987 7680 -2975
rect 7780 -2199 7838 -2187
rect 7780 -2975 7792 -2199
rect 7826 -2975 7838 -2199
rect 7780 -2987 7838 -2975
rect 7938 -2199 7996 -2187
rect 7938 -2975 7950 -2199
rect 7984 -2975 7996 -2199
rect 7938 -2987 7996 -2975
rect 8096 -2199 8154 -2187
rect 8096 -2975 8108 -2199
rect 8142 -2975 8154 -2199
rect 8096 -2987 8154 -2975
rect 8254 -2199 8312 -2187
rect 8254 -2975 8266 -2199
rect 8300 -2975 8312 -2199
rect 8254 -2987 8312 -2975
rect 8412 -2199 8470 -2187
rect 8412 -2975 8424 -2199
rect 8458 -2975 8470 -2199
rect 8412 -2987 8470 -2975
rect 8570 -2199 8628 -2187
rect 8570 -2975 8582 -2199
rect 8616 -2975 8628 -2199
rect 8570 -2987 8628 -2975
rect 8728 -2199 8786 -2187
rect 8728 -2975 8740 -2199
rect 8774 -2975 8786 -2199
rect 8728 -2987 8786 -2975
rect 8886 -2199 8944 -2187
rect 8886 -2975 8898 -2199
rect 8932 -2975 8944 -2199
rect 8886 -2987 8944 -2975
rect 9044 -2199 9102 -2187
rect 9044 -2975 9056 -2199
rect 9090 -2975 9102 -2199
rect 9044 -2987 9102 -2975
rect 14285 -1987 14363 -1953
rect 14397 -1987 14485 -1953
rect 14285 -1997 14485 -1987
rect 14285 -2037 14485 -2027
rect 14285 -2071 14439 -2037
rect 14473 -2071 14485 -2037
rect 14285 -2079 14485 -2071
rect 14285 -2141 14485 -2133
rect 14285 -2175 14431 -2141
rect 14465 -2175 14485 -2141
rect 14285 -2185 14485 -2175
rect 15197 -2133 15295 -2119
rect 15197 -2163 15248 -2133
rect 14285 -2230 14485 -2215
rect 15000 -2201 15053 -2163
rect 14285 -2264 14361 -2230
rect 14395 -2264 14431 -2230
rect 14465 -2264 14485 -2230
rect 15000 -2235 15008 -2201
rect 15042 -2235 15053 -2201
rect 15000 -2247 15053 -2235
rect 15083 -2193 15141 -2163
rect 15083 -2227 15096 -2193
rect 15130 -2227 15141 -2193
rect 15083 -2247 15141 -2227
rect 15171 -2167 15248 -2163
rect 15282 -2167 15295 -2133
rect 15171 -2201 15295 -2167
rect 15171 -2235 15182 -2201
rect 15216 -2235 15250 -2201
rect 15284 -2235 15295 -2201
rect 15171 -2247 15295 -2235
rect 15325 -2133 15378 -2119
rect 15325 -2167 15336 -2133
rect 15370 -2167 15378 -2133
rect 15325 -2201 15378 -2167
rect 15325 -2235 15336 -2201
rect 15370 -2235 15378 -2201
rect 15539 -2125 15591 -2113
rect 15539 -2159 15547 -2125
rect 15581 -2159 15591 -2125
rect 15539 -2193 15591 -2159
rect 15539 -2227 15547 -2193
rect 15581 -2227 15591 -2193
rect 15325 -2247 15378 -2235
rect 15539 -2241 15591 -2227
rect 15621 -2177 15675 -2113
rect 15621 -2211 15631 -2177
rect 15665 -2211 15675 -2177
rect 15621 -2241 15675 -2211
rect 15705 -2125 15757 -2113
rect 15705 -2159 15715 -2125
rect 15749 -2159 15757 -2125
rect 15705 -2193 15757 -2159
rect 15705 -2227 15715 -2193
rect 15749 -2227 15757 -2193
rect 15705 -2241 15757 -2227
rect 15890 -2201 15942 -2163
rect 15890 -2235 15898 -2201
rect 15932 -2235 15942 -2201
rect 14285 -2281 14485 -2264
rect 15890 -2247 15942 -2235
rect 15972 -2193 16034 -2163
rect 15972 -2227 15982 -2193
rect 16016 -2227 16034 -2193
rect 15972 -2247 16034 -2227
rect 16064 -2199 16133 -2163
rect 16064 -2233 16075 -2199
rect 16109 -2233 16133 -2199
rect 16064 -2247 16133 -2233
rect 16163 -2175 16273 -2163
rect 16163 -2209 16229 -2175
rect 16263 -2209 16273 -2175
rect 16163 -2247 16273 -2209
rect 16303 -2191 16370 -2163
rect 16303 -2225 16326 -2191
rect 16360 -2225 16370 -2191
rect 16303 -2247 16370 -2225
rect 16400 -2175 16452 -2163
rect 16400 -2209 16410 -2175
rect 16444 -2209 16452 -2175
rect 16400 -2247 16452 -2209
rect 16515 -2201 16567 -2079
rect 16515 -2235 16523 -2201
rect 16557 -2235 16567 -2201
rect 16515 -2247 16567 -2235
rect 16597 -2163 16651 -2079
rect 17142 -2163 17192 -2047
rect 16597 -2193 16666 -2163
rect 16597 -2227 16611 -2193
rect 16645 -2227 16666 -2193
rect 16597 -2247 16666 -2227
rect 16696 -2200 16752 -2163
rect 16696 -2234 16708 -2200
rect 16742 -2234 16752 -2200
rect 16696 -2247 16752 -2234
rect 16782 -2247 16836 -2163
rect 16866 -2201 16944 -2163
rect 16866 -2235 16900 -2201
rect 16934 -2235 16944 -2201
rect 16866 -2247 16944 -2235
rect 16974 -2175 17028 -2163
rect 16974 -2209 16984 -2175
rect 17018 -2209 17028 -2175
rect 16974 -2247 17028 -2209
rect 17058 -2201 17192 -2163
rect 17058 -2235 17070 -2201
rect 17104 -2235 17148 -2201
rect 17182 -2235 17192 -2201
rect 17058 -2247 17192 -2235
rect 17222 -2057 17278 -2047
rect 17222 -2091 17232 -2057
rect 17266 -2091 17278 -2057
rect 17222 -2125 17278 -2091
rect 17456 -2065 17508 -2047
rect 17456 -2099 17464 -2065
rect 17498 -2099 17508 -2065
rect 17456 -2119 17508 -2099
rect 17222 -2159 17232 -2125
rect 17266 -2159 17278 -2125
rect 17222 -2193 17278 -2159
rect 17222 -2227 17232 -2193
rect 17266 -2227 17278 -2193
rect 17222 -2247 17278 -2227
rect 17359 -2133 17411 -2119
rect 17359 -2167 17367 -2133
rect 17401 -2167 17411 -2133
rect 17359 -2201 17411 -2167
rect 17359 -2235 17367 -2201
rect 17401 -2235 17411 -2201
rect 17359 -2247 17411 -2235
rect 17441 -2133 17508 -2119
rect 17441 -2167 17464 -2133
rect 17498 -2167 17508 -2133
rect 17441 -2201 17508 -2167
rect 17441 -2235 17464 -2201
rect 17498 -2235 17508 -2201
rect 17441 -2247 17508 -2235
rect 17538 -2097 17590 -2047
rect 17538 -2131 17548 -2097
rect 17582 -2131 17590 -2097
rect 17538 -2165 17590 -2131
rect 17538 -2199 17548 -2165
rect 17582 -2199 17590 -2165
rect 17538 -2247 17590 -2199
rect 17747 -2125 17799 -2113
rect 17747 -2159 17755 -2125
rect 17789 -2159 17799 -2125
rect 17747 -2193 17799 -2159
rect 17747 -2227 17755 -2193
rect 17789 -2227 17799 -2193
rect 17747 -2241 17799 -2227
rect 17829 -2177 17883 -2113
rect 17829 -2211 17839 -2177
rect 17873 -2211 17883 -2177
rect 17829 -2241 17883 -2211
rect 17913 -2125 17965 -2113
rect 17913 -2159 17923 -2125
rect 17957 -2159 17965 -2125
rect 17913 -2193 17965 -2159
rect 17913 -2227 17923 -2193
rect 17957 -2227 17965 -2193
rect 17913 -2241 17965 -2227
rect 18098 -2201 18150 -2163
rect 18098 -2235 18106 -2201
rect 18140 -2235 18150 -2201
rect 18098 -2247 18150 -2235
rect 18180 -2193 18242 -2163
rect 18180 -2227 18190 -2193
rect 18224 -2227 18242 -2193
rect 18180 -2247 18242 -2227
rect 18272 -2199 18341 -2163
rect 18272 -2233 18283 -2199
rect 18317 -2233 18341 -2199
rect 18272 -2247 18341 -2233
rect 18371 -2175 18481 -2163
rect 18371 -2209 18437 -2175
rect 18471 -2209 18481 -2175
rect 18371 -2247 18481 -2209
rect 18511 -2191 18578 -2163
rect 18511 -2225 18534 -2191
rect 18568 -2225 18578 -2191
rect 18511 -2247 18578 -2225
rect 18608 -2175 18660 -2163
rect 18608 -2209 18618 -2175
rect 18652 -2209 18660 -2175
rect 18608 -2247 18660 -2209
rect 18723 -2201 18775 -2079
rect 18723 -2235 18731 -2201
rect 18765 -2235 18775 -2201
rect 18723 -2247 18775 -2235
rect 18805 -2163 18859 -2079
rect 19350 -2163 19400 -2047
rect 18805 -2193 18874 -2163
rect 18805 -2227 18819 -2193
rect 18853 -2227 18874 -2193
rect 18805 -2247 18874 -2227
rect 18904 -2200 18960 -2163
rect 18904 -2234 18916 -2200
rect 18950 -2234 18960 -2200
rect 18904 -2247 18960 -2234
rect 18990 -2247 19044 -2163
rect 19074 -2201 19152 -2163
rect 19074 -2235 19108 -2201
rect 19142 -2235 19152 -2201
rect 19074 -2247 19152 -2235
rect 19182 -2175 19236 -2163
rect 19182 -2209 19192 -2175
rect 19226 -2209 19236 -2175
rect 19182 -2247 19236 -2209
rect 19266 -2201 19400 -2163
rect 19266 -2235 19278 -2201
rect 19312 -2235 19356 -2201
rect 19390 -2235 19400 -2201
rect 19266 -2247 19400 -2235
rect 19430 -2057 19486 -2047
rect 19430 -2091 19440 -2057
rect 19474 -2091 19486 -2057
rect 19430 -2125 19486 -2091
rect 19664 -2065 19716 -2047
rect 19664 -2099 19672 -2065
rect 19706 -2099 19716 -2065
rect 19664 -2119 19716 -2099
rect 19430 -2159 19440 -2125
rect 19474 -2159 19486 -2125
rect 19430 -2193 19486 -2159
rect 19430 -2227 19440 -2193
rect 19474 -2227 19486 -2193
rect 19430 -2247 19486 -2227
rect 19567 -2133 19619 -2119
rect 19567 -2167 19575 -2133
rect 19609 -2167 19619 -2133
rect 19567 -2201 19619 -2167
rect 19567 -2235 19575 -2201
rect 19609 -2235 19619 -2201
rect 19567 -2247 19619 -2235
rect 19649 -2133 19716 -2119
rect 19649 -2167 19672 -2133
rect 19706 -2167 19716 -2133
rect 19649 -2201 19716 -2167
rect 19649 -2235 19672 -2201
rect 19706 -2235 19716 -2201
rect 19649 -2247 19716 -2235
rect 19746 -2097 19798 -2047
rect 19746 -2131 19756 -2097
rect 19790 -2131 19798 -2097
rect 19746 -2165 19798 -2131
rect 19746 -2199 19756 -2165
rect 19790 -2199 19798 -2165
rect 19746 -2247 19798 -2199
rect 19955 -2125 20007 -2113
rect 19955 -2159 19963 -2125
rect 19997 -2159 20007 -2125
rect 19955 -2193 20007 -2159
rect 19955 -2227 19963 -2193
rect 19997 -2227 20007 -2193
rect 19955 -2241 20007 -2227
rect 20037 -2177 20091 -2113
rect 20037 -2211 20047 -2177
rect 20081 -2211 20091 -2177
rect 20037 -2241 20091 -2211
rect 20121 -2125 20173 -2113
rect 20121 -2159 20131 -2125
rect 20165 -2159 20173 -2125
rect 20121 -2193 20173 -2159
rect 20121 -2227 20131 -2193
rect 20165 -2227 20173 -2193
rect 20121 -2241 20173 -2227
rect 20306 -2201 20358 -2163
rect 20306 -2235 20314 -2201
rect 20348 -2235 20358 -2201
rect 20306 -2247 20358 -2235
rect 20388 -2193 20450 -2163
rect 20388 -2227 20398 -2193
rect 20432 -2227 20450 -2193
rect 20388 -2247 20450 -2227
rect 20480 -2199 20549 -2163
rect 20480 -2233 20491 -2199
rect 20525 -2233 20549 -2199
rect 20480 -2247 20549 -2233
rect 20579 -2175 20689 -2163
rect 20579 -2209 20645 -2175
rect 20679 -2209 20689 -2175
rect 20579 -2247 20689 -2209
rect 20719 -2191 20786 -2163
rect 20719 -2225 20742 -2191
rect 20776 -2225 20786 -2191
rect 20719 -2247 20786 -2225
rect 20816 -2175 20868 -2163
rect 20816 -2209 20826 -2175
rect 20860 -2209 20868 -2175
rect 20816 -2247 20868 -2209
rect 20931 -2201 20983 -2079
rect 20931 -2235 20939 -2201
rect 20973 -2235 20983 -2201
rect 20931 -2247 20983 -2235
rect 21013 -2163 21067 -2079
rect 21558 -2163 21608 -2047
rect 21013 -2193 21082 -2163
rect 21013 -2227 21027 -2193
rect 21061 -2227 21082 -2193
rect 21013 -2247 21082 -2227
rect 21112 -2200 21168 -2163
rect 21112 -2234 21124 -2200
rect 21158 -2234 21168 -2200
rect 21112 -2247 21168 -2234
rect 21198 -2247 21252 -2163
rect 21282 -2201 21360 -2163
rect 21282 -2235 21316 -2201
rect 21350 -2235 21360 -2201
rect 21282 -2247 21360 -2235
rect 21390 -2175 21444 -2163
rect 21390 -2209 21400 -2175
rect 21434 -2209 21444 -2175
rect 21390 -2247 21444 -2209
rect 21474 -2201 21608 -2163
rect 21474 -2235 21486 -2201
rect 21520 -2235 21564 -2201
rect 21598 -2235 21608 -2201
rect 21474 -2247 21608 -2235
rect 21638 -2057 21694 -2047
rect 21638 -2091 21648 -2057
rect 21682 -2091 21694 -2057
rect 21638 -2125 21694 -2091
rect 21872 -2065 21924 -2047
rect 21872 -2099 21880 -2065
rect 21914 -2099 21924 -2065
rect 21872 -2119 21924 -2099
rect 21638 -2159 21648 -2125
rect 21682 -2159 21694 -2125
rect 21638 -2193 21694 -2159
rect 21638 -2227 21648 -2193
rect 21682 -2227 21694 -2193
rect 21638 -2247 21694 -2227
rect 21775 -2133 21827 -2119
rect 21775 -2167 21783 -2133
rect 21817 -2167 21827 -2133
rect 21775 -2201 21827 -2167
rect 21775 -2235 21783 -2201
rect 21817 -2235 21827 -2201
rect 21775 -2247 21827 -2235
rect 21857 -2133 21924 -2119
rect 21857 -2167 21880 -2133
rect 21914 -2167 21924 -2133
rect 21857 -2201 21924 -2167
rect 21857 -2235 21880 -2201
rect 21914 -2235 21924 -2201
rect 21857 -2247 21924 -2235
rect 21954 -2097 22006 -2047
rect 21954 -2131 21964 -2097
rect 21998 -2131 22006 -2097
rect 21954 -2165 22006 -2131
rect 21954 -2199 21964 -2165
rect 21998 -2199 22006 -2165
rect 21954 -2247 22006 -2199
rect 14285 -2330 14485 -2311
rect 14285 -2364 14363 -2330
rect 14397 -2364 14431 -2330
rect 14465 -2364 14485 -2330
rect 15000 -2353 15053 -2341
rect 14285 -2374 14485 -2364
rect 14285 -2414 14485 -2404
rect 14285 -2448 14363 -2414
rect 14397 -2448 14431 -2414
rect 14465 -2448 14485 -2414
rect 14285 -2456 14485 -2448
rect 15000 -2387 15008 -2353
rect 15042 -2387 15053 -2353
rect 15000 -2425 15053 -2387
rect 15083 -2361 15141 -2341
rect 15083 -2395 15096 -2361
rect 15130 -2395 15141 -2361
rect 15083 -2425 15141 -2395
rect 15171 -2353 15295 -2341
rect 15171 -2387 15182 -2353
rect 15216 -2387 15250 -2353
rect 15284 -2387 15295 -2353
rect 15171 -2421 15295 -2387
rect 15171 -2425 15248 -2421
rect 14401 -2524 14485 -2516
rect 14401 -2558 14426 -2524
rect 14460 -2558 14485 -2524
rect 15197 -2455 15248 -2425
rect 15282 -2455 15295 -2421
rect 15197 -2469 15295 -2455
rect 15325 -2353 15378 -2341
rect 15325 -2387 15336 -2353
rect 15370 -2387 15378 -2353
rect 15325 -2421 15378 -2387
rect 15325 -2455 15336 -2421
rect 15370 -2455 15378 -2421
rect 15325 -2469 15378 -2455
rect 14401 -2568 14485 -2558
rect 14401 -2613 14485 -2598
rect 14357 -2618 14485 -2613
rect 14357 -2652 14443 -2618
rect 14477 -2652 14485 -2618
rect 14357 -2671 14485 -2652
rect 14357 -2743 14485 -2701
rect 15539 -2361 15591 -2347
rect 15539 -2395 15547 -2361
rect 15581 -2395 15591 -2361
rect 15539 -2429 15591 -2395
rect 15539 -2463 15547 -2429
rect 15581 -2463 15591 -2429
rect 15539 -2475 15591 -2463
rect 15621 -2377 15675 -2347
rect 15621 -2411 15631 -2377
rect 15665 -2411 15675 -2377
rect 15621 -2475 15675 -2411
rect 15705 -2361 15757 -2347
rect 15705 -2395 15715 -2361
rect 15749 -2395 15757 -2361
rect 15705 -2429 15757 -2395
rect 15890 -2353 15942 -2341
rect 15890 -2387 15898 -2353
rect 15932 -2387 15942 -2353
rect 15890 -2425 15942 -2387
rect 15972 -2361 16034 -2341
rect 15972 -2395 15982 -2361
rect 16016 -2395 16034 -2361
rect 15972 -2425 16034 -2395
rect 16064 -2355 16133 -2341
rect 16064 -2389 16075 -2355
rect 16109 -2389 16133 -2355
rect 16064 -2425 16133 -2389
rect 16163 -2379 16273 -2341
rect 16163 -2413 16229 -2379
rect 16263 -2413 16273 -2379
rect 16163 -2425 16273 -2413
rect 16303 -2363 16370 -2341
rect 16303 -2397 16326 -2363
rect 16360 -2397 16370 -2363
rect 16303 -2425 16370 -2397
rect 16400 -2379 16452 -2341
rect 16400 -2413 16410 -2379
rect 16444 -2413 16452 -2379
rect 16400 -2425 16452 -2413
rect 16515 -2353 16567 -2341
rect 16515 -2387 16523 -2353
rect 16557 -2387 16567 -2353
rect 15705 -2463 15715 -2429
rect 15749 -2463 15757 -2429
rect 15705 -2475 15757 -2463
rect 14357 -2783 14485 -2773
rect 14357 -2817 14431 -2783
rect 14465 -2817 14485 -2783
rect 16515 -2509 16567 -2387
rect 16597 -2361 16666 -2341
rect 16597 -2395 16611 -2361
rect 16645 -2395 16666 -2361
rect 16597 -2425 16666 -2395
rect 16696 -2354 16752 -2341
rect 16696 -2388 16708 -2354
rect 16742 -2388 16752 -2354
rect 16696 -2425 16752 -2388
rect 16782 -2425 16836 -2341
rect 16866 -2353 16944 -2341
rect 16866 -2387 16900 -2353
rect 16934 -2387 16944 -2353
rect 16866 -2425 16944 -2387
rect 16974 -2379 17028 -2341
rect 16974 -2413 16984 -2379
rect 17018 -2413 17028 -2379
rect 16974 -2425 17028 -2413
rect 17058 -2353 17192 -2341
rect 17058 -2387 17070 -2353
rect 17104 -2387 17148 -2353
rect 17182 -2387 17192 -2353
rect 17058 -2425 17192 -2387
rect 16597 -2509 16651 -2425
rect 17142 -2541 17192 -2425
rect 17222 -2361 17278 -2341
rect 17222 -2395 17232 -2361
rect 17266 -2395 17278 -2361
rect 17222 -2429 17278 -2395
rect 17222 -2463 17232 -2429
rect 17266 -2463 17278 -2429
rect 17222 -2497 17278 -2463
rect 17359 -2353 17411 -2341
rect 17359 -2387 17367 -2353
rect 17401 -2387 17411 -2353
rect 17359 -2421 17411 -2387
rect 17359 -2455 17367 -2421
rect 17401 -2455 17411 -2421
rect 17359 -2469 17411 -2455
rect 17441 -2353 17508 -2341
rect 17441 -2387 17464 -2353
rect 17498 -2387 17508 -2353
rect 17441 -2421 17508 -2387
rect 17441 -2455 17464 -2421
rect 17498 -2455 17508 -2421
rect 17441 -2469 17508 -2455
rect 17222 -2531 17232 -2497
rect 17266 -2531 17278 -2497
rect 17222 -2541 17278 -2531
rect 17456 -2489 17508 -2469
rect 17456 -2523 17464 -2489
rect 17498 -2523 17508 -2489
rect 17456 -2541 17508 -2523
rect 17538 -2389 17590 -2341
rect 17538 -2423 17548 -2389
rect 17582 -2423 17590 -2389
rect 17538 -2457 17590 -2423
rect 17538 -2491 17548 -2457
rect 17582 -2491 17590 -2457
rect 17538 -2541 17590 -2491
rect 17747 -2361 17799 -2347
rect 17747 -2395 17755 -2361
rect 17789 -2395 17799 -2361
rect 17747 -2429 17799 -2395
rect 17747 -2463 17755 -2429
rect 17789 -2463 17799 -2429
rect 17747 -2475 17799 -2463
rect 17829 -2377 17883 -2347
rect 17829 -2411 17839 -2377
rect 17873 -2411 17883 -2377
rect 17829 -2475 17883 -2411
rect 17913 -2361 17965 -2347
rect 17913 -2395 17923 -2361
rect 17957 -2395 17965 -2361
rect 17913 -2429 17965 -2395
rect 18098 -2353 18150 -2341
rect 18098 -2387 18106 -2353
rect 18140 -2387 18150 -2353
rect 18098 -2425 18150 -2387
rect 18180 -2361 18242 -2341
rect 18180 -2395 18190 -2361
rect 18224 -2395 18242 -2361
rect 18180 -2425 18242 -2395
rect 18272 -2355 18341 -2341
rect 18272 -2389 18283 -2355
rect 18317 -2389 18341 -2355
rect 18272 -2425 18341 -2389
rect 18371 -2379 18481 -2341
rect 18371 -2413 18437 -2379
rect 18471 -2413 18481 -2379
rect 18371 -2425 18481 -2413
rect 18511 -2363 18578 -2341
rect 18511 -2397 18534 -2363
rect 18568 -2397 18578 -2363
rect 18511 -2425 18578 -2397
rect 18608 -2379 18660 -2341
rect 18608 -2413 18618 -2379
rect 18652 -2413 18660 -2379
rect 18608 -2425 18660 -2413
rect 18723 -2353 18775 -2341
rect 18723 -2387 18731 -2353
rect 18765 -2387 18775 -2353
rect 17913 -2463 17923 -2429
rect 17957 -2463 17965 -2429
rect 17913 -2475 17965 -2463
rect 18723 -2509 18775 -2387
rect 18805 -2361 18874 -2341
rect 18805 -2395 18819 -2361
rect 18853 -2395 18874 -2361
rect 18805 -2425 18874 -2395
rect 18904 -2354 18960 -2341
rect 18904 -2388 18916 -2354
rect 18950 -2388 18960 -2354
rect 18904 -2425 18960 -2388
rect 18990 -2425 19044 -2341
rect 19074 -2353 19152 -2341
rect 19074 -2387 19108 -2353
rect 19142 -2387 19152 -2353
rect 19074 -2425 19152 -2387
rect 19182 -2379 19236 -2341
rect 19182 -2413 19192 -2379
rect 19226 -2413 19236 -2379
rect 19182 -2425 19236 -2413
rect 19266 -2353 19400 -2341
rect 19266 -2387 19278 -2353
rect 19312 -2387 19356 -2353
rect 19390 -2387 19400 -2353
rect 19266 -2425 19400 -2387
rect 18805 -2509 18859 -2425
rect 19350 -2541 19400 -2425
rect 19430 -2361 19486 -2341
rect 19430 -2395 19440 -2361
rect 19474 -2395 19486 -2361
rect 19430 -2429 19486 -2395
rect 19430 -2463 19440 -2429
rect 19474 -2463 19486 -2429
rect 19430 -2497 19486 -2463
rect 19567 -2353 19619 -2341
rect 19567 -2387 19575 -2353
rect 19609 -2387 19619 -2353
rect 19567 -2421 19619 -2387
rect 19567 -2455 19575 -2421
rect 19609 -2455 19619 -2421
rect 19567 -2469 19619 -2455
rect 19649 -2353 19716 -2341
rect 19649 -2387 19672 -2353
rect 19706 -2387 19716 -2353
rect 19649 -2421 19716 -2387
rect 19649 -2455 19672 -2421
rect 19706 -2455 19716 -2421
rect 19649 -2469 19716 -2455
rect 19430 -2531 19440 -2497
rect 19474 -2531 19486 -2497
rect 19430 -2541 19486 -2531
rect 19664 -2489 19716 -2469
rect 19664 -2523 19672 -2489
rect 19706 -2523 19716 -2489
rect 19664 -2541 19716 -2523
rect 19746 -2389 19798 -2341
rect 19746 -2423 19756 -2389
rect 19790 -2423 19798 -2389
rect 19746 -2457 19798 -2423
rect 19746 -2491 19756 -2457
rect 19790 -2491 19798 -2457
rect 19746 -2541 19798 -2491
rect 19955 -2361 20007 -2347
rect 19955 -2395 19963 -2361
rect 19997 -2395 20007 -2361
rect 19955 -2429 20007 -2395
rect 19955 -2463 19963 -2429
rect 19997 -2463 20007 -2429
rect 19955 -2475 20007 -2463
rect 20037 -2377 20091 -2347
rect 20037 -2411 20047 -2377
rect 20081 -2411 20091 -2377
rect 20037 -2475 20091 -2411
rect 20121 -2361 20173 -2347
rect 20121 -2395 20131 -2361
rect 20165 -2395 20173 -2361
rect 20121 -2429 20173 -2395
rect 20306 -2353 20358 -2341
rect 20306 -2387 20314 -2353
rect 20348 -2387 20358 -2353
rect 20306 -2425 20358 -2387
rect 20388 -2361 20450 -2341
rect 20388 -2395 20398 -2361
rect 20432 -2395 20450 -2361
rect 20388 -2425 20450 -2395
rect 20480 -2355 20549 -2341
rect 20480 -2389 20491 -2355
rect 20525 -2389 20549 -2355
rect 20480 -2425 20549 -2389
rect 20579 -2379 20689 -2341
rect 20579 -2413 20645 -2379
rect 20679 -2413 20689 -2379
rect 20579 -2425 20689 -2413
rect 20719 -2363 20786 -2341
rect 20719 -2397 20742 -2363
rect 20776 -2397 20786 -2363
rect 20719 -2425 20786 -2397
rect 20816 -2379 20868 -2341
rect 20816 -2413 20826 -2379
rect 20860 -2413 20868 -2379
rect 20816 -2425 20868 -2413
rect 20931 -2353 20983 -2341
rect 20931 -2387 20939 -2353
rect 20973 -2387 20983 -2353
rect 20121 -2463 20131 -2429
rect 20165 -2463 20173 -2429
rect 20121 -2475 20173 -2463
rect 20931 -2509 20983 -2387
rect 21013 -2361 21082 -2341
rect 21013 -2395 21027 -2361
rect 21061 -2395 21082 -2361
rect 21013 -2425 21082 -2395
rect 21112 -2354 21168 -2341
rect 21112 -2388 21124 -2354
rect 21158 -2388 21168 -2354
rect 21112 -2425 21168 -2388
rect 21198 -2425 21252 -2341
rect 21282 -2353 21360 -2341
rect 21282 -2387 21316 -2353
rect 21350 -2387 21360 -2353
rect 21282 -2425 21360 -2387
rect 21390 -2379 21444 -2341
rect 21390 -2413 21400 -2379
rect 21434 -2413 21444 -2379
rect 21390 -2425 21444 -2413
rect 21474 -2353 21608 -2341
rect 21474 -2387 21486 -2353
rect 21520 -2387 21564 -2353
rect 21598 -2387 21608 -2353
rect 21474 -2425 21608 -2387
rect 21013 -2509 21067 -2425
rect 21558 -2541 21608 -2425
rect 21638 -2361 21694 -2341
rect 21638 -2395 21648 -2361
rect 21682 -2395 21694 -2361
rect 21638 -2429 21694 -2395
rect 21638 -2463 21648 -2429
rect 21682 -2463 21694 -2429
rect 21638 -2497 21694 -2463
rect 21775 -2353 21827 -2341
rect 21775 -2387 21783 -2353
rect 21817 -2387 21827 -2353
rect 21775 -2421 21827 -2387
rect 21775 -2455 21783 -2421
rect 21817 -2455 21827 -2421
rect 21775 -2469 21827 -2455
rect 21857 -2353 21924 -2341
rect 21857 -2387 21880 -2353
rect 21914 -2387 21924 -2353
rect 21857 -2421 21924 -2387
rect 21857 -2455 21880 -2421
rect 21914 -2455 21924 -2421
rect 21857 -2469 21924 -2455
rect 21638 -2531 21648 -2497
rect 21682 -2531 21694 -2497
rect 21638 -2541 21694 -2531
rect 21872 -2489 21924 -2469
rect 21872 -2523 21880 -2489
rect 21914 -2523 21924 -2489
rect 21872 -2541 21924 -2523
rect 21954 -2389 22006 -2341
rect 21954 -2423 21964 -2389
rect 21998 -2423 22006 -2389
rect 21954 -2457 22006 -2423
rect 21954 -2491 21964 -2457
rect 21998 -2491 22006 -2457
rect 21954 -2541 22006 -2491
rect 14357 -2825 14485 -2817
rect 10624 -6001 10682 -5989
rect 10624 -6377 10636 -6001
rect 10670 -6377 10682 -6001
rect 10624 -6389 10682 -6377
rect 11082 -6001 11140 -5989
rect 11082 -6377 11094 -6001
rect 11128 -6377 11140 -6001
rect 11082 -6389 11140 -6377
rect 11196 -6001 11254 -5989
rect 11196 -6377 11208 -6001
rect 11242 -6377 11254 -6001
rect 11196 -6389 11254 -6377
rect 11654 -6001 11712 -5989
rect 11654 -6377 11666 -6001
rect 11700 -6377 11712 -6001
rect 11654 -6389 11712 -6377
rect 11768 -6001 11826 -5989
rect 11768 -6377 11780 -6001
rect 11814 -6377 11826 -6001
rect 11768 -6389 11826 -6377
rect 12226 -6001 12284 -5989
rect 12226 -6377 12238 -6001
rect 12272 -6377 12284 -6001
rect 12226 -6389 12284 -6377
rect 12340 -6001 12398 -5989
rect 12340 -6377 12352 -6001
rect 12386 -6377 12398 -6001
rect 12340 -6389 12398 -6377
rect 12798 -6001 12856 -5989
rect 12798 -6377 12810 -6001
rect 12844 -6377 12856 -6001
rect 12798 -6389 12856 -6377
rect 12912 -6001 12970 -5989
rect 12912 -6377 12924 -6001
rect 12958 -6377 12970 -6001
rect 12912 -6389 12970 -6377
rect 13370 -6001 13428 -5989
rect 13370 -6377 13382 -6001
rect 13416 -6377 13428 -6001
rect 13370 -6389 13428 -6377
rect 13484 -6001 13542 -5989
rect 13484 -6377 13496 -6001
rect 13530 -6377 13542 -6001
rect 13484 -6389 13542 -6377
rect 13942 -6001 14000 -5989
rect 13942 -6377 13954 -6001
rect 13988 -6377 14000 -6001
rect 13942 -6389 14000 -6377
rect 14056 -6001 14114 -5989
rect 14056 -6377 14068 -6001
rect 14102 -6377 14114 -6001
rect 14056 -6389 14114 -6377
rect 14514 -6001 14572 -5989
rect 14514 -6377 14526 -6001
rect 14560 -6377 14572 -6001
rect 14514 -6389 14572 -6377
rect 14628 -6001 14686 -5989
rect 14628 -6377 14640 -6001
rect 14674 -6377 14686 -6001
rect 14628 -6389 14686 -6377
rect 15086 -6001 15144 -5989
rect 15086 -6377 15098 -6001
rect 15132 -6377 15144 -6001
rect 15086 -6389 15144 -6377
rect 10624 -6529 10682 -6517
rect 10624 -6905 10636 -6529
rect 10670 -6905 10682 -6529
rect 10624 -6917 10682 -6905
rect 11082 -6529 11140 -6517
rect 11082 -6905 11094 -6529
rect 11128 -6905 11140 -6529
rect 11082 -6917 11140 -6905
rect 11196 -6529 11254 -6517
rect 11196 -6905 11208 -6529
rect 11242 -6905 11254 -6529
rect 11196 -6917 11254 -6905
rect 11654 -6529 11712 -6517
rect 11654 -6905 11666 -6529
rect 11700 -6905 11712 -6529
rect 11654 -6917 11712 -6905
rect 11768 -6529 11826 -6517
rect 11768 -6905 11780 -6529
rect 11814 -6905 11826 -6529
rect 11768 -6917 11826 -6905
rect 12226 -6529 12284 -6517
rect 12226 -6905 12238 -6529
rect 12272 -6905 12284 -6529
rect 12226 -6917 12284 -6905
rect 12340 -6529 12398 -6517
rect 12340 -6905 12352 -6529
rect 12386 -6905 12398 -6529
rect 12340 -6917 12398 -6905
rect 12798 -6529 12856 -6517
rect 12798 -6905 12810 -6529
rect 12844 -6905 12856 -6529
rect 12798 -6917 12856 -6905
rect 12912 -6529 12970 -6517
rect 12912 -6905 12924 -6529
rect 12958 -6905 12970 -6529
rect 12912 -6917 12970 -6905
rect 13370 -6529 13428 -6517
rect 13370 -6905 13382 -6529
rect 13416 -6905 13428 -6529
rect 13370 -6917 13428 -6905
rect 13484 -6529 13542 -6517
rect 13484 -6905 13496 -6529
rect 13530 -6905 13542 -6529
rect 13484 -6917 13542 -6905
rect 13942 -6529 14000 -6517
rect 13942 -6905 13954 -6529
rect 13988 -6905 14000 -6529
rect 13942 -6917 14000 -6905
rect 14056 -6529 14114 -6517
rect 14056 -6905 14068 -6529
rect 14102 -6905 14114 -6529
rect 14056 -6917 14114 -6905
rect 14514 -6529 14572 -6517
rect 14514 -6905 14526 -6529
rect 14560 -6905 14572 -6529
rect 14514 -6917 14572 -6905
rect 14628 -6529 14686 -6517
rect 14628 -6905 14640 -6529
rect 14674 -6905 14686 -6529
rect 14628 -6917 14686 -6905
rect 15086 -6529 15144 -6517
rect 15086 -6905 15098 -6529
rect 15132 -6905 15144 -6529
rect 15086 -6917 15144 -6905
rect 18870 -6559 18928 -6547
rect 18870 -6635 18882 -6559
rect 18916 -6635 18928 -6559
rect 18870 -6647 18928 -6635
rect 20528 -6559 20586 -6547
rect 20528 -6635 20540 -6559
rect 20574 -6635 20586 -6559
rect 20528 -6647 20586 -6635
rect 21354 -6423 21412 -6411
rect 21354 -6499 21366 -6423
rect 21400 -6499 21412 -6423
rect 21354 -6511 21412 -6499
rect 21612 -6423 21670 -6411
rect 21612 -6499 21624 -6423
rect 21658 -6499 21670 -6423
rect 21612 -6511 21670 -6499
rect 21870 -6423 21928 -6411
rect 21870 -6499 21882 -6423
rect 21916 -6499 21928 -6423
rect 21870 -6511 21928 -6499
rect 21354 -6651 21412 -6639
rect 21354 -6727 21366 -6651
rect 21400 -6727 21412 -6651
rect 21354 -6739 21412 -6727
rect 21612 -6651 21670 -6639
rect 21612 -6727 21624 -6651
rect 21658 -6727 21670 -6651
rect 21612 -6739 21670 -6727
rect 21870 -6651 21928 -6639
rect 21870 -6727 21882 -6651
rect 21916 -6727 21928 -6651
rect 21870 -6739 21928 -6727
rect 23131 -6404 23931 -6392
rect 23131 -6438 23143 -6404
rect 23919 -6438 23931 -6404
rect 23131 -6450 23931 -6438
rect 23131 -6662 23931 -6650
rect 23131 -6696 23143 -6662
rect 23919 -6696 23931 -6662
rect 23131 -6708 23931 -6696
rect 9797 -7434 9897 -7422
rect 9797 -7468 9809 -7434
rect 9885 -7468 9897 -7434
rect 9797 -7480 9897 -7468
rect 9797 -9092 9897 -9080
rect 9797 -9126 9809 -9092
rect 9885 -9126 9897 -9092
rect 9797 -9138 9897 -9126
<< mvndiff >>
rect 2670 -4138 2728 -4126
rect 2670 -4714 2682 -4138
rect 2716 -4714 2728 -4138
rect 2670 -4726 2728 -4714
rect 2828 -4138 2886 -4126
rect 2828 -4714 2840 -4138
rect 2874 -4714 2886 -4138
rect 2828 -4726 2886 -4714
rect 2986 -4138 3044 -4126
rect 2986 -4714 2998 -4138
rect 3032 -4714 3044 -4138
rect 2986 -4726 3044 -4714
rect 3376 -4138 3434 -4126
rect 3376 -4714 3388 -4138
rect 3422 -4714 3434 -4138
rect 3376 -4726 3434 -4714
rect 3534 -4138 3592 -4126
rect 3534 -4714 3546 -4138
rect 3580 -4714 3592 -4138
rect 3534 -4726 3592 -4714
rect 3692 -4138 3750 -4126
rect 3692 -4714 3704 -4138
rect 3738 -4714 3750 -4138
rect 3692 -4726 3750 -4714
rect 4586 -4138 4644 -4126
rect 4586 -4714 4598 -4138
rect 4632 -4714 4644 -4138
rect 4586 -4726 4644 -4714
rect 4744 -4138 4802 -4126
rect 4744 -4714 4756 -4138
rect 4790 -4714 4802 -4138
rect 4744 -4726 4802 -4714
rect 4902 -4138 4960 -4126
rect 4902 -4714 4914 -4138
rect 4948 -4714 4960 -4138
rect 4902 -4726 4960 -4714
rect 5292 -4138 5350 -4126
rect 5292 -4714 5304 -4138
rect 5338 -4714 5350 -4138
rect 5292 -4726 5350 -4714
rect 5450 -4138 5508 -4126
rect 5450 -4714 5462 -4138
rect 5496 -4714 5508 -4138
rect 5450 -4726 5508 -4714
rect 5608 -4138 5666 -4126
rect 5608 -4714 5620 -4138
rect 5654 -4714 5666 -4138
rect 5608 -4726 5666 -4714
rect 2439 -7265 2497 -7253
rect 2439 -8041 2451 -7265
rect 2485 -8041 2497 -7265
rect 2439 -8053 2497 -8041
rect 2597 -7265 2655 -7253
rect 2597 -8041 2609 -7265
rect 2643 -8041 2655 -7265
rect 2597 -8053 2655 -8041
rect 2755 -7265 2813 -7253
rect 2755 -8041 2767 -7265
rect 2801 -8041 2813 -7265
rect 2755 -8053 2813 -8041
rect 2913 -7265 2971 -7253
rect 2913 -8041 2925 -7265
rect 2959 -8041 2971 -7265
rect 2913 -8053 2971 -8041
rect 3071 -7265 3129 -7253
rect 3071 -8041 3083 -7265
rect 3117 -8041 3129 -7265
rect 3071 -8053 3129 -8041
rect 3229 -7265 3287 -7253
rect 3229 -8041 3241 -7265
rect 3275 -8041 3287 -7265
rect 3229 -8053 3287 -8041
rect 10600 -4970 10658 -4958
rect 10600 -5346 10612 -4970
rect 10646 -5346 10658 -4970
rect 10600 -5358 10658 -5346
rect 11058 -4970 11116 -4958
rect 11058 -5346 11070 -4970
rect 11104 -5346 11116 -4970
rect 11058 -5358 11116 -5346
rect 11178 -4970 11236 -4958
rect 11178 -5346 11190 -4970
rect 11224 -5346 11236 -4970
rect 11178 -5358 11236 -5346
rect 11636 -4970 11694 -4958
rect 11636 -5346 11648 -4970
rect 11682 -5346 11694 -4970
rect 11636 -5358 11694 -5346
rect 11756 -4970 11814 -4958
rect 11756 -5346 11768 -4970
rect 11802 -5346 11814 -4970
rect 11756 -5358 11814 -5346
rect 12214 -4970 12272 -4958
rect 12214 -5346 12226 -4970
rect 12260 -5346 12272 -4970
rect 12214 -5358 12272 -5346
rect 12334 -4970 12392 -4958
rect 12334 -5346 12346 -4970
rect 12380 -5346 12392 -4970
rect 12334 -5358 12392 -5346
rect 12792 -4970 12850 -4958
rect 12792 -5346 12804 -4970
rect 12838 -5346 12850 -4970
rect 12792 -5358 12850 -5346
rect 12912 -4970 12970 -4958
rect 12912 -5346 12924 -4970
rect 12958 -5346 12970 -4970
rect 12912 -5358 12970 -5346
rect 13370 -4970 13428 -4958
rect 13370 -5346 13382 -4970
rect 13416 -5346 13428 -4970
rect 13370 -5358 13428 -5346
rect 13490 -4970 13548 -4958
rect 13490 -5346 13502 -4970
rect 13536 -5346 13548 -4970
rect 13490 -5358 13548 -5346
rect 13948 -4970 14006 -4958
rect 13948 -5346 13960 -4970
rect 13994 -5346 14006 -4970
rect 13948 -5358 14006 -5346
rect 14068 -4970 14126 -4958
rect 14068 -5346 14080 -4970
rect 14114 -5346 14126 -4970
rect 14068 -5358 14126 -5346
rect 14526 -4970 14584 -4958
rect 14526 -5346 14538 -4970
rect 14572 -5346 14584 -4970
rect 14526 -5358 14584 -5346
rect 14646 -4970 14704 -4958
rect 14646 -5346 14658 -4970
rect 14692 -5346 14704 -4970
rect 14646 -5358 14704 -5346
rect 15104 -4970 15162 -4958
rect 15104 -5346 15116 -4970
rect 15150 -5346 15162 -4970
rect 15104 -5358 15162 -5346
rect 7268 -12262 7326 -12250
rect 7268 -12438 7280 -12262
rect 7314 -12438 7326 -12262
rect 7268 -12450 7326 -12438
rect 7526 -12262 7584 -12250
rect 7526 -12438 7538 -12262
rect 7572 -12438 7584 -12262
rect 7526 -12450 7584 -12438
rect 8210 -12322 8268 -12310
rect 8210 -12382 8222 -12322
rect 8256 -12382 8268 -12322
rect 8210 -12394 8268 -12382
rect 9868 -12322 9926 -12310
rect 9868 -12382 9880 -12322
rect 9914 -12382 9926 -12322
rect 9868 -12394 9926 -12382
rect 11526 -12322 11584 -12310
rect 11526 -12382 11538 -12322
rect 11572 -12382 11584 -12322
rect 11526 -12394 11584 -12382
rect 13184 -12322 13242 -12310
rect 13184 -12382 13196 -12322
rect 13230 -12382 13242 -12322
rect 13184 -12394 13242 -12382
rect 19998 -12700 20798 -12688
rect 19998 -12734 20010 -12700
rect 20786 -12734 20798 -12700
rect 19998 -12746 20798 -12734
rect 20908 -12700 21708 -12688
rect 20908 -12734 20920 -12700
rect 21696 -12734 21708 -12700
rect 20908 -12746 21708 -12734
rect 19998 -13158 20798 -13146
rect 19998 -13192 20010 -13158
rect 20786 -13192 20798 -13158
rect 19998 -13204 20798 -13192
rect 20908 -13158 21708 -13146
rect 20908 -13192 20920 -13158
rect 21696 -13192 21708 -13158
rect 20908 -13204 21708 -13192
rect 19998 -13278 20798 -13266
rect 19998 -13312 20010 -13278
rect 20786 -13312 20798 -13278
rect 19998 -13324 20798 -13312
rect 20908 -13278 21708 -13266
rect 20908 -13312 20920 -13278
rect 21696 -13312 21708 -13278
rect 20908 -13324 21708 -13312
rect 19998 -13736 20798 -13724
rect 19998 -13770 20010 -13736
rect 20786 -13770 20798 -13736
rect 19998 -13782 20798 -13770
rect 20908 -13736 21708 -13724
rect 20908 -13770 20920 -13736
rect 21696 -13770 21708 -13736
rect 20908 -13782 21708 -13770
rect 19998 -13856 20798 -13844
rect 19998 -13890 20010 -13856
rect 20786 -13890 20798 -13856
rect 19998 -13902 20798 -13890
rect 20908 -13856 21708 -13844
rect 20908 -13890 20920 -13856
rect 21696 -13890 21708 -13856
rect 20908 -13902 21708 -13890
rect 19998 -14314 20798 -14302
rect 19998 -14348 20010 -14314
rect 20786 -14348 20798 -14314
rect 19998 -14360 20798 -14348
rect 20908 -14314 21708 -14302
rect 20908 -14348 20920 -14314
rect 21696 -14348 21708 -14314
rect 20908 -14360 21708 -14348
rect 19998 -14434 20798 -14422
rect 19998 -14468 20010 -14434
rect 20786 -14468 20798 -14434
rect 19998 -14480 20798 -14468
rect 20908 -14434 21708 -14422
rect 20908 -14468 20920 -14434
rect 21696 -14468 21708 -14434
rect 20908 -14480 21708 -14468
rect 19998 -14892 20798 -14880
rect 19998 -14926 20010 -14892
rect 20786 -14926 20798 -14892
rect 19998 -14938 20798 -14926
rect 20908 -14892 21708 -14880
rect 20908 -14926 20920 -14892
rect 21696 -14926 21708 -14892
rect 20908 -14938 21708 -14926
rect 19998 -15012 20798 -15000
rect 19998 -15046 20010 -15012
rect 20786 -15046 20798 -15012
rect 19998 -15058 20798 -15046
rect 20908 -15012 21708 -15000
rect 20908 -15046 20920 -15012
rect 21696 -15046 21708 -15012
rect 20908 -15058 21708 -15046
rect 19998 -15470 20798 -15458
rect 19998 -15504 20010 -15470
rect 20786 -15504 20798 -15470
rect 19998 -15516 20798 -15504
rect 20908 -15470 21708 -15458
rect 20908 -15504 20920 -15470
rect 21696 -15504 21708 -15470
rect 20908 -15516 21708 -15504
rect 20464 -16044 21264 -16032
rect 20464 -16078 20476 -16044
rect 21252 -16078 21264 -16044
rect 20464 -16090 21264 -16078
rect 20464 -16202 21264 -16190
rect 20464 -16236 20476 -16202
rect 21252 -16236 21264 -16202
rect 20464 -16248 21264 -16236
rect 20464 -16360 21264 -16348
rect 20464 -16394 20476 -16360
rect 21252 -16394 21264 -16360
rect 20464 -16406 21264 -16394
rect 20464 -16518 21264 -16506
rect 20464 -16552 20476 -16518
rect 21252 -16552 21264 -16518
rect 20464 -16564 21264 -16552
rect 20464 -16676 21264 -16664
rect 20464 -16710 20476 -16676
rect 21252 -16710 21264 -16676
rect 20464 -16722 21264 -16710
rect 20464 -16834 21264 -16822
rect 20464 -16868 20476 -16834
rect 21252 -16868 21264 -16834
rect 20464 -16880 21264 -16868
rect 20464 -16992 21264 -16980
rect 20464 -17026 20476 -16992
rect 21252 -17026 21264 -16992
rect 20464 -17038 21264 -17026
rect 20464 -17150 21264 -17138
rect 20464 -17184 20476 -17150
rect 21252 -17184 21264 -17150
rect 20464 -17196 21264 -17184
rect 20464 -17308 21264 -17296
rect 20464 -17342 20476 -17308
rect 21252 -17342 21264 -17308
rect 20464 -17354 21264 -17342
rect 20464 -17466 21264 -17454
rect 20464 -17500 20476 -17466
rect 21252 -17500 21264 -17466
rect 20464 -17512 21264 -17500
rect 20464 -17624 21264 -17612
rect 20464 -17658 20476 -17624
rect 21252 -17658 21264 -17624
rect 20464 -17670 21264 -17658
rect 20464 -17782 21264 -17770
rect 20464 -17816 20476 -17782
rect 21252 -17816 21264 -17782
rect 20464 -17828 21264 -17816
rect 20464 -17940 21264 -17928
rect 20464 -17974 20476 -17940
rect 21252 -17974 21264 -17940
rect 20464 -17986 21264 -17974
<< mvpdiff >>
rect 11422 -2181 11480 -2169
rect 11422 -2957 11434 -2181
rect 11468 -2957 11480 -2181
rect 11422 -2969 11480 -2957
rect 11580 -2181 11638 -2169
rect 11580 -2957 11592 -2181
rect 11626 -2957 11638 -2181
rect 11580 -2969 11638 -2957
rect 2752 -5441 2810 -5429
rect 2752 -5617 2764 -5441
rect 2798 -5617 2810 -5441
rect 2752 -5629 2810 -5617
rect 3610 -5441 3668 -5429
rect 3610 -5617 3622 -5441
rect 3656 -5617 3668 -5441
rect 3610 -5629 3668 -5617
rect 2752 -6045 2810 -6033
rect 2752 -6221 2764 -6045
rect 2798 -6221 2810 -6045
rect 2752 -6233 2810 -6221
rect 3610 -6045 3668 -6033
rect 3610 -6221 3622 -6045
rect 3656 -6221 3668 -6045
rect 3610 -6233 3668 -6221
rect 4668 -5441 4726 -5429
rect 4668 -5617 4680 -5441
rect 4714 -5617 4726 -5441
rect 4668 -5629 4726 -5617
rect 5526 -5441 5584 -5429
rect 5526 -5617 5538 -5441
rect 5572 -5617 5584 -5441
rect 5526 -5629 5584 -5617
rect 4668 -6045 4726 -6033
rect 4668 -6221 4680 -6045
rect 4714 -6221 4726 -6045
rect 4668 -6233 4726 -6221
rect 5526 -6045 5584 -6033
rect 5526 -6221 5538 -6045
rect 5572 -6221 5584 -6045
rect 5526 -6233 5584 -6221
rect 3814 -7267 3872 -7255
rect 3814 -8043 3826 -7267
rect 3860 -8043 3872 -7267
rect 3814 -8055 3872 -8043
rect 3972 -7267 4030 -7255
rect 3972 -8043 3984 -7267
rect 4018 -8043 4030 -7267
rect 3972 -8055 4030 -8043
rect 4130 -7267 4188 -7255
rect 4130 -8043 4142 -7267
rect 4176 -8043 4188 -7267
rect 4130 -8055 4188 -8043
rect 4288 -7267 4346 -7255
rect 4288 -8043 4300 -7267
rect 4334 -8043 4346 -7267
rect 4288 -8055 4346 -8043
rect 4446 -7267 4504 -7255
rect 4446 -8043 4458 -7267
rect 4492 -8043 4504 -7267
rect 4446 -8055 4504 -8043
rect 4604 -7267 4662 -7255
rect 4604 -8043 4616 -7267
rect 4650 -8043 4662 -7267
rect 4604 -8055 4662 -8043
rect 16202 -6109 16260 -6097
rect 16202 -6885 16214 -6109
rect 16248 -6885 16260 -6109
rect 16202 -6897 16260 -6885
rect 16660 -6109 16718 -6097
rect 16660 -6885 16672 -6109
rect 16706 -6885 16718 -6109
rect 16660 -6897 16718 -6885
rect 17118 -6109 17176 -6097
rect 17118 -6885 17130 -6109
rect 17164 -6885 17176 -6109
rect 17118 -6897 17176 -6885
rect 17576 -6109 17634 -6097
rect 17576 -6885 17588 -6109
rect 17622 -6885 17634 -6109
rect 17576 -6897 17634 -6885
rect 18034 -6109 18092 -6097
rect 18034 -6885 18046 -6109
rect 18080 -6885 18092 -6109
rect 18034 -6897 18092 -6885
rect 22601 -12708 23401 -12696
rect 22601 -12742 22613 -12708
rect 23389 -12742 23401 -12708
rect 22601 -12754 23401 -12742
rect 23529 -12708 24329 -12696
rect 23529 -12742 23541 -12708
rect 24317 -12742 24329 -12708
rect 23529 -12754 24329 -12742
rect 22601 -13166 23401 -13154
rect 22601 -13200 22613 -13166
rect 23389 -13200 23401 -13166
rect 22601 -13212 23401 -13200
rect 23529 -13166 24329 -13154
rect 23529 -13200 23541 -13166
rect 24317 -13200 24329 -13166
rect 23529 -13212 24329 -13200
rect 22601 -13286 23401 -13274
rect 22601 -13320 22613 -13286
rect 23389 -13320 23401 -13286
rect 22601 -13332 23401 -13320
rect 23529 -13286 24329 -13274
rect 23529 -13320 23541 -13286
rect 24317 -13320 24329 -13286
rect 23529 -13332 24329 -13320
rect 22601 -13744 23401 -13732
rect 22601 -13778 22613 -13744
rect 23389 -13778 23401 -13744
rect 22601 -13790 23401 -13778
rect 23529 -13744 24329 -13732
rect 23529 -13778 23541 -13744
rect 24317 -13778 24329 -13744
rect 23529 -13790 24329 -13778
rect 22601 -13864 23401 -13852
rect 22601 -13898 22613 -13864
rect 23389 -13898 23401 -13864
rect 22601 -13910 23401 -13898
rect 23529 -13864 24329 -13852
rect 23529 -13898 23541 -13864
rect 24317 -13898 24329 -13864
rect 23529 -13910 24329 -13898
rect 22601 -14322 23401 -14310
rect 22601 -14356 22613 -14322
rect 23389 -14356 23401 -14322
rect 22601 -14368 23401 -14356
rect 23529 -14322 24329 -14310
rect 23529 -14356 23541 -14322
rect 24317 -14356 24329 -14322
rect 23529 -14368 24329 -14356
rect 22601 -14442 23401 -14430
rect 22601 -14476 22613 -14442
rect 23389 -14476 23401 -14442
rect 22601 -14488 23401 -14476
rect 23529 -14442 24329 -14430
rect 23529 -14476 23541 -14442
rect 24317 -14476 24329 -14442
rect 23529 -14488 24329 -14476
rect 22601 -14900 23401 -14888
rect 22601 -14934 22613 -14900
rect 23389 -14934 23401 -14900
rect 22601 -14946 23401 -14934
rect 23529 -14900 24329 -14888
rect 23529 -14934 23541 -14900
rect 24317 -14934 24329 -14900
rect 23529 -14946 24329 -14934
rect 22601 -15020 23401 -15008
rect 22601 -15054 22613 -15020
rect 23389 -15054 23401 -15020
rect 22601 -15066 23401 -15054
rect 23529 -15020 24329 -15008
rect 23529 -15054 23541 -15020
rect 24317 -15054 24329 -15020
rect 23529 -15066 24329 -15054
rect 22601 -15478 23401 -15466
rect 22601 -15512 22613 -15478
rect 23389 -15512 23401 -15478
rect 22601 -15524 23401 -15512
rect 23529 -15478 24329 -15466
rect 23529 -15512 23541 -15478
rect 24317 -15512 24329 -15478
rect 23529 -15524 24329 -15512
rect 22601 -15598 23401 -15586
rect 22601 -15632 22613 -15598
rect 23389 -15632 23401 -15598
rect 22601 -15644 23401 -15632
rect 23529 -15598 24329 -15586
rect 23529 -15632 23541 -15598
rect 24317 -15632 24329 -15598
rect 23529 -15644 24329 -15632
rect 22601 -16056 23401 -16044
rect 22601 -16090 22613 -16056
rect 23389 -16090 23401 -16056
rect 22601 -16102 23401 -16090
rect 23529 -16056 24329 -16044
rect 23529 -16090 23541 -16056
rect 24317 -16090 24329 -16056
rect 23529 -16102 24329 -16090
rect 22601 -16176 23401 -16164
rect 22601 -16210 22613 -16176
rect 23389 -16210 23401 -16176
rect 22601 -16222 23401 -16210
rect 23529 -16176 24329 -16164
rect 23529 -16210 23541 -16176
rect 24317 -16210 24329 -16176
rect 23529 -16222 24329 -16210
rect 22601 -16634 23401 -16622
rect 22601 -16668 22613 -16634
rect 23389 -16668 23401 -16634
rect 22601 -16680 23401 -16668
rect 23529 -16634 24329 -16622
rect 23529 -16668 23541 -16634
rect 24317 -16668 24329 -16634
rect 23529 -16680 24329 -16668
rect 22601 -16754 23401 -16742
rect 22601 -16788 22613 -16754
rect 23389 -16788 23401 -16754
rect 22601 -16800 23401 -16788
rect 23529 -16754 24329 -16742
rect 23529 -16788 23541 -16754
rect 24317 -16788 24329 -16754
rect 23529 -16800 24329 -16788
rect 22601 -17212 23401 -17200
rect 22601 -17246 22613 -17212
rect 23389 -17246 23401 -17212
rect 22601 -17258 23401 -17246
rect 23529 -17212 24329 -17200
rect 23529 -17246 23541 -17212
rect 24317 -17246 24329 -17212
rect 23529 -17258 24329 -17246
rect 22601 -17332 23401 -17320
rect 22601 -17366 22613 -17332
rect 23389 -17366 23401 -17332
rect 22601 -17378 23401 -17366
rect 23529 -17332 24329 -17320
rect 23529 -17366 23541 -17332
rect 24317 -17366 24329 -17332
rect 23529 -17378 24329 -17366
rect 22601 -17790 23401 -17778
rect 22601 -17824 22613 -17790
rect 23389 -17824 23401 -17790
rect 22601 -17836 23401 -17824
rect 23529 -17790 24329 -17778
rect 23529 -17824 23541 -17790
rect 24317 -17824 24329 -17790
rect 23529 -17836 24329 -17824
<< ndiffc >>
rect 3022 -1393 3056 -1359
rect 5274 -1393 5308 -1359
rect 3009 -1479 3043 -1445
rect 5287 -1479 5321 -1445
rect 3039 -1565 3073 -1531
rect 5257 -1565 5291 -1531
rect 14083 -1819 14117 -1785
rect 14059 -1903 14093 -1869
rect 2766 -2310 2800 -2134
rect 3024 -2310 3058 -2134
rect 15008 -1856 15042 -1822
rect 15179 -1839 15213 -1805
rect 15288 -1843 15322 -1809
rect 5278 -2310 5312 -2134
rect 5536 -2310 5570 -2134
rect 9402 -2980 9436 -2204
rect 9560 -2980 9594 -2204
rect 9718 -2980 9752 -2204
rect 9876 -2980 9910 -2204
rect 10034 -2980 10068 -2204
rect 10192 -2980 10226 -2204
rect 10350 -2980 10384 -2204
rect 10508 -2980 10542 -2204
rect 10666 -2980 10700 -2204
rect 10824 -2980 10858 -2204
rect 10982 -2980 11016 -2204
rect 14055 -2071 14089 -2037
rect 14055 -2175 14089 -2141
rect 12786 -2240 12862 -2206
rect 12786 -3098 12862 -3064
rect 15547 -1869 15581 -1835
rect 15631 -1843 15665 -1809
rect 15715 -1869 15749 -1835
rect 15837 -1839 15871 -1805
rect 15970 -1845 16004 -1811
rect 16077 -1845 16111 -1811
rect 16423 -1843 16457 -1809
rect 16535 -1839 16569 -1805
rect 16645 -1843 16679 -1809
rect 16857 -1839 16891 -1805
rect 17075 -1859 17109 -1825
rect 17179 -1882 17213 -1848
rect 17263 -1847 17297 -1813
rect 17367 -1869 17401 -1835
rect 17464 -1863 17498 -1829
rect 17263 -1915 17297 -1881
rect 17548 -1893 17582 -1859
rect 17755 -1869 17789 -1835
rect 17839 -1843 17873 -1809
rect 17923 -1869 17957 -1835
rect 18045 -1839 18079 -1805
rect 18178 -1845 18212 -1811
rect 18285 -1845 18319 -1811
rect 18631 -1843 18665 -1809
rect 18743 -1839 18777 -1805
rect 18853 -1843 18887 -1809
rect 19065 -1839 19099 -1805
rect 19283 -1859 19317 -1825
rect 19387 -1882 19421 -1848
rect 19471 -1847 19505 -1813
rect 19575 -1869 19609 -1835
rect 19672 -1863 19706 -1829
rect 19471 -1915 19505 -1881
rect 19756 -1893 19790 -1859
rect 19963 -1869 19997 -1835
rect 20047 -1843 20081 -1809
rect 20131 -1869 20165 -1835
rect 20253 -1839 20287 -1805
rect 20386 -1845 20420 -1811
rect 20493 -1845 20527 -1811
rect 20839 -1843 20873 -1809
rect 20951 -1839 20985 -1805
rect 21061 -1843 21095 -1809
rect 21273 -1839 21307 -1805
rect 21491 -1859 21525 -1825
rect 21595 -1882 21629 -1848
rect 21679 -1847 21713 -1813
rect 21783 -1869 21817 -1835
rect 21880 -1863 21914 -1829
rect 21679 -1915 21713 -1881
rect 21964 -1893 21998 -1859
rect 14051 -2355 14085 -2321
rect 14055 -2448 14089 -2414
rect 14060 -2558 14094 -2524
rect 14043 -2651 14077 -2617
rect 14055 -2817 14089 -2783
rect 15008 -2766 15042 -2732
rect 15179 -2783 15213 -2749
rect 15288 -2779 15322 -2745
rect 15547 -2753 15581 -2719
rect 15631 -2779 15665 -2745
rect 15715 -2753 15749 -2719
rect 15837 -2783 15871 -2749
rect 15970 -2777 16004 -2743
rect 16077 -2777 16111 -2743
rect 16423 -2779 16457 -2745
rect 16535 -2783 16569 -2749
rect 16645 -2779 16679 -2745
rect 16857 -2783 16891 -2749
rect 17075 -2763 17109 -2729
rect 17179 -2740 17213 -2706
rect 17263 -2707 17297 -2673
rect 17263 -2775 17297 -2741
rect 17367 -2753 17401 -2719
rect 17464 -2759 17498 -2725
rect 17548 -2729 17582 -2695
rect 17755 -2753 17789 -2719
rect 17839 -2779 17873 -2745
rect 17923 -2753 17957 -2719
rect 18045 -2783 18079 -2749
rect 18178 -2777 18212 -2743
rect 18285 -2777 18319 -2743
rect 18631 -2779 18665 -2745
rect 18743 -2783 18777 -2749
rect 18853 -2779 18887 -2745
rect 19065 -2783 19099 -2749
rect 19283 -2763 19317 -2729
rect 19387 -2740 19421 -2706
rect 19471 -2707 19505 -2673
rect 19471 -2775 19505 -2741
rect 19575 -2753 19609 -2719
rect 19672 -2759 19706 -2725
rect 19756 -2729 19790 -2695
rect 19963 -2753 19997 -2719
rect 20047 -2779 20081 -2745
rect 20131 -2753 20165 -2719
rect 20253 -2783 20287 -2749
rect 20386 -2777 20420 -2743
rect 20493 -2777 20527 -2743
rect 20839 -2779 20873 -2745
rect 20951 -2783 20985 -2749
rect 21061 -2779 21095 -2745
rect 21273 -2783 21307 -2749
rect 21491 -2763 21525 -2729
rect 21595 -2740 21629 -2706
rect 21679 -2707 21713 -2673
rect 21679 -2775 21713 -2741
rect 21783 -2753 21817 -2719
rect 21880 -2759 21914 -2725
rect 21964 -2729 21998 -2695
rect 15110 -3254 15144 -3178
rect 15968 -3254 16002 -3178
rect 16214 -5526 16248 -4750
rect 16672 -5526 16706 -4750
rect 17130 -5526 17164 -4750
rect 17588 -5526 17622 -4750
rect 18046 -5526 18080 -4750
rect 18902 -5622 18936 -5546
rect 20560 -5622 20594 -5546
rect 21366 -5494 21400 -5418
rect 21624 -5494 21658 -5418
rect 21882 -5494 21916 -5418
rect 21366 -5704 21400 -5628
rect 21624 -5704 21658 -5628
rect 21882 -5704 21916 -5628
rect 23446 -5436 23572 -5402
rect 23446 -5694 23572 -5660
rect 9220 -7734 9296 -7700
rect 9220 -9392 9296 -9358
<< pdiffc >>
rect 3325 -1393 3359 -1359
rect 3393 -1393 3427 -1359
rect 4903 -1393 4937 -1359
rect 4971 -1393 5005 -1359
rect 3325 -1479 3359 -1445
rect 3393 -1479 3427 -1445
rect 4903 -1479 4937 -1445
rect 4971 -1479 5005 -1445
rect 3312 -1565 3346 -1531
rect 3393 -1565 3427 -1531
rect 4903 -1565 4937 -1531
rect 4984 -1565 5018 -1531
rect 14301 -1819 14335 -1785
rect 14431 -1819 14465 -1785
rect 3366 -2311 3400 -2135
rect 3624 -2311 3658 -2135
rect 4678 -2311 4712 -2135
rect 4936 -2311 4970 -2135
rect 14363 -1903 14397 -1869
rect 14431 -1903 14465 -1869
rect 7476 -2975 7510 -2199
rect 7634 -2975 7668 -2199
rect 7792 -2975 7826 -2199
rect 7950 -2975 7984 -2199
rect 8108 -2975 8142 -2199
rect 8266 -2975 8300 -2199
rect 8424 -2975 8458 -2199
rect 8582 -2975 8616 -2199
rect 8740 -2975 8774 -2199
rect 8898 -2975 8932 -2199
rect 9056 -2975 9090 -2199
rect 14363 -1987 14397 -1953
rect 14439 -2071 14473 -2037
rect 14431 -2175 14465 -2141
rect 14361 -2264 14395 -2230
rect 14431 -2264 14465 -2230
rect 15008 -2235 15042 -2201
rect 15096 -2227 15130 -2193
rect 15248 -2167 15282 -2133
rect 15182 -2235 15216 -2201
rect 15250 -2235 15284 -2201
rect 15336 -2167 15370 -2133
rect 15336 -2235 15370 -2201
rect 15547 -2159 15581 -2125
rect 15547 -2227 15581 -2193
rect 15631 -2211 15665 -2177
rect 15715 -2159 15749 -2125
rect 15715 -2227 15749 -2193
rect 15898 -2235 15932 -2201
rect 15982 -2227 16016 -2193
rect 16075 -2233 16109 -2199
rect 16229 -2209 16263 -2175
rect 16326 -2225 16360 -2191
rect 16410 -2209 16444 -2175
rect 16523 -2235 16557 -2201
rect 16611 -2227 16645 -2193
rect 16708 -2234 16742 -2200
rect 16900 -2235 16934 -2201
rect 16984 -2209 17018 -2175
rect 17070 -2235 17104 -2201
rect 17148 -2235 17182 -2201
rect 17232 -2091 17266 -2057
rect 17464 -2099 17498 -2065
rect 17232 -2159 17266 -2125
rect 17232 -2227 17266 -2193
rect 17367 -2167 17401 -2133
rect 17367 -2235 17401 -2201
rect 17464 -2167 17498 -2133
rect 17464 -2235 17498 -2201
rect 17548 -2131 17582 -2097
rect 17548 -2199 17582 -2165
rect 17755 -2159 17789 -2125
rect 17755 -2227 17789 -2193
rect 17839 -2211 17873 -2177
rect 17923 -2159 17957 -2125
rect 17923 -2227 17957 -2193
rect 18106 -2235 18140 -2201
rect 18190 -2227 18224 -2193
rect 18283 -2233 18317 -2199
rect 18437 -2209 18471 -2175
rect 18534 -2225 18568 -2191
rect 18618 -2209 18652 -2175
rect 18731 -2235 18765 -2201
rect 18819 -2227 18853 -2193
rect 18916 -2234 18950 -2200
rect 19108 -2235 19142 -2201
rect 19192 -2209 19226 -2175
rect 19278 -2235 19312 -2201
rect 19356 -2235 19390 -2201
rect 19440 -2091 19474 -2057
rect 19672 -2099 19706 -2065
rect 19440 -2159 19474 -2125
rect 19440 -2227 19474 -2193
rect 19575 -2167 19609 -2133
rect 19575 -2235 19609 -2201
rect 19672 -2167 19706 -2133
rect 19672 -2235 19706 -2201
rect 19756 -2131 19790 -2097
rect 19756 -2199 19790 -2165
rect 19963 -2159 19997 -2125
rect 19963 -2227 19997 -2193
rect 20047 -2211 20081 -2177
rect 20131 -2159 20165 -2125
rect 20131 -2227 20165 -2193
rect 20314 -2235 20348 -2201
rect 20398 -2227 20432 -2193
rect 20491 -2233 20525 -2199
rect 20645 -2209 20679 -2175
rect 20742 -2225 20776 -2191
rect 20826 -2209 20860 -2175
rect 20939 -2235 20973 -2201
rect 21027 -2227 21061 -2193
rect 21124 -2234 21158 -2200
rect 21316 -2235 21350 -2201
rect 21400 -2209 21434 -2175
rect 21486 -2235 21520 -2201
rect 21564 -2235 21598 -2201
rect 21648 -2091 21682 -2057
rect 21880 -2099 21914 -2065
rect 21648 -2159 21682 -2125
rect 21648 -2227 21682 -2193
rect 21783 -2167 21817 -2133
rect 21783 -2235 21817 -2201
rect 21880 -2167 21914 -2133
rect 21880 -2235 21914 -2201
rect 21964 -2131 21998 -2097
rect 21964 -2199 21998 -2165
rect 14363 -2364 14397 -2330
rect 14431 -2364 14465 -2330
rect 14363 -2448 14397 -2414
rect 14431 -2448 14465 -2414
rect 15008 -2387 15042 -2353
rect 15096 -2395 15130 -2361
rect 15182 -2387 15216 -2353
rect 15250 -2387 15284 -2353
rect 14426 -2558 14460 -2524
rect 15248 -2455 15282 -2421
rect 15336 -2387 15370 -2353
rect 15336 -2455 15370 -2421
rect 14443 -2652 14477 -2618
rect 15547 -2395 15581 -2361
rect 15547 -2463 15581 -2429
rect 15631 -2411 15665 -2377
rect 15715 -2395 15749 -2361
rect 15898 -2387 15932 -2353
rect 15982 -2395 16016 -2361
rect 16075 -2389 16109 -2355
rect 16229 -2413 16263 -2379
rect 16326 -2397 16360 -2363
rect 16410 -2413 16444 -2379
rect 16523 -2387 16557 -2353
rect 15715 -2463 15749 -2429
rect 14431 -2817 14465 -2783
rect 16611 -2395 16645 -2361
rect 16708 -2388 16742 -2354
rect 16900 -2387 16934 -2353
rect 16984 -2413 17018 -2379
rect 17070 -2387 17104 -2353
rect 17148 -2387 17182 -2353
rect 17232 -2395 17266 -2361
rect 17232 -2463 17266 -2429
rect 17367 -2387 17401 -2353
rect 17367 -2455 17401 -2421
rect 17464 -2387 17498 -2353
rect 17464 -2455 17498 -2421
rect 17232 -2531 17266 -2497
rect 17464 -2523 17498 -2489
rect 17548 -2423 17582 -2389
rect 17548 -2491 17582 -2457
rect 17755 -2395 17789 -2361
rect 17755 -2463 17789 -2429
rect 17839 -2411 17873 -2377
rect 17923 -2395 17957 -2361
rect 18106 -2387 18140 -2353
rect 18190 -2395 18224 -2361
rect 18283 -2389 18317 -2355
rect 18437 -2413 18471 -2379
rect 18534 -2397 18568 -2363
rect 18618 -2413 18652 -2379
rect 18731 -2387 18765 -2353
rect 17923 -2463 17957 -2429
rect 18819 -2395 18853 -2361
rect 18916 -2388 18950 -2354
rect 19108 -2387 19142 -2353
rect 19192 -2413 19226 -2379
rect 19278 -2387 19312 -2353
rect 19356 -2387 19390 -2353
rect 19440 -2395 19474 -2361
rect 19440 -2463 19474 -2429
rect 19575 -2387 19609 -2353
rect 19575 -2455 19609 -2421
rect 19672 -2387 19706 -2353
rect 19672 -2455 19706 -2421
rect 19440 -2531 19474 -2497
rect 19672 -2523 19706 -2489
rect 19756 -2423 19790 -2389
rect 19756 -2491 19790 -2457
rect 19963 -2395 19997 -2361
rect 19963 -2463 19997 -2429
rect 20047 -2411 20081 -2377
rect 20131 -2395 20165 -2361
rect 20314 -2387 20348 -2353
rect 20398 -2395 20432 -2361
rect 20491 -2389 20525 -2355
rect 20645 -2413 20679 -2379
rect 20742 -2397 20776 -2363
rect 20826 -2413 20860 -2379
rect 20939 -2387 20973 -2353
rect 20131 -2463 20165 -2429
rect 21027 -2395 21061 -2361
rect 21124 -2388 21158 -2354
rect 21316 -2387 21350 -2353
rect 21400 -2413 21434 -2379
rect 21486 -2387 21520 -2353
rect 21564 -2387 21598 -2353
rect 21648 -2395 21682 -2361
rect 21648 -2463 21682 -2429
rect 21783 -2387 21817 -2353
rect 21783 -2455 21817 -2421
rect 21880 -2387 21914 -2353
rect 21880 -2455 21914 -2421
rect 21648 -2531 21682 -2497
rect 21880 -2523 21914 -2489
rect 21964 -2423 21998 -2389
rect 21964 -2491 21998 -2457
rect 10636 -6377 10670 -6001
rect 11094 -6377 11128 -6001
rect 11208 -6377 11242 -6001
rect 11666 -6377 11700 -6001
rect 11780 -6377 11814 -6001
rect 12238 -6377 12272 -6001
rect 12352 -6377 12386 -6001
rect 12810 -6377 12844 -6001
rect 12924 -6377 12958 -6001
rect 13382 -6377 13416 -6001
rect 13496 -6377 13530 -6001
rect 13954 -6377 13988 -6001
rect 14068 -6377 14102 -6001
rect 14526 -6377 14560 -6001
rect 14640 -6377 14674 -6001
rect 15098 -6377 15132 -6001
rect 10636 -6905 10670 -6529
rect 11094 -6905 11128 -6529
rect 11208 -6905 11242 -6529
rect 11666 -6905 11700 -6529
rect 11780 -6905 11814 -6529
rect 12238 -6905 12272 -6529
rect 12352 -6905 12386 -6529
rect 12810 -6905 12844 -6529
rect 12924 -6905 12958 -6529
rect 13382 -6905 13416 -6529
rect 13496 -6905 13530 -6529
rect 13954 -6905 13988 -6529
rect 14068 -6905 14102 -6529
rect 14526 -6905 14560 -6529
rect 14640 -6905 14674 -6529
rect 15098 -6905 15132 -6529
rect 18882 -6635 18916 -6559
rect 20540 -6635 20574 -6559
rect 21366 -6499 21400 -6423
rect 21624 -6499 21658 -6423
rect 21882 -6499 21916 -6423
rect 21366 -6727 21400 -6651
rect 21624 -6727 21658 -6651
rect 21882 -6727 21916 -6651
rect 23143 -6438 23919 -6404
rect 23143 -6696 23919 -6662
rect 9809 -7468 9885 -7434
rect 9809 -9126 9885 -9092
<< mvndiffc >>
rect 2682 -4714 2716 -4138
rect 2840 -4714 2874 -4138
rect 2998 -4714 3032 -4138
rect 3388 -4714 3422 -4138
rect 3546 -4714 3580 -4138
rect 3704 -4714 3738 -4138
rect 4598 -4714 4632 -4138
rect 4756 -4714 4790 -4138
rect 4914 -4714 4948 -4138
rect 5304 -4714 5338 -4138
rect 5462 -4714 5496 -4138
rect 5620 -4714 5654 -4138
rect 2451 -8041 2485 -7265
rect 2609 -8041 2643 -7265
rect 2767 -8041 2801 -7265
rect 2925 -8041 2959 -7265
rect 3083 -8041 3117 -7265
rect 3241 -8041 3275 -7265
rect 10612 -5346 10646 -4970
rect 11070 -5346 11104 -4970
rect 11190 -5346 11224 -4970
rect 11648 -5346 11682 -4970
rect 11768 -5346 11802 -4970
rect 12226 -5346 12260 -4970
rect 12346 -5346 12380 -4970
rect 12804 -5346 12838 -4970
rect 12924 -5346 12958 -4970
rect 13382 -5346 13416 -4970
rect 13502 -5346 13536 -4970
rect 13960 -5346 13994 -4970
rect 14080 -5346 14114 -4970
rect 14538 -5346 14572 -4970
rect 14658 -5346 14692 -4970
rect 15116 -5346 15150 -4970
rect 7280 -12438 7314 -12262
rect 7538 -12438 7572 -12262
rect 8222 -12382 8256 -12322
rect 9880 -12382 9914 -12322
rect 11538 -12382 11572 -12322
rect 13196 -12382 13230 -12322
rect 20010 -12734 20786 -12700
rect 20920 -12734 21696 -12700
rect 20010 -13192 20786 -13158
rect 20920 -13192 21696 -13158
rect 20010 -13312 20786 -13278
rect 20920 -13312 21696 -13278
rect 20010 -13770 20786 -13736
rect 20920 -13770 21696 -13736
rect 20010 -13890 20786 -13856
rect 20920 -13890 21696 -13856
rect 20010 -14348 20786 -14314
rect 20920 -14348 21696 -14314
rect 20010 -14468 20786 -14434
rect 20920 -14468 21696 -14434
rect 20010 -14926 20786 -14892
rect 20920 -14926 21696 -14892
rect 20010 -15046 20786 -15012
rect 20920 -15046 21696 -15012
rect 20010 -15504 20786 -15470
rect 20920 -15504 21696 -15470
rect 20476 -16078 21252 -16044
rect 20476 -16236 21252 -16202
rect 20476 -16394 21252 -16360
rect 20476 -16552 21252 -16518
rect 20476 -16710 21252 -16676
rect 20476 -16868 21252 -16834
rect 20476 -17026 21252 -16992
rect 20476 -17184 21252 -17150
rect 20476 -17342 21252 -17308
rect 20476 -17500 21252 -17466
rect 20476 -17658 21252 -17624
rect 20476 -17816 21252 -17782
rect 20476 -17974 21252 -17940
<< mvpdiffc >>
rect 11434 -2957 11468 -2181
rect 11592 -2957 11626 -2181
rect 2764 -5617 2798 -5441
rect 3622 -5617 3656 -5441
rect 2764 -6221 2798 -6045
rect 3622 -6221 3656 -6045
rect 4680 -5617 4714 -5441
rect 5538 -5617 5572 -5441
rect 4680 -6221 4714 -6045
rect 5538 -6221 5572 -6045
rect 3826 -8043 3860 -7267
rect 3984 -8043 4018 -7267
rect 4142 -8043 4176 -7267
rect 4300 -8043 4334 -7267
rect 4458 -8043 4492 -7267
rect 4616 -8043 4650 -7267
rect 16214 -6885 16248 -6109
rect 16672 -6885 16706 -6109
rect 17130 -6885 17164 -6109
rect 17588 -6885 17622 -6109
rect 18046 -6885 18080 -6109
rect 22613 -12742 23389 -12708
rect 23541 -12742 24317 -12708
rect 22613 -13200 23389 -13166
rect 23541 -13200 24317 -13166
rect 22613 -13320 23389 -13286
rect 23541 -13320 24317 -13286
rect 22613 -13778 23389 -13744
rect 23541 -13778 24317 -13744
rect 22613 -13898 23389 -13864
rect 23541 -13898 24317 -13864
rect 22613 -14356 23389 -14322
rect 23541 -14356 24317 -14322
rect 22613 -14476 23389 -14442
rect 23541 -14476 24317 -14442
rect 22613 -14934 23389 -14900
rect 23541 -14934 24317 -14900
rect 22613 -15054 23389 -15020
rect 23541 -15054 24317 -15020
rect 22613 -15512 23389 -15478
rect 23541 -15512 24317 -15478
rect 22613 -15632 23389 -15598
rect 23541 -15632 24317 -15598
rect 22613 -16090 23389 -16056
rect 23541 -16090 24317 -16056
rect 22613 -16210 23389 -16176
rect 23541 -16210 24317 -16176
rect 22613 -16668 23389 -16634
rect 23541 -16668 24317 -16634
rect 22613 -16788 23389 -16754
rect 23541 -16788 24317 -16754
rect 22613 -17246 23389 -17212
rect 23541 -17246 24317 -17212
rect 22613 -17366 23389 -17332
rect 23541 -17366 24317 -17332
rect 22613 -17824 23389 -17790
rect 23541 -17824 24317 -17790
<< psubdiff >>
rect 2786 -884 2882 -850
rect 2984 -884 3080 -850
rect 2786 -946 2820 -884
rect 3046 -946 3080 -884
rect 2786 -1110 2820 -1048
rect 3046 -1110 3080 -1048
rect 2786 -1144 2882 -1110
rect 2984 -1144 3080 -1110
rect 5256 -884 5352 -850
rect 5454 -884 5550 -850
rect 5256 -946 5290 -884
rect 5516 -946 5550 -884
rect 5256 -1110 5290 -1048
rect 5516 -1110 5550 -1048
rect 5256 -1144 5352 -1110
rect 5454 -1144 5550 -1110
rect 3014 -1295 3061 -1261
rect 3095 -1295 3119 -1261
rect 5211 -1295 5235 -1261
rect 5269 -1295 5316 -1261
rect 14052 -1721 14099 -1687
rect 14133 -1721 14157 -1687
rect 2652 -1982 2748 -1948
rect 3076 -1982 3172 -1948
rect 2652 -2044 2686 -1982
rect 3138 -2044 3172 -1982
rect 2652 -2462 2686 -2400
rect 3138 -2462 3172 -2400
rect 2652 -2496 2748 -2462
rect 3076 -2496 3172 -2462
rect 5164 -1982 5260 -1948
rect 5588 -1982 5684 -1948
rect 5164 -2044 5198 -1982
rect 5650 -2044 5684 -1982
rect 14897 -1861 14931 -1814
rect 15449 -1861 15483 -1814
rect 14897 -1919 14931 -1895
rect 5164 -2462 5198 -2400
rect 5650 -2462 5684 -2400
rect 5164 -2496 5260 -2462
rect 5588 -2496 5684 -2462
rect 9288 -2052 9384 -2018
rect 11034 -2052 11130 -2018
rect 9288 -2114 9322 -2052
rect 11096 -2114 11130 -2052
rect 9288 -3132 9322 -3070
rect 11096 -3132 11130 -3070
rect 9288 -3166 9384 -3132
rect 11034 -3166 11130 -3132
rect 12600 -2126 12696 -2092
rect 12952 -2126 13048 -2092
rect 12600 -2188 12634 -2126
rect 13014 -2188 13048 -2126
rect 12600 -3178 12634 -3116
rect 15449 -1919 15483 -1895
rect 17657 -1861 17691 -1814
rect 17657 -1919 17691 -1895
rect 19865 -1861 19899 -1814
rect 19865 -1919 19899 -1895
rect 22073 -1861 22107 -1814
rect 22073 -1919 22107 -1895
rect 14897 -2693 14931 -2669
rect 13918 -2754 13978 -2730
rect 15449 -2693 15483 -2669
rect 13918 -2838 13978 -2814
rect 14897 -2774 14931 -2727
rect 15449 -2774 15483 -2727
rect 17657 -2693 17691 -2669
rect 17657 -2774 17691 -2727
rect 19865 -2693 19899 -2669
rect 19865 -2774 19899 -2727
rect 22073 -2693 22107 -2669
rect 22073 -2774 22107 -2727
rect 13014 -3178 13048 -3116
rect 12600 -3212 12696 -3178
rect 12952 -3212 13048 -3178
rect 14996 -3026 15092 -2992
rect 16020 -3026 16116 -2992
rect 14996 -3088 15030 -3026
rect 16082 -3088 16116 -3026
rect 14996 -3406 15030 -3344
rect 16082 -3406 16116 -3344
rect 14996 -3440 15092 -3406
rect 16020 -3440 16116 -3406
rect 16100 -4598 16196 -4564
rect 18098 -4598 18194 -4564
rect 16100 -4660 16134 -4598
rect 18160 -4660 18194 -4598
rect 16100 -5678 16134 -5616
rect 21252 -5266 21348 -5232
rect 21934 -5266 22030 -5232
rect 21252 -5328 21286 -5266
rect 18160 -5678 18194 -5616
rect 16100 -5712 16196 -5678
rect 18098 -5712 18194 -5678
rect 18788 -5394 18884 -5360
rect 20612 -5394 20708 -5360
rect 18788 -5456 18822 -5394
rect 20674 -5456 20708 -5394
rect 18788 -5774 18822 -5712
rect 20674 -5774 20708 -5712
rect 18788 -5808 18884 -5774
rect 20612 -5808 20708 -5774
rect 21996 -5328 22030 -5266
rect 21252 -5856 21286 -5794
rect 21996 -5856 22030 -5794
rect 23260 -5322 23356 -5288
rect 23662 -5322 23758 -5288
rect 23260 -5384 23294 -5322
rect 23724 -5384 23758 -5322
rect 23260 -5774 23294 -5712
rect 23724 -5774 23758 -5712
rect 23260 -5808 23356 -5774
rect 23662 -5808 23758 -5774
rect 21252 -5890 21348 -5856
rect 21934 -5890 22030 -5856
rect 9034 -7620 9130 -7586
rect 9386 -7620 9482 -7586
rect 9034 -7682 9068 -7620
rect 9448 -7682 9482 -7620
rect 9034 -9472 9068 -9410
rect 10490 -7342 10586 -7308
rect 24686 -7342 24782 -7308
rect 10490 -7404 10524 -7342
rect 9448 -9472 9482 -9410
rect 9034 -9506 9130 -9472
rect 9386 -9506 9482 -9472
rect 24748 -7404 24782 -7342
rect 10490 -9928 10524 -9866
rect 24748 -9928 24782 -9866
rect 10490 -9962 10586 -9928
rect 24686 -9962 24782 -9928
rect 3004 -12826 3100 -12792
rect 19000 -12826 19096 -12792
rect 3004 -12888 3038 -12826
rect 19062 -12888 19096 -12826
rect 3004 -13586 3038 -13524
rect 19062 -13586 19096 -13524
rect 3004 -13620 3100 -13586
rect 19000 -13620 19096 -13586
rect 2002 -13764 2098 -13730
rect 19398 -13764 19494 -13730
rect 2002 -13826 2036 -13764
rect 19460 -13826 19494 -13764
rect 2002 -18176 2036 -18114
rect 19460 -18176 19494 -18114
rect 2002 -18210 2098 -18176
rect 19398 -18210 19494 -18176
rect 2000 -18354 2096 -18320
rect 24996 -18354 25092 -18320
rect 2000 -18416 2034 -18354
rect 25058 -18416 25092 -18354
rect 2000 -22600 2034 -22538
rect 25058 -22600 25092 -22538
rect 2000 -22634 2096 -22600
rect 24996 -22634 25092 -22600
rect 21076 -22724 21172 -22690
rect 21550 -22724 21646 -22690
rect 21076 -22786 21110 -22724
rect 20358 -22872 20454 -22838
rect 20556 -22872 20652 -22838
rect 20358 -22934 20392 -22872
rect 20618 -22934 20652 -22872
rect 20358 -23098 20392 -23036
rect 20618 -23098 20652 -23036
rect 20358 -23132 20454 -23098
rect 20556 -23132 20652 -23098
rect 21612 -22786 21646 -22724
rect 21076 -23226 21110 -23164
rect 21612 -23226 21646 -23164
rect 21076 -23260 21172 -23226
rect 21550 -23260 21646 -23226
rect 22502 -22726 22598 -22692
rect 22976 -22726 23072 -22692
rect 22502 -22788 22536 -22726
rect 23038 -22788 23072 -22726
rect 22502 -23228 22536 -23166
rect 23466 -22874 23562 -22840
rect 23664 -22874 23760 -22840
rect 23466 -22936 23500 -22874
rect 23726 -22936 23760 -22874
rect 23466 -23100 23500 -23038
rect 23726 -23100 23760 -23038
rect 23466 -23134 23562 -23100
rect 23664 -23134 23760 -23100
rect 23038 -23228 23072 -23166
rect 22502 -23262 22598 -23228
rect 22976 -23262 23072 -23228
<< nsubdiff >>
rect 3255 -1295 3279 -1261
rect 3313 -1295 3372 -1261
rect 3406 -1295 3430 -1261
rect 4900 -1295 4924 -1261
rect 4958 -1295 5017 -1261
rect 5051 -1295 5075 -1261
rect 14293 -1721 14317 -1687
rect 14351 -1721 14410 -1687
rect 14444 -1721 14468 -1687
rect 3252 -1974 3348 -1940
rect 3676 -1974 3772 -1940
rect 3252 -2036 3286 -1974
rect 3738 -2036 3772 -1974
rect 3252 -2472 3286 -2410
rect 3738 -2472 3772 -2410
rect 3252 -2506 3348 -2472
rect 3676 -2506 3772 -2472
rect 4564 -1974 4660 -1940
rect 4988 -1974 5084 -1940
rect 4564 -2036 4598 -1974
rect 5050 -2036 5084 -1974
rect 4564 -2472 4598 -2410
rect 5050 -2472 5084 -2410
rect 4564 -2506 4660 -2472
rect 4988 -2506 5084 -2472
rect 7362 -2038 7458 -2004
rect 9108 -2038 9204 -2004
rect 7362 -2100 7396 -2038
rect 9170 -2100 9204 -2038
rect 7362 -3136 7396 -3074
rect 9170 -3136 9204 -3074
rect 7362 -3170 7458 -3136
rect 9108 -3170 9204 -3136
rect 14897 -2079 14931 -2055
rect 14897 -2172 14931 -2113
rect 15449 -2079 15483 -2055
rect 14897 -2230 14931 -2206
rect 15449 -2172 15483 -2113
rect 15449 -2230 15483 -2206
rect 17657 -2079 17691 -2055
rect 17657 -2172 17691 -2113
rect 17657 -2230 17691 -2206
rect 19865 -2079 19899 -2055
rect 19865 -2172 19899 -2113
rect 19865 -2230 19899 -2206
rect 22073 -2079 22107 -2055
rect 22073 -2172 22107 -2113
rect 22073 -2230 22107 -2206
rect 14897 -2382 14931 -2358
rect 14897 -2475 14931 -2416
rect 14897 -2533 14931 -2509
rect 15449 -2382 15483 -2358
rect 15449 -2475 15483 -2416
rect 15449 -2533 15483 -2509
rect 17657 -2382 17691 -2358
rect 17657 -2475 17691 -2416
rect 17657 -2533 17691 -2509
rect 19865 -2382 19899 -2358
rect 19865 -2475 19899 -2416
rect 19865 -2533 19899 -2509
rect 22073 -2382 22107 -2358
rect 22073 -2475 22107 -2416
rect 22073 -2533 22107 -2509
rect 1883 -3423 6465 -3403
rect 1883 -3457 1963 -3423
rect 6385 -3457 6465 -3423
rect 1883 -3477 6465 -3457
rect 1883 -3483 1957 -3477
rect 1883 -8969 1903 -3483
rect 1937 -8969 1957 -3483
rect 6391 -3483 6465 -3477
rect 1883 -8975 1957 -8969
rect 6391 -8969 6411 -3483
rect 6445 -8969 6465 -3483
rect 6391 -8975 6465 -8969
rect 1883 -8995 6465 -8975
rect 1883 -9029 1963 -8995
rect 6385 -9029 6465 -8995
rect 1883 -9049 6465 -9029
rect 8737 -4197 25291 -4177
rect 8737 -4231 8817 -4197
rect 25211 -4231 25291 -4197
rect 8737 -4251 25291 -4231
rect 8737 -4257 8811 -4251
rect 8737 -10275 8757 -4257
rect 8791 -10275 8811 -4257
rect 25217 -4257 25291 -4251
rect 10522 -5840 10618 -5806
rect 15150 -5840 15246 -5806
rect 10522 -5902 10556 -5840
rect 15212 -5902 15246 -5840
rect 10522 -7066 10556 -7004
rect 15212 -7066 15246 -7004
rect 10522 -7100 10618 -7066
rect 15150 -7100 15246 -7066
rect 21252 -6262 21348 -6228
rect 21934 -6262 22030 -6228
rect 21252 -6324 21286 -6262
rect 18768 -6398 18864 -6364
rect 20592 -6398 20688 -6364
rect 18768 -6460 18802 -6398
rect 20654 -6460 20688 -6398
rect 18768 -6796 18802 -6734
rect 20654 -6796 20688 -6734
rect 18768 -6830 18864 -6796
rect 20592 -6830 20688 -6796
rect 21996 -6324 22030 -6262
rect 21252 -6888 21286 -6826
rect 22948 -6324 23044 -6290
rect 24018 -6324 24114 -6290
rect 22948 -6386 22982 -6324
rect 24080 -6386 24114 -6324
rect 22948 -6776 22982 -6714
rect 24080 -6776 24114 -6714
rect 22948 -6810 23044 -6776
rect 24018 -6810 24114 -6776
rect 21996 -6888 22030 -6826
rect 21252 -6922 21348 -6888
rect 21934 -6922 22030 -6888
rect 9614 -7354 9710 -7320
rect 9984 -7354 10080 -7320
rect 9614 -7416 9648 -7354
rect 10046 -7416 10080 -7354
rect 9614 -9206 9648 -9144
rect 10046 -9206 10080 -9144
rect 9614 -9240 9710 -9206
rect 9984 -9240 10080 -9206
rect 8737 -10281 8811 -10275
rect 25217 -10275 25237 -4257
rect 25271 -10275 25291 -4257
rect 25217 -10281 25291 -10275
rect 8737 -10301 25291 -10281
rect 8737 -10335 8817 -10301
rect 25211 -10335 25291 -10301
rect 8737 -10355 25291 -10335
rect 1663 -11595 25533 -11575
rect 1663 -11629 1743 -11595
rect 25453 -11629 25533 -11595
rect 1663 -11649 25533 -11629
rect 1663 -11655 1737 -11649
rect 1663 -23587 1683 -11655
rect 1717 -23587 1737 -11655
rect 25459 -11655 25533 -11649
rect 21214 -22862 21310 -22828
rect 21412 -22862 21508 -22828
rect 21214 -22924 21248 -22862
rect 21474 -22924 21508 -22862
rect 21214 -23088 21248 -23026
rect 21474 -23088 21508 -23026
rect 21214 -23122 21310 -23088
rect 21412 -23122 21508 -23088
rect 22640 -22864 22736 -22830
rect 22838 -22864 22934 -22830
rect 22640 -22926 22674 -22864
rect 22900 -22926 22934 -22864
rect 22640 -23090 22674 -23028
rect 22900 -23090 22934 -23028
rect 22640 -23124 22736 -23090
rect 22838 -23124 22934 -23090
rect 1663 -23593 1737 -23587
rect 25459 -23587 25479 -11655
rect 25513 -23587 25533 -11655
rect 25459 -23593 25533 -23587
rect 1663 -23613 25533 -23593
rect 1663 -23647 1743 -23613
rect 25453 -23647 25533 -23613
rect 1663 -23667 25533 -23647
<< mvpsubdiff >>
rect 2536 -3916 3178 -3904
rect 2536 -3950 2644 -3916
rect 3070 -3950 3178 -3916
rect 2536 -3962 3178 -3950
rect 2536 -4012 2594 -3962
rect 2536 -4840 2548 -4012
rect 2582 -4840 2594 -4012
rect 3120 -4012 3178 -3962
rect 2536 -4890 2594 -4840
rect 3120 -4840 3132 -4012
rect 3166 -4840 3178 -4012
rect 3120 -4890 3178 -4840
rect 2536 -4902 3178 -4890
rect 2536 -4936 2644 -4902
rect 3070 -4936 3178 -4902
rect 2536 -4948 3178 -4936
rect 3242 -3916 3884 -3904
rect 3242 -3950 3350 -3916
rect 3776 -3950 3884 -3916
rect 3242 -3962 3884 -3950
rect 3242 -4012 3300 -3962
rect 3242 -4840 3254 -4012
rect 3288 -4840 3300 -4012
rect 3826 -4012 3884 -3962
rect 3242 -4890 3300 -4840
rect 3826 -4840 3838 -4012
rect 3872 -4840 3884 -4012
rect 3826 -4890 3884 -4840
rect 3242 -4902 3884 -4890
rect 3242 -4936 3350 -4902
rect 3776 -4936 3884 -4902
rect 3242 -4948 3884 -4936
rect 4452 -3916 5094 -3904
rect 4452 -3950 4560 -3916
rect 4986 -3950 5094 -3916
rect 4452 -3962 5094 -3950
rect 4452 -4012 4510 -3962
rect 4452 -4840 4464 -4012
rect 4498 -4840 4510 -4012
rect 5036 -4012 5094 -3962
rect 4452 -4890 4510 -4840
rect 5036 -4840 5048 -4012
rect 5082 -4840 5094 -4012
rect 5036 -4890 5094 -4840
rect 4452 -4902 5094 -4890
rect 4452 -4936 4560 -4902
rect 4986 -4936 5094 -4902
rect 4452 -4948 5094 -4936
rect 5158 -3916 5800 -3904
rect 5158 -3950 5266 -3916
rect 5692 -3950 5800 -3916
rect 5158 -3962 5800 -3950
rect 5158 -4012 5216 -3962
rect 5158 -4840 5170 -4012
rect 5204 -4840 5216 -4012
rect 5742 -4012 5800 -3962
rect 5158 -4890 5216 -4840
rect 5742 -4840 5754 -4012
rect 5788 -4840 5800 -4012
rect 5742 -4890 5800 -4840
rect 5158 -4902 5800 -4890
rect 5158 -4936 5266 -4902
rect 5692 -4936 5800 -4902
rect 5158 -4948 5800 -4936
rect 2305 -7043 3421 -7031
rect 2305 -7077 2413 -7043
rect 3313 -7077 3421 -7043
rect 2305 -7089 3421 -7077
rect 2305 -7139 2363 -7089
rect 2305 -8167 2317 -7139
rect 2351 -8167 2363 -7139
rect 3363 -7139 3421 -7089
rect 2305 -8217 2363 -8167
rect 3363 -8167 3375 -7139
rect 3409 -8167 3421 -7139
rect 3363 -8217 3421 -8167
rect 2305 -8229 3421 -8217
rect 2305 -8263 2413 -8229
rect 3313 -8263 3421 -8229
rect 2305 -8275 3421 -8263
rect 10466 -4748 15296 -4736
rect 10466 -4782 10574 -4748
rect 15188 -4782 15296 -4748
rect 10466 -4794 15296 -4782
rect 10466 -4844 10524 -4794
rect 10466 -5472 10478 -4844
rect 10512 -5472 10524 -4844
rect 15238 -4844 15296 -4794
rect 10466 -5522 10524 -5472
rect 15238 -5472 15250 -4844
rect 15284 -5472 15296 -4844
rect 15238 -5522 15296 -5472
rect 10466 -5534 15296 -5522
rect 10466 -5568 10574 -5534
rect 15188 -5568 15296 -5534
rect 10466 -5580 15296 -5568
rect 7134 -12040 7718 -12028
rect 7134 -12074 7242 -12040
rect 7610 -12074 7718 -12040
rect 7134 -12086 7718 -12074
rect 7134 -12136 7192 -12086
rect 7134 -12564 7146 -12136
rect 7180 -12564 7192 -12136
rect 7660 -12136 7718 -12086
rect 7134 -12614 7192 -12564
rect 7660 -12564 7672 -12136
rect 7706 -12564 7718 -12136
rect 7660 -12614 7718 -12564
rect 7134 -12626 7718 -12614
rect 8076 -12100 13376 -12088
rect 8076 -12134 8184 -12100
rect 13268 -12134 13376 -12100
rect 8076 -12146 13376 -12134
rect 8076 -12196 8134 -12146
rect 8076 -12508 8088 -12196
rect 8122 -12508 8134 -12196
rect 13318 -12196 13376 -12146
rect 8076 -12558 8134 -12508
rect 13318 -12508 13330 -12196
rect 13364 -12508 13376 -12196
rect 13318 -12558 13376 -12508
rect 8076 -12570 13376 -12558
rect 8076 -12604 8184 -12570
rect 13268 -12604 13376 -12570
rect 8076 -12616 13376 -12604
rect 19776 -12566 21930 -12554
rect 19776 -12600 19884 -12566
rect 21822 -12600 21930 -12566
rect 19776 -12612 21930 -12600
rect 7134 -12660 7242 -12626
rect 7610 -12660 7718 -12626
rect 7134 -12672 7718 -12660
rect 19776 -12662 19834 -12612
rect 19776 -15542 19788 -12662
rect 19822 -15542 19834 -12662
rect 21872 -12662 21930 -12612
rect 19776 -15592 19834 -15542
rect 21872 -15542 21884 -12662
rect 21918 -15542 21930 -12662
rect 21872 -15592 21930 -15542
rect 19776 -15604 21930 -15592
rect 19776 -15638 19884 -15604
rect 21822 -15638 21930 -15604
rect 19776 -15650 21930 -15638
rect 20242 -15910 21486 -15898
rect 20242 -15944 20350 -15910
rect 21378 -15944 21486 -15910
rect 20242 -15956 21486 -15944
rect 20242 -16006 20300 -15956
rect 20242 -18012 20254 -16006
rect 20288 -18012 20300 -16006
rect 21428 -16006 21486 -15956
rect 20242 -18062 20300 -18012
rect 21428 -18012 21440 -16006
rect 21474 -18012 21486 -16006
rect 21428 -18062 21486 -18012
rect 20242 -18074 21486 -18062
rect 20242 -18108 20350 -18074
rect 21378 -18108 21486 -18074
rect 20242 -18120 21486 -18108
<< mvnsubdiff >>
rect 11288 -1950 11772 -1938
rect 11288 -1984 11396 -1950
rect 11664 -1984 11772 -1950
rect 11288 -1996 11772 -1984
rect 11288 -2046 11346 -1996
rect 11288 -3092 11300 -2046
rect 11334 -3092 11346 -2046
rect 11714 -2046 11772 -1996
rect 11288 -3142 11346 -3092
rect 11714 -3092 11726 -2046
rect 11760 -3092 11772 -2046
rect 11714 -3142 11772 -3092
rect 11288 -3154 11772 -3142
rect 11288 -3188 11396 -3154
rect 11664 -3188 11772 -3154
rect 11288 -3200 11772 -3188
rect 2618 -5210 3802 -5198
rect 2618 -5244 2726 -5210
rect 3694 -5244 3802 -5210
rect 2618 -5256 3802 -5244
rect 2618 -5306 2676 -5256
rect 2618 -5752 2630 -5306
rect 2664 -5752 2676 -5306
rect 3744 -5306 3802 -5256
rect 2618 -5802 2676 -5752
rect 3744 -5752 3756 -5306
rect 3790 -5752 3802 -5306
rect 3744 -5802 3802 -5752
rect 2618 -5814 3802 -5802
rect 2618 -5848 2726 -5814
rect 3694 -5848 3802 -5814
rect 2618 -5860 3802 -5848
rect 2618 -5910 2676 -5860
rect 2618 -6356 2630 -5910
rect 2664 -6356 2676 -5910
rect 3744 -5910 3802 -5860
rect 2618 -6406 2676 -6356
rect 3744 -6356 3756 -5910
rect 3790 -6356 3802 -5910
rect 3744 -6406 3802 -6356
rect 2618 -6418 3802 -6406
rect 2618 -6452 2726 -6418
rect 3694 -6452 3802 -6418
rect 2618 -6464 3802 -6452
rect 4534 -5210 5718 -5198
rect 4534 -5244 4642 -5210
rect 5610 -5244 5718 -5210
rect 4534 -5256 5718 -5244
rect 4534 -5306 4592 -5256
rect 4534 -5752 4546 -5306
rect 4580 -5752 4592 -5306
rect 5660 -5306 5718 -5256
rect 4534 -5802 4592 -5752
rect 5660 -5752 5672 -5306
rect 5706 -5752 5718 -5306
rect 5660 -5802 5718 -5752
rect 4534 -5814 5718 -5802
rect 4534 -5848 4642 -5814
rect 5610 -5848 5718 -5814
rect 4534 -5860 5718 -5848
rect 4534 -5910 4592 -5860
rect 4534 -6356 4546 -5910
rect 4580 -6356 4592 -5910
rect 5660 -5910 5718 -5860
rect 4534 -6406 4592 -6356
rect 5660 -6356 5672 -5910
rect 5706 -6356 5718 -5910
rect 5660 -6406 5718 -6356
rect 4534 -6418 5718 -6406
rect 4534 -6452 4642 -6418
rect 5610 -6452 5718 -6418
rect 4534 -6464 5718 -6452
rect 3680 -7036 4796 -7024
rect 3680 -7070 3788 -7036
rect 4688 -7070 4796 -7036
rect 3680 -7082 4796 -7070
rect 3680 -7132 3738 -7082
rect 3680 -8178 3692 -7132
rect 3726 -8178 3738 -7132
rect 4738 -7132 4796 -7082
rect 3680 -8228 3738 -8178
rect 4738 -8178 4750 -7132
rect 4784 -8178 4796 -7132
rect 4738 -8228 4796 -8178
rect 3680 -8240 4796 -8228
rect 3680 -8274 3788 -8240
rect 4688 -8274 4796 -8240
rect 3680 -8286 4796 -8274
rect 16068 -5878 18226 -5866
rect 16068 -5912 16176 -5878
rect 18118 -5912 18226 -5878
rect 16068 -5924 18226 -5912
rect 16068 -5974 16126 -5924
rect 16068 -7020 16080 -5974
rect 16114 -7020 16126 -5974
rect 18168 -5974 18226 -5924
rect 16068 -7070 16126 -7020
rect 18168 -7020 18180 -5974
rect 18214 -7020 18226 -5974
rect 18168 -7070 18226 -7020
rect 16068 -7082 18226 -7070
rect 16068 -7116 16176 -7082
rect 18118 -7116 18226 -7082
rect 16068 -7128 18226 -7116
rect 22370 -12574 24560 -12562
rect 22370 -12608 22478 -12574
rect 24452 -12608 24560 -12574
rect 22370 -12620 24560 -12608
rect 22370 -12670 22428 -12620
rect 22370 -17862 22382 -12670
rect 22416 -17862 22428 -12670
rect 24502 -12670 24560 -12620
rect 22370 -17912 22428 -17862
rect 24502 -17862 24514 -12670
rect 24548 -17862 24560 -12670
rect 24502 -17912 24560 -17862
rect 22370 -17924 24560 -17912
rect 22370 -17958 22478 -17924
rect 24452 -17958 24560 -17924
rect 22370 -17970 24560 -17958
<< psubdiffcont >>
rect 2882 -884 2984 -850
rect 2786 -1048 2820 -946
rect 3046 -1048 3080 -946
rect 2882 -1144 2984 -1110
rect 5352 -884 5454 -850
rect 5256 -1048 5290 -946
rect 5516 -1048 5550 -946
rect 5352 -1144 5454 -1110
rect 3061 -1295 3095 -1261
rect 5235 -1295 5269 -1261
rect 14099 -1721 14133 -1687
rect 2748 -1982 3076 -1948
rect 2652 -2400 2686 -2044
rect 3138 -2400 3172 -2044
rect 2748 -2496 3076 -2462
rect 5260 -1982 5588 -1948
rect 5164 -2400 5198 -2044
rect 14897 -1895 14931 -1861
rect 5650 -2400 5684 -2044
rect 5260 -2496 5588 -2462
rect 9384 -2052 11034 -2018
rect 9288 -3070 9322 -2114
rect 11096 -3070 11130 -2114
rect 9384 -3166 11034 -3132
rect 12696 -2126 12952 -2092
rect 12600 -3116 12634 -2188
rect 13014 -3116 13048 -2188
rect 15449 -1895 15483 -1861
rect 17657 -1895 17691 -1861
rect 19865 -1895 19899 -1861
rect 22073 -1895 22107 -1861
rect 14897 -2727 14931 -2693
rect 13918 -2814 13978 -2754
rect 15449 -2727 15483 -2693
rect 17657 -2727 17691 -2693
rect 19865 -2727 19899 -2693
rect 22073 -2727 22107 -2693
rect 12696 -3212 12952 -3178
rect 15092 -3026 16020 -2992
rect 14996 -3344 15030 -3088
rect 16082 -3344 16116 -3088
rect 15092 -3440 16020 -3406
rect 16196 -4598 18098 -4564
rect 16100 -5616 16134 -4660
rect 18160 -5616 18194 -4660
rect 21348 -5266 21934 -5232
rect 16196 -5712 18098 -5678
rect 18884 -5394 20612 -5360
rect 18788 -5712 18822 -5456
rect 20674 -5712 20708 -5456
rect 18884 -5808 20612 -5774
rect 21252 -5794 21286 -5328
rect 21996 -5794 22030 -5328
rect 23356 -5322 23662 -5288
rect 23260 -5712 23294 -5384
rect 23724 -5712 23758 -5384
rect 23356 -5808 23662 -5774
rect 21348 -5890 21934 -5856
rect 9130 -7620 9386 -7586
rect 9034 -9410 9068 -7682
rect 9448 -9410 9482 -7682
rect 10586 -7342 24686 -7308
rect 9130 -9506 9386 -9472
rect 10490 -9866 10524 -7404
rect 24748 -9866 24782 -7404
rect 10586 -9962 24686 -9928
rect 3100 -12826 19000 -12792
rect 3004 -13524 3038 -12888
rect 19062 -13524 19096 -12888
rect 3100 -13620 19000 -13586
rect 2098 -13764 19398 -13730
rect 2002 -18114 2036 -13826
rect 19460 -18114 19494 -13826
rect 2098 -18210 19398 -18176
rect 2096 -18354 24996 -18320
rect 2000 -22538 2034 -18416
rect 25058 -22538 25092 -18416
rect 2096 -22634 24996 -22600
rect 21172 -22724 21550 -22690
rect 20454 -22872 20556 -22838
rect 20358 -23036 20392 -22934
rect 20618 -23036 20652 -22934
rect 20454 -23132 20556 -23098
rect 21076 -23164 21110 -22786
rect 21612 -23164 21646 -22786
rect 21172 -23260 21550 -23226
rect 22598 -22726 22976 -22692
rect 22502 -23166 22536 -22788
rect 23038 -23166 23072 -22788
rect 23562 -22874 23664 -22840
rect 23466 -23038 23500 -22936
rect 23726 -23038 23760 -22936
rect 23562 -23134 23664 -23100
rect 22598 -23262 22976 -23228
<< nsubdiffcont >>
rect 3279 -1295 3313 -1261
rect 3372 -1295 3406 -1261
rect 4924 -1295 4958 -1261
rect 5017 -1295 5051 -1261
rect 14317 -1721 14351 -1687
rect 14410 -1721 14444 -1687
rect 3348 -1974 3676 -1940
rect 3252 -2410 3286 -2036
rect 3738 -2410 3772 -2036
rect 3348 -2506 3676 -2472
rect 4660 -1974 4988 -1940
rect 4564 -2410 4598 -2036
rect 5050 -2410 5084 -2036
rect 4660 -2506 4988 -2472
rect 7458 -2038 9108 -2004
rect 7362 -3074 7396 -2100
rect 9170 -3074 9204 -2100
rect 7458 -3170 9108 -3136
rect 14897 -2113 14931 -2079
rect 15449 -2113 15483 -2079
rect 14897 -2206 14931 -2172
rect 15449 -2206 15483 -2172
rect 17657 -2113 17691 -2079
rect 17657 -2206 17691 -2172
rect 19865 -2113 19899 -2079
rect 19865 -2206 19899 -2172
rect 22073 -2113 22107 -2079
rect 22073 -2206 22107 -2172
rect 14897 -2416 14931 -2382
rect 14897 -2509 14931 -2475
rect 15449 -2416 15483 -2382
rect 15449 -2509 15483 -2475
rect 17657 -2416 17691 -2382
rect 17657 -2509 17691 -2475
rect 19865 -2416 19899 -2382
rect 19865 -2509 19899 -2475
rect 22073 -2416 22107 -2382
rect 22073 -2509 22107 -2475
rect 1963 -3457 6385 -3423
rect 1903 -8969 1937 -3483
rect 6411 -8969 6445 -3483
rect 1963 -9029 6385 -8995
rect 8817 -4231 25211 -4197
rect 8757 -10275 8791 -4257
rect 10618 -5840 15150 -5806
rect 10522 -7004 10556 -5902
rect 15212 -7004 15246 -5902
rect 10618 -7100 15150 -7066
rect 21348 -6262 21934 -6228
rect 18864 -6398 20592 -6364
rect 18768 -6734 18802 -6460
rect 20654 -6734 20688 -6460
rect 18864 -6830 20592 -6796
rect 21252 -6826 21286 -6324
rect 21996 -6826 22030 -6324
rect 23044 -6324 24018 -6290
rect 22948 -6714 22982 -6386
rect 24080 -6714 24114 -6386
rect 23044 -6810 24018 -6776
rect 21348 -6922 21934 -6888
rect 9710 -7354 9984 -7320
rect 9614 -9144 9648 -7416
rect 10046 -9144 10080 -7416
rect 9710 -9240 9984 -9206
rect 25237 -10275 25271 -4257
rect 8817 -10335 25211 -10301
rect 1743 -11629 25453 -11595
rect 1683 -23587 1717 -11655
rect 21310 -22862 21412 -22828
rect 21214 -23026 21248 -22924
rect 21474 -23026 21508 -22924
rect 21310 -23122 21412 -23088
rect 22736 -22864 22838 -22830
rect 22640 -23028 22674 -22926
rect 22900 -23028 22934 -22926
rect 22736 -23124 22838 -23090
rect 25479 -23587 25513 -11655
rect 1743 -23647 25453 -23613
<< mvpsubdiffcont >>
rect 2644 -3950 3070 -3916
rect 2548 -4840 2582 -4012
rect 3132 -4840 3166 -4012
rect 2644 -4936 3070 -4902
rect 3350 -3950 3776 -3916
rect 3254 -4840 3288 -4012
rect 3838 -4840 3872 -4012
rect 3350 -4936 3776 -4902
rect 4560 -3950 4986 -3916
rect 4464 -4840 4498 -4012
rect 5048 -4840 5082 -4012
rect 4560 -4936 4986 -4902
rect 5266 -3950 5692 -3916
rect 5170 -4840 5204 -4012
rect 5754 -4840 5788 -4012
rect 5266 -4936 5692 -4902
rect 2413 -7077 3313 -7043
rect 2317 -8167 2351 -7139
rect 3375 -8167 3409 -7139
rect 2413 -8263 3313 -8229
rect 10574 -4782 15188 -4748
rect 10478 -5472 10512 -4844
rect 15250 -5472 15284 -4844
rect 10574 -5568 15188 -5534
rect 7242 -12074 7610 -12040
rect 7146 -12564 7180 -12136
rect 7672 -12564 7706 -12136
rect 8184 -12134 13268 -12100
rect 8088 -12508 8122 -12196
rect 13330 -12508 13364 -12196
rect 8184 -12604 13268 -12570
rect 19884 -12600 21822 -12566
rect 7242 -12660 7610 -12626
rect 19788 -15542 19822 -12662
rect 21884 -15542 21918 -12662
rect 19884 -15638 21822 -15604
rect 20350 -15944 21378 -15910
rect 20254 -18012 20288 -16006
rect 21440 -18012 21474 -16006
rect 20350 -18108 21378 -18074
<< mvnsubdiffcont >>
rect 11396 -1984 11664 -1950
rect 11300 -3092 11334 -2046
rect 11726 -3092 11760 -2046
rect 11396 -3188 11664 -3154
rect 2726 -5244 3694 -5210
rect 2630 -5752 2664 -5306
rect 3756 -5752 3790 -5306
rect 2726 -5848 3694 -5814
rect 2630 -6356 2664 -5910
rect 3756 -6356 3790 -5910
rect 2726 -6452 3694 -6418
rect 4642 -5244 5610 -5210
rect 4546 -5752 4580 -5306
rect 5672 -5752 5706 -5306
rect 4642 -5848 5610 -5814
rect 4546 -6356 4580 -5910
rect 5672 -6356 5706 -5910
rect 4642 -6452 5610 -6418
rect 3788 -7070 4688 -7036
rect 3692 -8178 3726 -7132
rect 4750 -8178 4784 -7132
rect 3788 -8274 4688 -8240
rect 16176 -5912 18118 -5878
rect 16080 -7020 16114 -5974
rect 18180 -7020 18214 -5974
rect 16176 -7116 18118 -7082
rect 22478 -12608 24452 -12574
rect 22382 -17862 22416 -12670
rect 24514 -17862 24548 -12670
rect 22478 -17958 24452 -17924
<< poly >>
rect 3149 -1361 3215 -1351
rect 3149 -1395 3165 -1361
rect 3199 -1395 3215 -1361
rect 3149 -1397 3215 -1395
rect 3116 -1403 3274 -1397
rect 5115 -1361 5181 -1351
rect 5115 -1395 5131 -1361
rect 5165 -1395 5181 -1361
rect 5115 -1397 5181 -1395
rect 5056 -1403 5214 -1397
rect 2971 -1433 2997 -1403
rect 3101 -1427 3289 -1403
rect 3101 -1433 3140 -1427
rect 3250 -1433 3289 -1427
rect 3447 -1433 3473 -1403
rect 4857 -1433 4883 -1403
rect 5041 -1427 5229 -1403
rect 5041 -1433 5080 -1427
rect 5190 -1433 5229 -1427
rect 5333 -1433 5359 -1403
rect 3162 -1479 3228 -1469
rect 3162 -1491 3178 -1479
rect 2971 -1521 2997 -1491
rect 3101 -1513 3178 -1491
rect 3212 -1491 3228 -1479
rect 5102 -1479 5168 -1469
rect 5102 -1491 5118 -1479
rect 3212 -1513 3289 -1491
rect 3101 -1521 3289 -1513
rect 3447 -1521 3473 -1491
rect 4857 -1521 4883 -1491
rect 5041 -1513 5118 -1491
rect 5152 -1491 5168 -1479
rect 5152 -1513 5229 -1491
rect 5041 -1521 5229 -1513
rect 5333 -1521 5359 -1491
rect 3162 -1523 3228 -1521
rect 5102 -1523 5168 -1521
rect 14187 -1788 14253 -1778
rect 14187 -1822 14203 -1788
rect 14237 -1822 14253 -1788
rect 14187 -1829 14253 -1822
rect 15053 -1797 15083 -1771
rect 15125 -1797 15155 -1771
rect 15247 -1797 15277 -1771
rect 15591 -1797 15621 -1771
rect 15675 -1797 15705 -1771
rect 15930 -1797 15960 -1771
rect 16025 -1797 16055 -1771
rect 16121 -1797 16151 -1771
rect 16287 -1797 16317 -1771
rect 16359 -1797 16389 -1771
rect 16491 -1797 16521 -1771
rect 16590 -1797 16620 -1771
rect 16699 -1797 16729 -1771
rect 16795 -1797 16825 -1771
rect 16944 -1797 16974 -1771
rect 17035 -1797 17065 -1771
rect 17223 -1797 17253 -1771
rect 17411 -1797 17441 -1771
rect 17508 -1797 17538 -1771
rect 17799 -1797 17829 -1771
rect 17883 -1797 17913 -1771
rect 18138 -1797 18168 -1771
rect 18233 -1797 18263 -1771
rect 18329 -1797 18359 -1771
rect 18495 -1797 18525 -1771
rect 18567 -1797 18597 -1771
rect 18699 -1797 18729 -1771
rect 18798 -1797 18828 -1771
rect 18907 -1797 18937 -1771
rect 19003 -1797 19033 -1771
rect 19152 -1797 19182 -1771
rect 19243 -1797 19273 -1771
rect 19431 -1797 19461 -1771
rect 19619 -1797 19649 -1771
rect 19716 -1797 19746 -1771
rect 20007 -1797 20037 -1771
rect 20091 -1797 20121 -1771
rect 20346 -1797 20376 -1771
rect 20441 -1797 20471 -1771
rect 20537 -1797 20567 -1771
rect 20703 -1797 20733 -1771
rect 20775 -1797 20805 -1771
rect 20907 -1797 20937 -1771
rect 21006 -1797 21036 -1771
rect 21115 -1797 21145 -1771
rect 21211 -1797 21241 -1771
rect 21360 -1797 21390 -1771
rect 21451 -1797 21481 -1771
rect 21639 -1797 21669 -1771
rect 21827 -1797 21857 -1771
rect 21924 -1797 21954 -1771
rect 14009 -1859 14035 -1829
rect 14165 -1859 14285 -1829
rect 14485 -1859 14511 -1829
rect 14187 -1911 14253 -1901
rect 14187 -1925 14203 -1911
rect 2812 -2050 3012 -2034
rect 2812 -2084 2828 -2050
rect 2996 -2084 3012 -2050
rect 2812 -2122 3012 -2084
rect 2812 -2360 3012 -2322
rect 2812 -2394 2828 -2360
rect 2996 -2394 3012 -2360
rect 2812 -2410 3012 -2394
rect 3412 -2042 3612 -2026
rect 3412 -2076 3428 -2042
rect 3596 -2076 3612 -2042
rect 3412 -2123 3612 -2076
rect 3412 -2370 3612 -2323
rect 3412 -2404 3428 -2370
rect 3596 -2404 3612 -2370
rect 3412 -2420 3612 -2404
rect 4724 -2042 4924 -2026
rect 4724 -2076 4740 -2042
rect 4908 -2076 4924 -2042
rect 4724 -2123 4924 -2076
rect 4724 -2370 4924 -2323
rect 4724 -2404 4740 -2370
rect 4908 -2404 4924 -2370
rect 4724 -2420 4924 -2404
rect 5324 -2050 5524 -2034
rect 5324 -2084 5340 -2050
rect 5508 -2084 5524 -2050
rect 5324 -2122 5524 -2084
rect 14009 -1955 14035 -1925
rect 14165 -1945 14203 -1925
rect 14237 -1913 14253 -1911
rect 14237 -1943 14285 -1913
rect 14485 -1943 14511 -1913
rect 14237 -1945 14253 -1943
rect 14165 -1955 14253 -1945
rect 5324 -2360 5524 -2322
rect 5324 -2394 5340 -2360
rect 5508 -2394 5524 -2360
rect 5324 -2410 5524 -2394
rect 7522 -2106 7622 -2090
rect 7522 -2140 7538 -2106
rect 7606 -2140 7622 -2106
rect 7522 -2187 7622 -2140
rect 7680 -2106 7780 -2090
rect 7680 -2140 7696 -2106
rect 7764 -2140 7780 -2106
rect 7680 -2187 7780 -2140
rect 7838 -2106 7938 -2090
rect 7838 -2140 7854 -2106
rect 7922 -2140 7938 -2106
rect 7838 -2187 7938 -2140
rect 7996 -2106 8096 -2090
rect 7996 -2140 8012 -2106
rect 8080 -2140 8096 -2106
rect 7996 -2187 8096 -2140
rect 8154 -2106 8254 -2090
rect 8154 -2140 8170 -2106
rect 8238 -2140 8254 -2106
rect 8154 -2187 8254 -2140
rect 8312 -2106 8412 -2090
rect 8312 -2140 8328 -2106
rect 8396 -2140 8412 -2106
rect 8312 -2187 8412 -2140
rect 8470 -2106 8570 -2090
rect 8470 -2140 8486 -2106
rect 8554 -2140 8570 -2106
rect 8470 -2187 8570 -2140
rect 8628 -2106 8728 -2090
rect 8628 -2140 8644 -2106
rect 8712 -2140 8728 -2106
rect 8628 -2187 8728 -2140
rect 8786 -2106 8886 -2090
rect 8786 -2140 8802 -2106
rect 8870 -2140 8886 -2106
rect 8786 -2187 8886 -2140
rect 8944 -2106 9044 -2090
rect 8944 -2140 8960 -2106
rect 9028 -2140 9044 -2106
rect 8944 -2187 9044 -2140
rect 7522 -3034 7622 -2987
rect 7522 -3068 7538 -3034
rect 7606 -3068 7622 -3034
rect 7522 -3084 7622 -3068
rect 7680 -3034 7780 -2987
rect 7680 -3068 7696 -3034
rect 7764 -3068 7780 -3034
rect 7680 -3084 7780 -3068
rect 7838 -3034 7938 -2987
rect 7838 -3068 7854 -3034
rect 7922 -3068 7938 -3034
rect 7838 -3084 7938 -3068
rect 7996 -3034 8096 -2987
rect 7996 -3068 8012 -3034
rect 8080 -3068 8096 -3034
rect 7996 -3084 8096 -3068
rect 8154 -3034 8254 -2987
rect 8154 -3068 8170 -3034
rect 8238 -3068 8254 -3034
rect 8154 -3084 8254 -3068
rect 8312 -3034 8412 -2987
rect 8312 -3068 8328 -3034
rect 8396 -3068 8412 -3034
rect 8312 -3084 8412 -3068
rect 8470 -3034 8570 -2987
rect 8470 -3068 8486 -3034
rect 8554 -3068 8570 -3034
rect 8470 -3084 8570 -3068
rect 8628 -3034 8728 -2987
rect 8628 -3068 8644 -3034
rect 8712 -3068 8728 -3034
rect 8628 -3084 8728 -3068
rect 8786 -3034 8886 -2987
rect 8786 -3068 8802 -3034
rect 8870 -3068 8886 -3034
rect 8786 -3084 8886 -3068
rect 8944 -3034 9044 -2987
rect 8944 -3068 8960 -3034
rect 9028 -3068 9044 -3034
rect 8944 -3084 9044 -3068
rect 9448 -2120 9548 -2104
rect 9448 -2154 9464 -2120
rect 9532 -2154 9548 -2120
rect 9448 -2192 9548 -2154
rect 9606 -2120 9706 -2104
rect 9606 -2154 9622 -2120
rect 9690 -2154 9706 -2120
rect 9606 -2192 9706 -2154
rect 9764 -2120 9864 -2104
rect 9764 -2154 9780 -2120
rect 9848 -2154 9864 -2120
rect 9764 -2192 9864 -2154
rect 9922 -2120 10022 -2104
rect 9922 -2154 9938 -2120
rect 10006 -2154 10022 -2120
rect 9922 -2192 10022 -2154
rect 10080 -2120 10180 -2104
rect 10080 -2154 10096 -2120
rect 10164 -2154 10180 -2120
rect 10080 -2192 10180 -2154
rect 10238 -2120 10338 -2104
rect 10238 -2154 10254 -2120
rect 10322 -2154 10338 -2120
rect 10238 -2192 10338 -2154
rect 10396 -2120 10496 -2104
rect 10396 -2154 10412 -2120
rect 10480 -2154 10496 -2120
rect 10396 -2192 10496 -2154
rect 10554 -2120 10654 -2104
rect 10554 -2154 10570 -2120
rect 10638 -2154 10654 -2120
rect 10554 -2192 10654 -2154
rect 10712 -2120 10812 -2104
rect 10712 -2154 10728 -2120
rect 10796 -2154 10812 -2120
rect 10712 -2192 10812 -2154
rect 10870 -2120 10970 -2104
rect 10870 -2154 10886 -2120
rect 10954 -2154 10970 -2120
rect 10870 -2192 10970 -2154
rect 9448 -3030 9548 -2992
rect 9448 -3064 9464 -3030
rect 9532 -3064 9548 -3030
rect 9448 -3080 9548 -3064
rect 9606 -3030 9706 -2992
rect 9606 -3064 9622 -3030
rect 9690 -3064 9706 -3030
rect 9606 -3080 9706 -3064
rect 9764 -3030 9864 -2992
rect 9764 -3064 9780 -3030
rect 9848 -3064 9864 -3030
rect 9764 -3080 9864 -3064
rect 9922 -3030 10022 -2992
rect 9922 -3064 9938 -3030
rect 10006 -3064 10022 -3030
rect 9922 -3080 10022 -3064
rect 10080 -3030 10180 -2992
rect 10080 -3064 10096 -3030
rect 10164 -3064 10180 -3030
rect 10080 -3080 10180 -3064
rect 10238 -3030 10338 -2992
rect 10238 -3064 10254 -3030
rect 10322 -3064 10338 -3030
rect 10238 -3080 10338 -3064
rect 10396 -3030 10496 -2992
rect 10396 -3064 10412 -3030
rect 10480 -3064 10496 -3030
rect 10396 -3080 10496 -3064
rect 10554 -3030 10654 -2992
rect 10554 -3064 10570 -3030
rect 10638 -3064 10654 -3030
rect 10554 -3080 10654 -3064
rect 10712 -3030 10812 -2992
rect 10712 -3064 10728 -3030
rect 10796 -3064 10812 -3030
rect 10712 -3080 10812 -3064
rect 10870 -3030 10970 -2992
rect 10870 -3064 10886 -3030
rect 10954 -3064 10970 -3030
rect 10870 -3080 10970 -3064
rect 15053 -1992 15083 -1881
rect 14009 -2027 14035 -1997
rect 14165 -2011 14285 -1997
rect 14165 -2027 14203 -2011
rect 11480 -2088 11580 -2072
rect 11480 -2122 11496 -2088
rect 11564 -2122 11580 -2088
rect 11480 -2169 11580 -2122
rect 11480 -3016 11580 -2969
rect 11480 -3050 11496 -3016
rect 11564 -3050 11580 -3016
rect 11480 -3066 11580 -3050
rect 14187 -2045 14203 -2027
rect 14237 -2027 14285 -2011
rect 14485 -2027 14511 -1997
rect 14996 -2008 15083 -1992
rect 14237 -2045 14253 -2027
rect 14187 -2055 14253 -2045
rect 14996 -2042 15012 -2008
rect 15046 -2042 15083 -2008
rect 14187 -2160 14253 -2150
rect 14187 -2185 14203 -2160
rect 12686 -2268 12774 -2252
rect 12686 -3036 12702 -2268
rect 12736 -3036 12774 -2268
rect 12686 -3052 12774 -3036
rect 12874 -2268 12962 -2252
rect 12874 -3036 12912 -2268
rect 12946 -3036 12962 -2268
rect 12874 -3052 12962 -3036
rect 14009 -2215 14035 -2185
rect 14165 -2194 14203 -2185
rect 14237 -2185 14253 -2160
rect 14996 -2076 15083 -2042
rect 14996 -2110 15012 -2076
rect 15046 -2110 15083 -2076
rect 15125 -1959 15155 -1881
rect 15247 -1903 15277 -1881
rect 15247 -1919 15325 -1903
rect 15591 -1896 15621 -1881
rect 15247 -1933 15266 -1919
rect 15256 -1953 15266 -1933
rect 15300 -1953 15325 -1919
rect 15558 -1926 15621 -1896
rect 15558 -1949 15588 -1926
rect 15125 -1969 15214 -1959
rect 15125 -2003 15164 -1969
rect 15198 -2003 15214 -1969
rect 15125 -2037 15214 -2003
rect 15256 -1987 15325 -1953
rect 15256 -2021 15266 -1987
rect 15300 -2021 15325 -1987
rect 15534 -1965 15588 -1949
rect 15534 -1999 15544 -1965
rect 15578 -1999 15588 -1965
rect 15675 -1970 15705 -1881
rect 15534 -2015 15588 -1999
rect 15256 -2037 15325 -2021
rect 15125 -2071 15164 -2037
rect 15198 -2071 15214 -2037
rect 15125 -2092 15214 -2071
rect 14996 -2126 15083 -2110
rect 15053 -2163 15083 -2126
rect 15141 -2163 15171 -2092
rect 15295 -2119 15325 -2037
rect 15558 -2068 15588 -2015
rect 15630 -1980 15705 -1970
rect 15630 -2014 15646 -1980
rect 15680 -2014 15705 -1980
rect 15930 -2010 15960 -1881
rect 16025 -1903 16055 -1869
rect 16121 -1903 16151 -1869
rect 16002 -1919 16056 -1903
rect 16002 -1953 16012 -1919
rect 16046 -1953 16056 -1919
rect 16002 -1969 16056 -1953
rect 16098 -1913 16164 -1903
rect 16098 -1947 16114 -1913
rect 16148 -1947 16164 -1913
rect 16098 -1957 16164 -1947
rect 15630 -2024 15705 -2014
rect 15558 -2098 15621 -2068
rect 15591 -2113 15621 -2098
rect 15675 -2113 15705 -2024
rect 15843 -2026 15960 -2010
rect 15843 -2060 15853 -2026
rect 15887 -2046 15960 -2026
rect 16025 -1999 16056 -1969
rect 16025 -2029 16163 -1999
rect 15887 -2060 15972 -2046
rect 15843 -2076 15972 -2060
rect 14237 -2194 14285 -2185
rect 14165 -2215 14285 -2194
rect 14485 -2215 14511 -2185
rect 14187 -2267 14253 -2257
rect 14187 -2281 14203 -2267
rect 14009 -2311 14035 -2281
rect 14165 -2301 14203 -2281
rect 14237 -2281 14253 -2267
rect 15942 -2163 15972 -2076
rect 16018 -2081 16084 -2071
rect 16018 -2115 16034 -2081
rect 16068 -2115 16084 -2081
rect 16018 -2125 16084 -2115
rect 16034 -2163 16064 -2125
rect 16133 -2163 16163 -2029
rect 16287 -2039 16317 -1881
rect 16359 -1903 16389 -1881
rect 16359 -1919 16413 -1903
rect 16359 -1953 16369 -1919
rect 16403 -1953 16413 -1919
rect 16590 -1891 16620 -1869
rect 16590 -1907 16657 -1891
rect 16491 -1951 16521 -1925
rect 16359 -1969 16413 -1953
rect 16455 -1967 16521 -1951
rect 16590 -1941 16613 -1907
rect 16647 -1941 16657 -1907
rect 16590 -1957 16657 -1941
rect 16699 -1939 16729 -1869
rect 16795 -1913 16825 -1881
rect 16795 -1929 16897 -1913
rect 16699 -1955 16753 -1939
rect 16795 -1943 16853 -1929
rect 16273 -2055 16328 -2039
rect 16273 -2089 16283 -2055
rect 16317 -2089 16328 -2055
rect 16273 -2105 16328 -2089
rect 16273 -2163 16303 -2105
rect 16370 -2163 16400 -1969
rect 16455 -2001 16465 -1967
rect 16499 -2001 16521 -1967
rect 16699 -1987 16709 -1955
rect 16687 -1989 16709 -1987
rect 16743 -1989 16753 -1955
rect 16687 -1999 16753 -1989
rect 16455 -2017 16521 -2001
rect 16491 -2034 16521 -2017
rect 16666 -2005 16753 -1999
rect 16836 -1963 16853 -1943
rect 16887 -1963 16897 -1929
rect 16944 -1941 16974 -1881
rect 16836 -1979 16897 -1963
rect 16939 -1957 16993 -1941
rect 16666 -2017 16729 -2005
rect 16666 -2029 16716 -2017
rect 16491 -2064 16597 -2034
rect 16567 -2079 16597 -2064
rect 15053 -2273 15083 -2247
rect 15141 -2273 15171 -2247
rect 15295 -2273 15325 -2247
rect 15591 -2267 15621 -2241
rect 15675 -2267 15705 -2241
rect 16666 -2163 16696 -2029
rect 16738 -2081 16792 -2065
rect 16738 -2115 16748 -2081
rect 16782 -2115 16792 -2081
rect 16738 -2131 16792 -2115
rect 16752 -2163 16782 -2131
rect 16836 -2163 16866 -1979
rect 16939 -1991 16949 -1957
rect 16983 -1991 16993 -1957
rect 16939 -2007 16993 -1991
rect 16944 -2163 16974 -2007
rect 17035 -2049 17065 -1881
rect 17411 -1896 17441 -1881
rect 17400 -1926 17441 -1896
rect 17223 -1949 17253 -1927
rect 17400 -1949 17430 -1926
rect 17799 -1896 17829 -1881
rect 17766 -1926 17829 -1896
rect 17508 -1949 17538 -1927
rect 17766 -1949 17796 -1926
rect 17121 -1965 17430 -1949
rect 17121 -1999 17149 -1965
rect 17183 -1999 17430 -1965
rect 17121 -2015 17430 -1999
rect 17479 -1965 17538 -1949
rect 17479 -1999 17489 -1965
rect 17523 -1999 17538 -1965
rect 17479 -2015 17538 -1999
rect 17742 -1965 17796 -1949
rect 17742 -1999 17752 -1965
rect 17786 -1999 17796 -1965
rect 17883 -1970 17913 -1881
rect 17742 -2015 17796 -1999
rect 17192 -2047 17222 -2015
rect 17016 -2065 17070 -2049
rect 17016 -2099 17026 -2065
rect 17060 -2099 17070 -2065
rect 17016 -2115 17070 -2099
rect 17028 -2163 17058 -2115
rect 17400 -2053 17430 -2015
rect 17508 -2047 17538 -2015
rect 17400 -2083 17441 -2053
rect 17411 -2119 17441 -2083
rect 17766 -2068 17796 -2015
rect 17838 -1980 17913 -1970
rect 17838 -2014 17854 -1980
rect 17888 -2014 17913 -1980
rect 18138 -2010 18168 -1881
rect 18233 -1903 18263 -1869
rect 18329 -1903 18359 -1869
rect 18210 -1919 18264 -1903
rect 18210 -1953 18220 -1919
rect 18254 -1953 18264 -1919
rect 18210 -1969 18264 -1953
rect 18306 -1913 18372 -1903
rect 18306 -1947 18322 -1913
rect 18356 -1947 18372 -1913
rect 18306 -1957 18372 -1947
rect 17838 -2024 17913 -2014
rect 17766 -2098 17829 -2068
rect 17799 -2113 17829 -2098
rect 17883 -2113 17913 -2024
rect 18051 -2026 18168 -2010
rect 18051 -2060 18061 -2026
rect 18095 -2046 18168 -2026
rect 18233 -1999 18264 -1969
rect 18233 -2029 18371 -1999
rect 18095 -2060 18180 -2046
rect 18051 -2076 18180 -2060
rect 18150 -2163 18180 -2076
rect 18226 -2081 18292 -2071
rect 18226 -2115 18242 -2081
rect 18276 -2115 18292 -2081
rect 18226 -2125 18292 -2115
rect 18242 -2163 18272 -2125
rect 18341 -2163 18371 -2029
rect 18495 -2039 18525 -1881
rect 18567 -1903 18597 -1881
rect 18567 -1919 18621 -1903
rect 18567 -1953 18577 -1919
rect 18611 -1953 18621 -1919
rect 18798 -1891 18828 -1869
rect 18798 -1907 18865 -1891
rect 18699 -1951 18729 -1925
rect 18567 -1969 18621 -1953
rect 18663 -1967 18729 -1951
rect 18798 -1941 18821 -1907
rect 18855 -1941 18865 -1907
rect 18798 -1957 18865 -1941
rect 18907 -1939 18937 -1869
rect 19003 -1913 19033 -1881
rect 19003 -1929 19105 -1913
rect 18907 -1955 18961 -1939
rect 19003 -1943 19061 -1929
rect 18481 -2055 18536 -2039
rect 18481 -2089 18491 -2055
rect 18525 -2089 18536 -2055
rect 18481 -2105 18536 -2089
rect 18481 -2163 18511 -2105
rect 18578 -2163 18608 -1969
rect 18663 -2001 18673 -1967
rect 18707 -2001 18729 -1967
rect 18907 -1987 18917 -1955
rect 18895 -1989 18917 -1987
rect 18951 -1989 18961 -1955
rect 18895 -1999 18961 -1989
rect 18663 -2017 18729 -2001
rect 18699 -2034 18729 -2017
rect 18874 -2005 18961 -1999
rect 19044 -1963 19061 -1943
rect 19095 -1963 19105 -1929
rect 19152 -1941 19182 -1881
rect 19044 -1979 19105 -1963
rect 19147 -1957 19201 -1941
rect 18874 -2017 18937 -2005
rect 18874 -2029 18924 -2017
rect 18699 -2064 18805 -2034
rect 18775 -2079 18805 -2064
rect 15942 -2273 15972 -2247
rect 16034 -2273 16064 -2247
rect 16133 -2273 16163 -2247
rect 16273 -2273 16303 -2247
rect 16370 -2273 16400 -2247
rect 16567 -2273 16597 -2247
rect 16666 -2273 16696 -2247
rect 16752 -2273 16782 -2247
rect 16836 -2273 16866 -2247
rect 16944 -2273 16974 -2247
rect 17028 -2273 17058 -2247
rect 17192 -2273 17222 -2247
rect 17411 -2273 17441 -2247
rect 17508 -2273 17538 -2247
rect 17799 -2267 17829 -2241
rect 17883 -2267 17913 -2241
rect 18874 -2163 18904 -2029
rect 18946 -2081 19000 -2065
rect 18946 -2115 18956 -2081
rect 18990 -2115 19000 -2081
rect 18946 -2131 19000 -2115
rect 18960 -2163 18990 -2131
rect 19044 -2163 19074 -1979
rect 19147 -1991 19157 -1957
rect 19191 -1991 19201 -1957
rect 19147 -2007 19201 -1991
rect 19152 -2163 19182 -2007
rect 19243 -2049 19273 -1881
rect 19619 -1896 19649 -1881
rect 19608 -1926 19649 -1896
rect 19431 -1949 19461 -1927
rect 19608 -1949 19638 -1926
rect 20007 -1896 20037 -1881
rect 19974 -1926 20037 -1896
rect 19716 -1949 19746 -1927
rect 19974 -1949 20004 -1926
rect 19329 -1965 19638 -1949
rect 19329 -1999 19357 -1965
rect 19391 -1999 19638 -1965
rect 19329 -2015 19638 -1999
rect 19687 -1965 19746 -1949
rect 19687 -1999 19697 -1965
rect 19731 -1999 19746 -1965
rect 19687 -2015 19746 -1999
rect 19950 -1965 20004 -1949
rect 19950 -1999 19960 -1965
rect 19994 -1999 20004 -1965
rect 20091 -1970 20121 -1881
rect 19950 -2015 20004 -1999
rect 19400 -2047 19430 -2015
rect 19224 -2065 19278 -2049
rect 19224 -2099 19234 -2065
rect 19268 -2099 19278 -2065
rect 19224 -2115 19278 -2099
rect 19236 -2163 19266 -2115
rect 19608 -2053 19638 -2015
rect 19716 -2047 19746 -2015
rect 19608 -2083 19649 -2053
rect 19619 -2119 19649 -2083
rect 19974 -2068 20004 -2015
rect 20046 -1980 20121 -1970
rect 20046 -2014 20062 -1980
rect 20096 -2014 20121 -1980
rect 20346 -2010 20376 -1881
rect 20441 -1903 20471 -1869
rect 20537 -1903 20567 -1869
rect 20418 -1919 20472 -1903
rect 20418 -1953 20428 -1919
rect 20462 -1953 20472 -1919
rect 20418 -1969 20472 -1953
rect 20514 -1913 20580 -1903
rect 20514 -1947 20530 -1913
rect 20564 -1947 20580 -1913
rect 20514 -1957 20580 -1947
rect 20046 -2024 20121 -2014
rect 19974 -2098 20037 -2068
rect 20007 -2113 20037 -2098
rect 20091 -2113 20121 -2024
rect 20259 -2026 20376 -2010
rect 20259 -2060 20269 -2026
rect 20303 -2046 20376 -2026
rect 20441 -1999 20472 -1969
rect 20441 -2029 20579 -1999
rect 20303 -2060 20388 -2046
rect 20259 -2076 20388 -2060
rect 20358 -2163 20388 -2076
rect 20434 -2081 20500 -2071
rect 20434 -2115 20450 -2081
rect 20484 -2115 20500 -2081
rect 20434 -2125 20500 -2115
rect 20450 -2163 20480 -2125
rect 20549 -2163 20579 -2029
rect 20703 -2039 20733 -1881
rect 20775 -1903 20805 -1881
rect 20775 -1919 20829 -1903
rect 20775 -1953 20785 -1919
rect 20819 -1953 20829 -1919
rect 21006 -1891 21036 -1869
rect 21006 -1907 21073 -1891
rect 20907 -1951 20937 -1925
rect 20775 -1969 20829 -1953
rect 20871 -1967 20937 -1951
rect 21006 -1941 21029 -1907
rect 21063 -1941 21073 -1907
rect 21006 -1957 21073 -1941
rect 21115 -1939 21145 -1869
rect 21211 -1913 21241 -1881
rect 21211 -1929 21313 -1913
rect 21115 -1955 21169 -1939
rect 21211 -1943 21269 -1929
rect 20689 -2055 20744 -2039
rect 20689 -2089 20699 -2055
rect 20733 -2089 20744 -2055
rect 20689 -2105 20744 -2089
rect 20689 -2163 20719 -2105
rect 20786 -2163 20816 -1969
rect 20871 -2001 20881 -1967
rect 20915 -2001 20937 -1967
rect 21115 -1987 21125 -1955
rect 21103 -1989 21125 -1987
rect 21159 -1989 21169 -1955
rect 21103 -1999 21169 -1989
rect 20871 -2017 20937 -2001
rect 20907 -2034 20937 -2017
rect 21082 -2005 21169 -1999
rect 21252 -1963 21269 -1943
rect 21303 -1963 21313 -1929
rect 21360 -1941 21390 -1881
rect 21252 -1979 21313 -1963
rect 21355 -1957 21409 -1941
rect 21082 -2017 21145 -2005
rect 21082 -2029 21132 -2017
rect 20907 -2064 21013 -2034
rect 20983 -2079 21013 -2064
rect 18150 -2273 18180 -2247
rect 18242 -2273 18272 -2247
rect 18341 -2273 18371 -2247
rect 18481 -2273 18511 -2247
rect 18578 -2273 18608 -2247
rect 18775 -2273 18805 -2247
rect 18874 -2273 18904 -2247
rect 18960 -2273 18990 -2247
rect 19044 -2273 19074 -2247
rect 19152 -2273 19182 -2247
rect 19236 -2273 19266 -2247
rect 19400 -2273 19430 -2247
rect 19619 -2273 19649 -2247
rect 19716 -2273 19746 -2247
rect 20007 -2267 20037 -2241
rect 20091 -2267 20121 -2241
rect 21082 -2163 21112 -2029
rect 21154 -2081 21208 -2065
rect 21154 -2115 21164 -2081
rect 21198 -2115 21208 -2081
rect 21154 -2131 21208 -2115
rect 21168 -2163 21198 -2131
rect 21252 -2163 21282 -1979
rect 21355 -1991 21365 -1957
rect 21399 -1991 21409 -1957
rect 21355 -2007 21409 -1991
rect 21360 -2163 21390 -2007
rect 21451 -2049 21481 -1881
rect 21827 -1896 21857 -1881
rect 21816 -1926 21857 -1896
rect 21639 -1949 21669 -1927
rect 21816 -1949 21846 -1926
rect 21924 -1949 21954 -1927
rect 21537 -1965 21846 -1949
rect 21537 -1999 21565 -1965
rect 21599 -1999 21846 -1965
rect 21537 -2015 21846 -1999
rect 21895 -1965 21954 -1949
rect 21895 -1999 21905 -1965
rect 21939 -1999 21954 -1965
rect 21895 -2015 21954 -1999
rect 21608 -2047 21638 -2015
rect 21432 -2065 21486 -2049
rect 21432 -2099 21442 -2065
rect 21476 -2099 21486 -2065
rect 21432 -2115 21486 -2099
rect 21444 -2163 21474 -2115
rect 21816 -2053 21846 -2015
rect 21924 -2047 21954 -2015
rect 21816 -2083 21857 -2053
rect 21827 -2119 21857 -2083
rect 20358 -2273 20388 -2247
rect 20450 -2273 20480 -2247
rect 20549 -2273 20579 -2247
rect 20689 -2273 20719 -2247
rect 20786 -2273 20816 -2247
rect 20983 -2273 21013 -2247
rect 21082 -2273 21112 -2247
rect 21168 -2273 21198 -2247
rect 21252 -2273 21282 -2247
rect 21360 -2273 21390 -2247
rect 21444 -2273 21474 -2247
rect 21608 -2273 21638 -2247
rect 21827 -2273 21857 -2247
rect 21924 -2273 21954 -2247
rect 14237 -2301 14285 -2281
rect 14165 -2311 14285 -2301
rect 14485 -2311 14511 -2281
rect 14187 -2363 14253 -2353
rect 14187 -2374 14203 -2363
rect 14009 -2404 14035 -2374
rect 14165 -2397 14203 -2374
rect 14237 -2374 14253 -2363
rect 15053 -2341 15083 -2315
rect 15141 -2341 15171 -2315
rect 15295 -2341 15325 -2315
rect 14237 -2397 14285 -2374
rect 14165 -2404 14285 -2397
rect 14485 -2404 14511 -2374
rect 14187 -2407 14253 -2404
rect 15053 -2462 15083 -2425
rect 14187 -2554 14253 -2544
rect 14187 -2568 14203 -2554
rect 14009 -2598 14035 -2568
rect 14119 -2588 14203 -2568
rect 14237 -2568 14253 -2554
rect 14996 -2478 15083 -2462
rect 14996 -2512 15012 -2478
rect 15046 -2512 15083 -2478
rect 15141 -2496 15171 -2425
rect 15591 -2347 15621 -2321
rect 15675 -2347 15705 -2321
rect 15942 -2341 15972 -2315
rect 16034 -2341 16064 -2315
rect 16133 -2341 16163 -2315
rect 16273 -2341 16303 -2315
rect 16370 -2341 16400 -2315
rect 16567 -2341 16597 -2315
rect 16666 -2341 16696 -2315
rect 16752 -2341 16782 -2315
rect 16836 -2341 16866 -2315
rect 16944 -2341 16974 -2315
rect 17028 -2341 17058 -2315
rect 17192 -2341 17222 -2315
rect 17411 -2341 17441 -2315
rect 17508 -2341 17538 -2315
rect 14996 -2546 15083 -2512
rect 14237 -2588 14401 -2568
rect 14119 -2598 14401 -2588
rect 14485 -2598 14511 -2568
rect 14996 -2580 15012 -2546
rect 15046 -2580 15083 -2546
rect 14996 -2596 15083 -2580
rect 14187 -2650 14253 -2640
rect 14187 -2671 14203 -2650
rect 14009 -2701 14035 -2671
rect 14119 -2684 14203 -2671
rect 14237 -2684 14253 -2650
rect 14119 -2701 14253 -2684
rect 14312 -2671 14342 -2598
rect 14312 -2701 14357 -2671
rect 14485 -2701 14511 -2671
rect 15053 -2707 15083 -2596
rect 15125 -2517 15214 -2496
rect 15125 -2551 15164 -2517
rect 15198 -2551 15214 -2517
rect 15295 -2551 15325 -2469
rect 15591 -2490 15621 -2475
rect 15558 -2520 15621 -2490
rect 15125 -2585 15214 -2551
rect 15125 -2619 15164 -2585
rect 15198 -2619 15214 -2585
rect 15125 -2629 15214 -2619
rect 15256 -2567 15325 -2551
rect 15256 -2601 15266 -2567
rect 15300 -2601 15325 -2567
rect 15558 -2573 15588 -2520
rect 15675 -2564 15705 -2475
rect 15942 -2512 15972 -2425
rect 16034 -2463 16064 -2425
rect 15125 -2707 15155 -2629
rect 15256 -2635 15325 -2601
rect 15256 -2655 15266 -2635
rect 15247 -2669 15266 -2655
rect 15300 -2669 15325 -2635
rect 15534 -2589 15588 -2573
rect 15534 -2623 15544 -2589
rect 15578 -2623 15588 -2589
rect 15630 -2574 15705 -2564
rect 15630 -2608 15646 -2574
rect 15680 -2608 15705 -2574
rect 15843 -2528 15972 -2512
rect 16018 -2473 16084 -2463
rect 16018 -2507 16034 -2473
rect 16068 -2507 16084 -2473
rect 16018 -2517 16084 -2507
rect 15843 -2562 15853 -2528
rect 15887 -2542 15972 -2528
rect 15887 -2562 15960 -2542
rect 16133 -2559 16163 -2425
rect 16273 -2483 16303 -2425
rect 16273 -2499 16328 -2483
rect 16273 -2533 16283 -2499
rect 16317 -2533 16328 -2499
rect 16273 -2549 16328 -2533
rect 15843 -2578 15960 -2562
rect 15630 -2618 15705 -2608
rect 15534 -2639 15588 -2623
rect 15558 -2662 15588 -2639
rect 15247 -2685 15325 -2669
rect 15247 -2707 15277 -2685
rect 15558 -2692 15621 -2662
rect 14009 -2773 14035 -2743
rect 14119 -2773 14357 -2743
rect 14485 -2773 14511 -2743
rect 14187 -2786 14253 -2773
rect 14187 -2820 14203 -2786
rect 14237 -2820 14253 -2786
rect 14187 -2830 14253 -2820
rect 15591 -2707 15621 -2692
rect 15675 -2707 15705 -2618
rect 15930 -2707 15960 -2578
rect 16025 -2589 16163 -2559
rect 16025 -2619 16056 -2589
rect 16002 -2635 16056 -2619
rect 16002 -2669 16012 -2635
rect 16046 -2669 16056 -2635
rect 16002 -2685 16056 -2669
rect 16098 -2641 16164 -2631
rect 16098 -2675 16114 -2641
rect 16148 -2675 16164 -2641
rect 16098 -2685 16164 -2675
rect 16025 -2719 16055 -2685
rect 16121 -2719 16151 -2685
rect 16287 -2707 16317 -2549
rect 16370 -2619 16400 -2425
rect 16567 -2524 16597 -2509
rect 16491 -2554 16597 -2524
rect 16491 -2571 16521 -2554
rect 16455 -2587 16521 -2571
rect 16359 -2635 16413 -2619
rect 16359 -2669 16369 -2635
rect 16403 -2669 16413 -2635
rect 16455 -2621 16465 -2587
rect 16499 -2621 16521 -2587
rect 16666 -2559 16696 -2425
rect 16752 -2457 16782 -2425
rect 16738 -2473 16792 -2457
rect 16738 -2507 16748 -2473
rect 16782 -2507 16792 -2473
rect 16738 -2523 16792 -2507
rect 16666 -2571 16716 -2559
rect 16666 -2583 16729 -2571
rect 16666 -2589 16753 -2583
rect 16687 -2599 16753 -2589
rect 16687 -2601 16709 -2599
rect 16455 -2637 16521 -2621
rect 16491 -2663 16521 -2637
rect 16590 -2647 16657 -2631
rect 16359 -2685 16413 -2669
rect 16359 -2707 16389 -2685
rect 16590 -2681 16613 -2647
rect 16647 -2681 16657 -2647
rect 16590 -2697 16657 -2681
rect 16699 -2633 16709 -2601
rect 16743 -2633 16753 -2599
rect 16699 -2649 16753 -2633
rect 16836 -2609 16866 -2425
rect 16944 -2581 16974 -2425
rect 17028 -2473 17058 -2425
rect 17016 -2489 17070 -2473
rect 17016 -2523 17026 -2489
rect 17060 -2523 17070 -2489
rect 17016 -2539 17070 -2523
rect 16939 -2597 16993 -2581
rect 16836 -2625 16897 -2609
rect 16836 -2645 16853 -2625
rect 16590 -2719 16620 -2697
rect 16699 -2719 16729 -2649
rect 16795 -2659 16853 -2645
rect 16887 -2659 16897 -2625
rect 16939 -2631 16949 -2597
rect 16983 -2631 16993 -2597
rect 16939 -2647 16993 -2631
rect 16795 -2675 16897 -2659
rect 16795 -2707 16825 -2675
rect 16944 -2707 16974 -2647
rect 17035 -2707 17065 -2539
rect 17411 -2505 17441 -2469
rect 17400 -2535 17441 -2505
rect 17192 -2573 17222 -2541
rect 17400 -2573 17430 -2535
rect 17799 -2347 17829 -2321
rect 17883 -2347 17913 -2321
rect 18150 -2341 18180 -2315
rect 18242 -2341 18272 -2315
rect 18341 -2341 18371 -2315
rect 18481 -2341 18511 -2315
rect 18578 -2341 18608 -2315
rect 18775 -2341 18805 -2315
rect 18874 -2341 18904 -2315
rect 18960 -2341 18990 -2315
rect 19044 -2341 19074 -2315
rect 19152 -2341 19182 -2315
rect 19236 -2341 19266 -2315
rect 19400 -2341 19430 -2315
rect 19619 -2341 19649 -2315
rect 19716 -2341 19746 -2315
rect 17799 -2490 17829 -2475
rect 17766 -2520 17829 -2490
rect 17508 -2573 17538 -2541
rect 17766 -2573 17796 -2520
rect 17883 -2564 17913 -2475
rect 18150 -2512 18180 -2425
rect 18242 -2463 18272 -2425
rect 17121 -2589 17430 -2573
rect 17121 -2623 17149 -2589
rect 17183 -2623 17430 -2589
rect 17121 -2639 17430 -2623
rect 17479 -2589 17538 -2573
rect 17479 -2623 17489 -2589
rect 17523 -2623 17538 -2589
rect 17479 -2639 17538 -2623
rect 17742 -2589 17796 -2573
rect 17742 -2623 17752 -2589
rect 17786 -2623 17796 -2589
rect 17838 -2574 17913 -2564
rect 17838 -2608 17854 -2574
rect 17888 -2608 17913 -2574
rect 18051 -2528 18180 -2512
rect 18226 -2473 18292 -2463
rect 18226 -2507 18242 -2473
rect 18276 -2507 18292 -2473
rect 18226 -2517 18292 -2507
rect 18051 -2562 18061 -2528
rect 18095 -2542 18180 -2528
rect 18095 -2562 18168 -2542
rect 18341 -2559 18371 -2425
rect 18481 -2483 18511 -2425
rect 18481 -2499 18536 -2483
rect 18481 -2533 18491 -2499
rect 18525 -2533 18536 -2499
rect 18481 -2549 18536 -2533
rect 18051 -2578 18168 -2562
rect 17838 -2618 17913 -2608
rect 17742 -2639 17796 -2623
rect 17223 -2661 17253 -2639
rect 17400 -2662 17430 -2639
rect 17508 -2661 17538 -2639
rect 17400 -2692 17441 -2662
rect 17411 -2707 17441 -2692
rect 17766 -2662 17796 -2639
rect 17766 -2692 17829 -2662
rect 17799 -2707 17829 -2692
rect 17883 -2707 17913 -2618
rect 18138 -2707 18168 -2578
rect 18233 -2589 18371 -2559
rect 18233 -2619 18264 -2589
rect 18210 -2635 18264 -2619
rect 18210 -2669 18220 -2635
rect 18254 -2669 18264 -2635
rect 18210 -2685 18264 -2669
rect 18306 -2641 18372 -2631
rect 18306 -2675 18322 -2641
rect 18356 -2675 18372 -2641
rect 18306 -2685 18372 -2675
rect 18233 -2719 18263 -2685
rect 18329 -2719 18359 -2685
rect 18495 -2707 18525 -2549
rect 18578 -2619 18608 -2425
rect 18775 -2524 18805 -2509
rect 18699 -2554 18805 -2524
rect 18699 -2571 18729 -2554
rect 18663 -2587 18729 -2571
rect 18567 -2635 18621 -2619
rect 18567 -2669 18577 -2635
rect 18611 -2669 18621 -2635
rect 18663 -2621 18673 -2587
rect 18707 -2621 18729 -2587
rect 18874 -2559 18904 -2425
rect 18960 -2457 18990 -2425
rect 18946 -2473 19000 -2457
rect 18946 -2507 18956 -2473
rect 18990 -2507 19000 -2473
rect 18946 -2523 19000 -2507
rect 18874 -2571 18924 -2559
rect 18874 -2583 18937 -2571
rect 18874 -2589 18961 -2583
rect 18895 -2599 18961 -2589
rect 18895 -2601 18917 -2599
rect 18663 -2637 18729 -2621
rect 18699 -2663 18729 -2637
rect 18798 -2647 18865 -2631
rect 18567 -2685 18621 -2669
rect 18567 -2707 18597 -2685
rect 18798 -2681 18821 -2647
rect 18855 -2681 18865 -2647
rect 18798 -2697 18865 -2681
rect 18907 -2633 18917 -2601
rect 18951 -2633 18961 -2599
rect 18907 -2649 18961 -2633
rect 19044 -2609 19074 -2425
rect 19152 -2581 19182 -2425
rect 19236 -2473 19266 -2425
rect 19224 -2489 19278 -2473
rect 19224 -2523 19234 -2489
rect 19268 -2523 19278 -2489
rect 19224 -2539 19278 -2523
rect 19147 -2597 19201 -2581
rect 19044 -2625 19105 -2609
rect 19044 -2645 19061 -2625
rect 18798 -2719 18828 -2697
rect 18907 -2719 18937 -2649
rect 19003 -2659 19061 -2645
rect 19095 -2659 19105 -2625
rect 19147 -2631 19157 -2597
rect 19191 -2631 19201 -2597
rect 19147 -2647 19201 -2631
rect 19003 -2675 19105 -2659
rect 19003 -2707 19033 -2675
rect 19152 -2707 19182 -2647
rect 19243 -2707 19273 -2539
rect 19619 -2505 19649 -2469
rect 19608 -2535 19649 -2505
rect 19400 -2573 19430 -2541
rect 19608 -2573 19638 -2535
rect 20007 -2347 20037 -2321
rect 20091 -2347 20121 -2321
rect 20358 -2341 20388 -2315
rect 20450 -2341 20480 -2315
rect 20549 -2341 20579 -2315
rect 20689 -2341 20719 -2315
rect 20786 -2341 20816 -2315
rect 20983 -2341 21013 -2315
rect 21082 -2341 21112 -2315
rect 21168 -2341 21198 -2315
rect 21252 -2341 21282 -2315
rect 21360 -2341 21390 -2315
rect 21444 -2341 21474 -2315
rect 21608 -2341 21638 -2315
rect 21827 -2341 21857 -2315
rect 21924 -2341 21954 -2315
rect 20007 -2490 20037 -2475
rect 19974 -2520 20037 -2490
rect 19716 -2573 19746 -2541
rect 19974 -2573 20004 -2520
rect 20091 -2564 20121 -2475
rect 20358 -2512 20388 -2425
rect 20450 -2463 20480 -2425
rect 19329 -2589 19638 -2573
rect 19329 -2623 19357 -2589
rect 19391 -2623 19638 -2589
rect 19329 -2639 19638 -2623
rect 19687 -2589 19746 -2573
rect 19687 -2623 19697 -2589
rect 19731 -2623 19746 -2589
rect 19687 -2639 19746 -2623
rect 19950 -2589 20004 -2573
rect 19950 -2623 19960 -2589
rect 19994 -2623 20004 -2589
rect 20046 -2574 20121 -2564
rect 20046 -2608 20062 -2574
rect 20096 -2608 20121 -2574
rect 20259 -2528 20388 -2512
rect 20434 -2473 20500 -2463
rect 20434 -2507 20450 -2473
rect 20484 -2507 20500 -2473
rect 20434 -2517 20500 -2507
rect 20259 -2562 20269 -2528
rect 20303 -2542 20388 -2528
rect 20303 -2562 20376 -2542
rect 20549 -2559 20579 -2425
rect 20689 -2483 20719 -2425
rect 20689 -2499 20744 -2483
rect 20689 -2533 20699 -2499
rect 20733 -2533 20744 -2499
rect 20689 -2549 20744 -2533
rect 20259 -2578 20376 -2562
rect 20046 -2618 20121 -2608
rect 19950 -2639 20004 -2623
rect 19431 -2661 19461 -2639
rect 19608 -2662 19638 -2639
rect 19716 -2661 19746 -2639
rect 19608 -2692 19649 -2662
rect 19619 -2707 19649 -2692
rect 19974 -2662 20004 -2639
rect 19974 -2692 20037 -2662
rect 20007 -2707 20037 -2692
rect 20091 -2707 20121 -2618
rect 20346 -2707 20376 -2578
rect 20441 -2589 20579 -2559
rect 20441 -2619 20472 -2589
rect 20418 -2635 20472 -2619
rect 20418 -2669 20428 -2635
rect 20462 -2669 20472 -2635
rect 20418 -2685 20472 -2669
rect 20514 -2641 20580 -2631
rect 20514 -2675 20530 -2641
rect 20564 -2675 20580 -2641
rect 20514 -2685 20580 -2675
rect 20441 -2719 20471 -2685
rect 20537 -2719 20567 -2685
rect 20703 -2707 20733 -2549
rect 20786 -2619 20816 -2425
rect 20983 -2524 21013 -2509
rect 20907 -2554 21013 -2524
rect 20907 -2571 20937 -2554
rect 20871 -2587 20937 -2571
rect 20775 -2635 20829 -2619
rect 20775 -2669 20785 -2635
rect 20819 -2669 20829 -2635
rect 20871 -2621 20881 -2587
rect 20915 -2621 20937 -2587
rect 21082 -2559 21112 -2425
rect 21168 -2457 21198 -2425
rect 21154 -2473 21208 -2457
rect 21154 -2507 21164 -2473
rect 21198 -2507 21208 -2473
rect 21154 -2523 21208 -2507
rect 21082 -2571 21132 -2559
rect 21082 -2583 21145 -2571
rect 21082 -2589 21169 -2583
rect 21103 -2599 21169 -2589
rect 21103 -2601 21125 -2599
rect 20871 -2637 20937 -2621
rect 20907 -2663 20937 -2637
rect 21006 -2647 21073 -2631
rect 20775 -2685 20829 -2669
rect 20775 -2707 20805 -2685
rect 21006 -2681 21029 -2647
rect 21063 -2681 21073 -2647
rect 21006 -2697 21073 -2681
rect 21115 -2633 21125 -2601
rect 21159 -2633 21169 -2599
rect 21115 -2649 21169 -2633
rect 21252 -2609 21282 -2425
rect 21360 -2581 21390 -2425
rect 21444 -2473 21474 -2425
rect 21432 -2489 21486 -2473
rect 21432 -2523 21442 -2489
rect 21476 -2523 21486 -2489
rect 21432 -2539 21486 -2523
rect 21355 -2597 21409 -2581
rect 21252 -2625 21313 -2609
rect 21252 -2645 21269 -2625
rect 21006 -2719 21036 -2697
rect 21115 -2719 21145 -2649
rect 21211 -2659 21269 -2645
rect 21303 -2659 21313 -2625
rect 21355 -2631 21365 -2597
rect 21399 -2631 21409 -2597
rect 21355 -2647 21409 -2631
rect 21211 -2675 21313 -2659
rect 21211 -2707 21241 -2675
rect 21360 -2707 21390 -2647
rect 21451 -2707 21481 -2539
rect 21827 -2505 21857 -2469
rect 21816 -2535 21857 -2505
rect 21608 -2573 21638 -2541
rect 21816 -2573 21846 -2535
rect 21924 -2573 21954 -2541
rect 21537 -2589 21846 -2573
rect 21537 -2623 21565 -2589
rect 21599 -2623 21846 -2589
rect 21537 -2639 21846 -2623
rect 21895 -2589 21954 -2573
rect 21895 -2623 21905 -2589
rect 21939 -2623 21954 -2589
rect 21895 -2639 21954 -2623
rect 21639 -2661 21669 -2639
rect 21816 -2662 21846 -2639
rect 21924 -2661 21954 -2639
rect 21816 -2692 21857 -2662
rect 21827 -2707 21857 -2692
rect 15053 -2817 15083 -2791
rect 15125 -2817 15155 -2791
rect 15247 -2817 15277 -2791
rect 15591 -2817 15621 -2791
rect 15675 -2817 15705 -2791
rect 15930 -2817 15960 -2791
rect 16025 -2817 16055 -2791
rect 16121 -2817 16151 -2791
rect 16287 -2817 16317 -2791
rect 16359 -2817 16389 -2791
rect 16491 -2817 16521 -2791
rect 16590 -2817 16620 -2791
rect 16699 -2817 16729 -2791
rect 16795 -2817 16825 -2791
rect 16944 -2817 16974 -2791
rect 17035 -2817 17065 -2791
rect 17223 -2817 17253 -2791
rect 17411 -2817 17441 -2791
rect 17508 -2817 17538 -2791
rect 17799 -2817 17829 -2791
rect 17883 -2817 17913 -2791
rect 18138 -2817 18168 -2791
rect 18233 -2817 18263 -2791
rect 18329 -2817 18359 -2791
rect 18495 -2817 18525 -2791
rect 18567 -2817 18597 -2791
rect 18699 -2817 18729 -2791
rect 18798 -2817 18828 -2791
rect 18907 -2817 18937 -2791
rect 19003 -2817 19033 -2791
rect 19152 -2817 19182 -2791
rect 19243 -2817 19273 -2791
rect 19431 -2817 19461 -2791
rect 19619 -2817 19649 -2791
rect 19716 -2817 19746 -2791
rect 20007 -2817 20037 -2791
rect 20091 -2817 20121 -2791
rect 20346 -2817 20376 -2791
rect 20441 -2817 20471 -2791
rect 20537 -2817 20567 -2791
rect 20703 -2817 20733 -2791
rect 20775 -2817 20805 -2791
rect 20907 -2817 20937 -2791
rect 21006 -2817 21036 -2791
rect 21115 -2817 21145 -2791
rect 21211 -2817 21241 -2791
rect 21360 -2817 21390 -2791
rect 21451 -2817 21481 -2791
rect 21639 -2817 21669 -2791
rect 21827 -2817 21857 -2791
rect 21924 -2817 21954 -2791
rect 15156 -3094 15956 -3078
rect 15156 -3128 15172 -3094
rect 15940 -3128 15956 -3094
rect 15156 -3166 15956 -3128
rect 15156 -3304 15956 -3266
rect 15156 -3338 15172 -3304
rect 15940 -3338 15956 -3304
rect 15156 -3354 15956 -3338
rect 2728 -4054 2828 -4038
rect 2728 -4088 2744 -4054
rect 2812 -4088 2828 -4054
rect 2728 -4126 2828 -4088
rect 2886 -4054 2986 -4038
rect 2886 -4088 2902 -4054
rect 2970 -4088 2986 -4054
rect 2886 -4126 2986 -4088
rect 2728 -4764 2828 -4726
rect 2728 -4798 2744 -4764
rect 2812 -4798 2828 -4764
rect 2728 -4814 2828 -4798
rect 2886 -4764 2986 -4726
rect 2886 -4798 2902 -4764
rect 2970 -4798 2986 -4764
rect 2886 -4814 2986 -4798
rect 3434 -4054 3534 -4038
rect 3434 -4088 3450 -4054
rect 3518 -4088 3534 -4054
rect 3434 -4126 3534 -4088
rect 3592 -4054 3692 -4038
rect 3592 -4088 3608 -4054
rect 3676 -4088 3692 -4054
rect 3592 -4126 3692 -4088
rect 3434 -4764 3534 -4726
rect 3434 -4798 3450 -4764
rect 3518 -4798 3534 -4764
rect 3434 -4814 3534 -4798
rect 3592 -4764 3692 -4726
rect 3592 -4798 3608 -4764
rect 3676 -4798 3692 -4764
rect 3592 -4814 3692 -4798
rect 4644 -4054 4744 -4038
rect 4644 -4088 4660 -4054
rect 4728 -4088 4744 -4054
rect 4644 -4126 4744 -4088
rect 4802 -4054 4902 -4038
rect 4802 -4088 4818 -4054
rect 4886 -4088 4902 -4054
rect 4802 -4126 4902 -4088
rect 4644 -4764 4744 -4726
rect 4644 -4798 4660 -4764
rect 4728 -4798 4744 -4764
rect 4644 -4814 4744 -4798
rect 4802 -4764 4902 -4726
rect 4802 -4798 4818 -4764
rect 4886 -4798 4902 -4764
rect 4802 -4814 4902 -4798
rect 5350 -4054 5450 -4038
rect 5350 -4088 5366 -4054
rect 5434 -4088 5450 -4054
rect 5350 -4126 5450 -4088
rect 5508 -4054 5608 -4038
rect 5508 -4088 5524 -4054
rect 5592 -4088 5608 -4054
rect 5508 -4126 5608 -4088
rect 5350 -4764 5450 -4726
rect 5350 -4798 5366 -4764
rect 5434 -4798 5450 -4764
rect 5350 -4814 5450 -4798
rect 5508 -4764 5608 -4726
rect 5508 -4798 5524 -4764
rect 5592 -4798 5608 -4764
rect 5508 -4814 5608 -4798
rect 2810 -5348 3610 -5332
rect 2810 -5382 2826 -5348
rect 3594 -5382 3610 -5348
rect 2810 -5429 3610 -5382
rect 2810 -5676 3610 -5629
rect 2810 -5710 2826 -5676
rect 3594 -5710 3610 -5676
rect 2810 -5726 3610 -5710
rect 2810 -5952 3610 -5936
rect 2810 -5986 2826 -5952
rect 3594 -5986 3610 -5952
rect 2810 -6033 3610 -5986
rect 2810 -6280 3610 -6233
rect 2810 -6314 2826 -6280
rect 3594 -6314 3610 -6280
rect 2810 -6330 3610 -6314
rect 4726 -5348 5526 -5332
rect 4726 -5382 4742 -5348
rect 5510 -5382 5526 -5348
rect 4726 -5429 5526 -5382
rect 4726 -5676 5526 -5629
rect 4726 -5710 4742 -5676
rect 5510 -5710 5526 -5676
rect 4726 -5726 5526 -5710
rect 4726 -5952 5526 -5936
rect 4726 -5986 4742 -5952
rect 5510 -5986 5526 -5952
rect 4726 -6033 5526 -5986
rect 4726 -6280 5526 -6233
rect 4726 -6314 4742 -6280
rect 5510 -6314 5526 -6280
rect 4726 -6330 5526 -6314
rect 2497 -7181 2597 -7165
rect 2497 -7215 2513 -7181
rect 2581 -7215 2597 -7181
rect 2497 -7253 2597 -7215
rect 2655 -7181 2755 -7165
rect 2655 -7215 2671 -7181
rect 2739 -7215 2755 -7181
rect 2655 -7253 2755 -7215
rect 2813 -7181 2913 -7165
rect 2813 -7215 2829 -7181
rect 2897 -7215 2913 -7181
rect 2813 -7253 2913 -7215
rect 2971 -7181 3071 -7165
rect 2971 -7215 2987 -7181
rect 3055 -7215 3071 -7181
rect 2971 -7253 3071 -7215
rect 3129 -7181 3229 -7165
rect 3129 -7215 3145 -7181
rect 3213 -7215 3229 -7181
rect 3129 -7253 3229 -7215
rect 2497 -8091 2597 -8053
rect 2497 -8125 2513 -8091
rect 2581 -8125 2597 -8091
rect 2497 -8141 2597 -8125
rect 2655 -8091 2755 -8053
rect 2655 -8125 2671 -8091
rect 2739 -8125 2755 -8091
rect 2655 -8141 2755 -8125
rect 2813 -8091 2913 -8053
rect 2813 -8125 2829 -8091
rect 2897 -8125 2913 -8091
rect 2813 -8141 2913 -8125
rect 2971 -8091 3071 -8053
rect 2971 -8125 2987 -8091
rect 3055 -8125 3071 -8091
rect 2971 -8141 3071 -8125
rect 3129 -8091 3229 -8053
rect 3129 -8125 3145 -8091
rect 3213 -8125 3229 -8091
rect 3129 -8141 3229 -8125
rect 3872 -7174 3972 -7158
rect 3872 -7208 3888 -7174
rect 3956 -7208 3972 -7174
rect 3872 -7255 3972 -7208
rect 4030 -7174 4130 -7158
rect 4030 -7208 4046 -7174
rect 4114 -7208 4130 -7174
rect 4030 -7255 4130 -7208
rect 4188 -7174 4288 -7158
rect 4188 -7208 4204 -7174
rect 4272 -7208 4288 -7174
rect 4188 -7255 4288 -7208
rect 4346 -7174 4446 -7158
rect 4346 -7208 4362 -7174
rect 4430 -7208 4446 -7174
rect 4346 -7255 4446 -7208
rect 4504 -7174 4604 -7158
rect 4504 -7208 4520 -7174
rect 4588 -7208 4604 -7174
rect 4504 -7255 4604 -7208
rect 3872 -8102 3972 -8055
rect 3872 -8136 3888 -8102
rect 3956 -8136 3972 -8102
rect 3872 -8152 3972 -8136
rect 4030 -8102 4130 -8055
rect 4030 -8136 4046 -8102
rect 4114 -8136 4130 -8102
rect 4030 -8152 4130 -8136
rect 4188 -8102 4288 -8055
rect 4188 -8136 4204 -8102
rect 4272 -8136 4288 -8102
rect 4188 -8152 4288 -8136
rect 4346 -8102 4446 -8055
rect 4346 -8136 4362 -8102
rect 4430 -8136 4446 -8102
rect 4346 -8152 4446 -8136
rect 4504 -8102 4604 -8055
rect 4504 -8136 4520 -8102
rect 4588 -8136 4604 -8102
rect 4504 -8152 4604 -8136
rect 10658 -4886 11058 -4870
rect 10658 -4920 10674 -4886
rect 11042 -4920 11058 -4886
rect 10658 -4958 11058 -4920
rect 11236 -4886 11636 -4870
rect 11236 -4920 11252 -4886
rect 11620 -4920 11636 -4886
rect 11236 -4958 11636 -4920
rect 11814 -4886 12214 -4870
rect 11814 -4920 11830 -4886
rect 12198 -4920 12214 -4886
rect 11814 -4958 12214 -4920
rect 12392 -4886 12792 -4870
rect 12392 -4920 12408 -4886
rect 12776 -4920 12792 -4886
rect 12392 -4958 12792 -4920
rect 12970 -4886 13370 -4870
rect 12970 -4920 12986 -4886
rect 13354 -4920 13370 -4886
rect 12970 -4958 13370 -4920
rect 13548 -4886 13948 -4870
rect 13548 -4920 13564 -4886
rect 13932 -4920 13948 -4886
rect 13548 -4958 13948 -4920
rect 14126 -4886 14526 -4870
rect 14126 -4920 14142 -4886
rect 14510 -4920 14526 -4886
rect 14126 -4958 14526 -4920
rect 14704 -4886 15104 -4870
rect 14704 -4920 14720 -4886
rect 15088 -4920 15104 -4886
rect 14704 -4958 15104 -4920
rect 10658 -5396 11058 -5358
rect 10658 -5430 10674 -5396
rect 11042 -5430 11058 -5396
rect 10658 -5446 11058 -5430
rect 11236 -5396 11636 -5358
rect 11236 -5430 11252 -5396
rect 11620 -5430 11636 -5396
rect 11236 -5446 11636 -5430
rect 11814 -5396 12214 -5358
rect 11814 -5430 11830 -5396
rect 12198 -5430 12214 -5396
rect 11814 -5446 12214 -5430
rect 12392 -5396 12792 -5358
rect 12392 -5430 12408 -5396
rect 12776 -5430 12792 -5396
rect 12392 -5446 12792 -5430
rect 12970 -5396 13370 -5358
rect 12970 -5430 12986 -5396
rect 13354 -5430 13370 -5396
rect 12970 -5446 13370 -5430
rect 13548 -5396 13948 -5358
rect 13548 -5430 13564 -5396
rect 13932 -5430 13948 -5396
rect 13548 -5446 13948 -5430
rect 14126 -5396 14526 -5358
rect 14126 -5430 14142 -5396
rect 14510 -5430 14526 -5396
rect 14126 -5446 14526 -5430
rect 14704 -5396 15104 -5358
rect 14704 -5430 14720 -5396
rect 15088 -5430 15104 -5396
rect 14704 -5446 15104 -5430
rect 16260 -4666 16660 -4650
rect 16260 -4700 16276 -4666
rect 16644 -4700 16660 -4666
rect 16260 -4738 16660 -4700
rect 16718 -4666 17118 -4650
rect 16718 -4700 16734 -4666
rect 17102 -4700 17118 -4666
rect 16718 -4738 17118 -4700
rect 17176 -4666 17576 -4650
rect 17176 -4700 17192 -4666
rect 17560 -4700 17576 -4666
rect 17176 -4738 17576 -4700
rect 17634 -4666 18034 -4650
rect 17634 -4700 17650 -4666
rect 18018 -4700 18034 -4666
rect 17634 -4738 18034 -4700
rect 16260 -5576 16660 -5538
rect 16260 -5610 16276 -5576
rect 16644 -5610 16660 -5576
rect 16260 -5626 16660 -5610
rect 16718 -5576 17118 -5538
rect 16718 -5610 16734 -5576
rect 17102 -5610 17118 -5576
rect 16718 -5626 17118 -5610
rect 17176 -5576 17576 -5538
rect 17176 -5610 17192 -5576
rect 17560 -5610 17576 -5576
rect 17176 -5626 17576 -5610
rect 17634 -5576 18034 -5538
rect 17634 -5610 17650 -5576
rect 18018 -5610 18034 -5576
rect 17634 -5626 18034 -5610
rect 18948 -5462 20548 -5446
rect 18948 -5496 18964 -5462
rect 20532 -5496 20548 -5462
rect 18948 -5534 20548 -5496
rect 18948 -5672 20548 -5634
rect 18948 -5706 18964 -5672
rect 20532 -5706 20548 -5672
rect 18948 -5722 20548 -5706
rect 21412 -5334 21612 -5318
rect 21412 -5368 21428 -5334
rect 21596 -5368 21612 -5334
rect 21412 -5406 21612 -5368
rect 21670 -5334 21870 -5318
rect 21670 -5368 21686 -5334
rect 21854 -5368 21870 -5334
rect 21670 -5406 21870 -5368
rect 21412 -5544 21612 -5506
rect 21412 -5578 21428 -5544
rect 21596 -5578 21612 -5544
rect 21412 -5616 21612 -5578
rect 21670 -5544 21870 -5506
rect 21670 -5578 21686 -5544
rect 21854 -5578 21870 -5544
rect 21670 -5616 21870 -5578
rect 10682 -5908 11082 -5892
rect 10682 -5942 10698 -5908
rect 11066 -5942 11082 -5908
rect 10682 -5989 11082 -5942
rect 11254 -5908 11654 -5892
rect 11254 -5942 11270 -5908
rect 11638 -5942 11654 -5908
rect 11254 -5989 11654 -5942
rect 11826 -5908 12226 -5892
rect 11826 -5942 11842 -5908
rect 12210 -5942 12226 -5908
rect 11826 -5989 12226 -5942
rect 12398 -5908 12798 -5892
rect 12398 -5942 12414 -5908
rect 12782 -5942 12798 -5908
rect 12398 -5989 12798 -5942
rect 12970 -5908 13370 -5892
rect 12970 -5942 12986 -5908
rect 13354 -5942 13370 -5908
rect 12970 -5989 13370 -5942
rect 13542 -5908 13942 -5892
rect 13542 -5942 13558 -5908
rect 13926 -5942 13942 -5908
rect 13542 -5989 13942 -5942
rect 14114 -5908 14514 -5892
rect 14114 -5942 14130 -5908
rect 14498 -5942 14514 -5908
rect 14114 -5989 14514 -5942
rect 14686 -5908 15086 -5892
rect 14686 -5942 14702 -5908
rect 15070 -5942 15086 -5908
rect 14686 -5989 15086 -5942
rect 21412 -5754 21612 -5716
rect 21412 -5788 21428 -5754
rect 21596 -5788 21612 -5754
rect 21412 -5804 21612 -5788
rect 21670 -5754 21870 -5716
rect 21670 -5788 21686 -5754
rect 21854 -5788 21870 -5754
rect 21670 -5804 21870 -5788
rect 23346 -5464 23434 -5448
rect 23346 -5632 23362 -5464
rect 23396 -5632 23434 -5464
rect 23346 -5648 23434 -5632
rect 23584 -5464 23672 -5448
rect 23584 -5632 23622 -5464
rect 23656 -5632 23672 -5464
rect 23584 -5648 23672 -5632
rect 10682 -6436 11082 -6389
rect 10682 -6470 10698 -6436
rect 11066 -6470 11082 -6436
rect 10682 -6517 11082 -6470
rect 11254 -6436 11654 -6389
rect 11254 -6470 11270 -6436
rect 11638 -6470 11654 -6436
rect 11254 -6517 11654 -6470
rect 11826 -6436 12226 -6389
rect 11826 -6470 11842 -6436
rect 12210 -6470 12226 -6436
rect 11826 -6517 12226 -6470
rect 12398 -6436 12798 -6389
rect 12398 -6470 12414 -6436
rect 12782 -6470 12798 -6436
rect 12398 -6517 12798 -6470
rect 12970 -6436 13370 -6389
rect 12970 -6470 12986 -6436
rect 13354 -6470 13370 -6436
rect 12970 -6517 13370 -6470
rect 13542 -6436 13942 -6389
rect 13542 -6470 13558 -6436
rect 13926 -6470 13942 -6436
rect 13542 -6517 13942 -6470
rect 14114 -6436 14514 -6389
rect 14114 -6470 14130 -6436
rect 14498 -6470 14514 -6436
rect 14114 -6517 14514 -6470
rect 14686 -6436 15086 -6389
rect 14686 -6470 14702 -6436
rect 15070 -6470 15086 -6436
rect 14686 -6517 15086 -6470
rect 10682 -6964 11082 -6917
rect 10682 -6998 10698 -6964
rect 11066 -6998 11082 -6964
rect 10682 -7014 11082 -6998
rect 11254 -6964 11654 -6917
rect 11254 -6998 11270 -6964
rect 11638 -6998 11654 -6964
rect 11254 -7014 11654 -6998
rect 11826 -6964 12226 -6917
rect 11826 -6998 11842 -6964
rect 12210 -6998 12226 -6964
rect 11826 -7014 12226 -6998
rect 12398 -6964 12798 -6917
rect 12398 -6998 12414 -6964
rect 12782 -6998 12798 -6964
rect 12398 -7014 12798 -6998
rect 12970 -6964 13370 -6917
rect 12970 -6998 12986 -6964
rect 13354 -6998 13370 -6964
rect 12970 -7014 13370 -6998
rect 13542 -6964 13942 -6917
rect 13542 -6998 13558 -6964
rect 13926 -6998 13942 -6964
rect 13542 -7014 13942 -6998
rect 14114 -6964 14514 -6917
rect 14114 -6998 14130 -6964
rect 14498 -6998 14514 -6964
rect 14114 -7014 14514 -6998
rect 14686 -6964 15086 -6917
rect 14686 -6998 14702 -6964
rect 15070 -6998 15086 -6964
rect 14686 -7014 15086 -6998
rect 16260 -6016 16660 -6000
rect 16260 -6050 16276 -6016
rect 16644 -6050 16660 -6016
rect 16260 -6097 16660 -6050
rect 16718 -6016 17118 -6000
rect 16718 -6050 16734 -6016
rect 17102 -6050 17118 -6016
rect 16718 -6097 17118 -6050
rect 17176 -6016 17576 -6000
rect 17176 -6050 17192 -6016
rect 17560 -6050 17576 -6016
rect 17176 -6097 17576 -6050
rect 17634 -6016 18034 -6000
rect 17634 -6050 17650 -6016
rect 18018 -6050 18034 -6016
rect 17634 -6097 18034 -6050
rect 16260 -6944 16660 -6897
rect 16260 -6978 16276 -6944
rect 16644 -6978 16660 -6944
rect 16260 -6994 16660 -6978
rect 16718 -6944 17118 -6897
rect 16718 -6978 16734 -6944
rect 17102 -6978 17118 -6944
rect 16718 -6994 17118 -6978
rect 17176 -6944 17576 -6897
rect 17176 -6978 17192 -6944
rect 17560 -6978 17576 -6944
rect 17176 -6994 17576 -6978
rect 17634 -6944 18034 -6897
rect 17634 -6978 17650 -6944
rect 18018 -6978 18034 -6944
rect 17634 -6994 18034 -6978
rect 18928 -6466 20528 -6450
rect 18928 -6500 18944 -6466
rect 20512 -6500 20528 -6466
rect 18928 -6547 20528 -6500
rect 18928 -6694 20528 -6647
rect 18928 -6728 18944 -6694
rect 20512 -6728 20528 -6694
rect 18928 -6744 20528 -6728
rect 21412 -6330 21612 -6314
rect 21412 -6364 21428 -6330
rect 21596 -6364 21612 -6330
rect 21412 -6411 21612 -6364
rect 21670 -6330 21870 -6314
rect 21670 -6364 21686 -6330
rect 21854 -6364 21870 -6330
rect 21670 -6411 21870 -6364
rect 21412 -6558 21612 -6511
rect 21412 -6592 21428 -6558
rect 21596 -6592 21612 -6558
rect 21412 -6639 21612 -6592
rect 21670 -6558 21870 -6511
rect 21670 -6592 21686 -6558
rect 21854 -6592 21870 -6558
rect 21670 -6639 21870 -6592
rect 21412 -6786 21612 -6739
rect 21412 -6820 21428 -6786
rect 21596 -6820 21612 -6786
rect 21412 -6836 21612 -6820
rect 21670 -6786 21870 -6739
rect 21670 -6820 21686 -6786
rect 21854 -6820 21870 -6786
rect 21670 -6836 21870 -6820
rect 23034 -6466 23131 -6450
rect 23034 -6634 23050 -6466
rect 23084 -6634 23131 -6466
rect 23034 -6650 23131 -6634
rect 23931 -6466 24028 -6450
rect 23931 -6634 23978 -6466
rect 24012 -6634 24028 -6466
rect 23931 -6650 24028 -6634
rect 9120 -7762 9208 -7746
rect 9120 -9330 9136 -7762
rect 9170 -9330 9208 -7762
rect 9120 -9346 9208 -9330
rect 9308 -7762 9396 -7746
rect 9308 -9330 9346 -7762
rect 9380 -9330 9396 -7762
rect 9308 -9346 9396 -9330
rect 9700 -7496 9797 -7480
rect 9700 -9064 9716 -7496
rect 9750 -9064 9797 -7496
rect 9700 -9080 9797 -9064
rect 9897 -7496 9994 -7480
rect 9897 -9064 9944 -7496
rect 9978 -9064 9994 -7496
rect 9897 -9080 9994 -9064
rect 7326 -12178 7526 -12162
rect 7326 -12212 7342 -12178
rect 7510 -12212 7526 -12178
rect 7326 -12250 7526 -12212
rect 7326 -12488 7526 -12450
rect 7326 -12522 7342 -12488
rect 7510 -12522 7526 -12488
rect 7326 -12538 7526 -12522
rect 8268 -12238 9868 -12222
rect 8268 -12272 8284 -12238
rect 9852 -12272 9868 -12238
rect 8268 -12310 9868 -12272
rect 9926 -12238 11526 -12222
rect 9926 -12272 9942 -12238
rect 11510 -12272 11526 -12238
rect 9926 -12310 11526 -12272
rect 11584 -12238 13184 -12222
rect 11584 -12272 11600 -12238
rect 13168 -12272 13184 -12238
rect 11584 -12310 13184 -12272
rect 8268 -12432 9868 -12394
rect 8268 -12466 8284 -12432
rect 9852 -12466 9868 -12432
rect 8268 -12482 9868 -12466
rect 9926 -12432 11526 -12394
rect 9926 -12466 9942 -12432
rect 11510 -12466 11526 -12432
rect 9926 -12482 11526 -12466
rect 11584 -12432 13184 -12394
rect 11584 -12466 11600 -12432
rect 13168 -12466 13184 -12432
rect 11584 -12482 13184 -12466
rect 19910 -12762 19998 -12746
rect 19910 -13130 19926 -12762
rect 19960 -13130 19998 -12762
rect 19910 -13146 19998 -13130
rect 20798 -12762 20908 -12746
rect 20798 -13130 20836 -12762
rect 20870 -13130 20908 -12762
rect 20798 -13146 20908 -13130
rect 21708 -12762 21796 -12746
rect 21708 -13130 21746 -12762
rect 21780 -13130 21796 -12762
rect 21708 -13146 21796 -13130
rect 19910 -13340 19998 -13324
rect 19910 -13708 19926 -13340
rect 19960 -13708 19998 -13340
rect 19910 -13724 19998 -13708
rect 20798 -13340 20908 -13324
rect 20798 -13708 20836 -13340
rect 20870 -13708 20908 -13340
rect 20798 -13724 20908 -13708
rect 21708 -13340 21796 -13324
rect 21708 -13708 21746 -13340
rect 21780 -13708 21796 -13340
rect 21708 -13724 21796 -13708
rect 19910 -13918 19998 -13902
rect 19910 -14286 19926 -13918
rect 19960 -14286 19998 -13918
rect 19910 -14302 19998 -14286
rect 20798 -13918 20908 -13902
rect 20798 -14286 20836 -13918
rect 20870 -14286 20908 -13918
rect 20798 -14302 20908 -14286
rect 21708 -13918 21796 -13902
rect 21708 -14286 21746 -13918
rect 21780 -14286 21796 -13918
rect 21708 -14302 21796 -14286
rect 19910 -14496 19998 -14480
rect 19910 -14864 19926 -14496
rect 19960 -14864 19998 -14496
rect 19910 -14880 19998 -14864
rect 20798 -14496 20908 -14480
rect 20798 -14864 20836 -14496
rect 20870 -14864 20908 -14496
rect 20798 -14880 20908 -14864
rect 21708 -14496 21796 -14480
rect 21708 -14864 21746 -14496
rect 21780 -14864 21796 -14496
rect 21708 -14880 21796 -14864
rect 19910 -15074 19998 -15058
rect 19910 -15442 19926 -15074
rect 19960 -15442 19998 -15074
rect 19910 -15458 19998 -15442
rect 20798 -15074 20908 -15058
rect 20798 -15442 20836 -15074
rect 20870 -15442 20908 -15074
rect 20798 -15458 20908 -15442
rect 21708 -15074 21796 -15058
rect 21708 -15442 21746 -15074
rect 21780 -15442 21796 -15074
rect 21708 -15458 21796 -15442
rect 20376 -16106 20464 -16090
rect 20376 -16174 20392 -16106
rect 20426 -16174 20464 -16106
rect 20376 -16190 20464 -16174
rect 21264 -16106 21352 -16090
rect 21264 -16174 21302 -16106
rect 21336 -16174 21352 -16106
rect 21264 -16190 21352 -16174
rect 20376 -16264 20464 -16248
rect 20376 -16332 20392 -16264
rect 20426 -16332 20464 -16264
rect 20376 -16348 20464 -16332
rect 21264 -16264 21352 -16248
rect 21264 -16332 21302 -16264
rect 21336 -16332 21352 -16264
rect 21264 -16348 21352 -16332
rect 20376 -16422 20464 -16406
rect 20376 -16490 20392 -16422
rect 20426 -16490 20464 -16422
rect 20376 -16506 20464 -16490
rect 21264 -16422 21352 -16406
rect 21264 -16490 21302 -16422
rect 21336 -16490 21352 -16422
rect 21264 -16506 21352 -16490
rect 20376 -16580 20464 -16564
rect 20376 -16648 20392 -16580
rect 20426 -16648 20464 -16580
rect 20376 -16664 20464 -16648
rect 21264 -16580 21352 -16564
rect 21264 -16648 21302 -16580
rect 21336 -16648 21352 -16580
rect 21264 -16664 21352 -16648
rect 20376 -16738 20464 -16722
rect 20376 -16806 20392 -16738
rect 20426 -16806 20464 -16738
rect 20376 -16822 20464 -16806
rect 21264 -16738 21352 -16722
rect 21264 -16806 21302 -16738
rect 21336 -16806 21352 -16738
rect 21264 -16822 21352 -16806
rect 20376 -16896 20464 -16880
rect 20376 -16964 20392 -16896
rect 20426 -16964 20464 -16896
rect 20376 -16980 20464 -16964
rect 21264 -16896 21352 -16880
rect 21264 -16964 21302 -16896
rect 21336 -16964 21352 -16896
rect 21264 -16980 21352 -16964
rect 20376 -17054 20464 -17038
rect 20376 -17122 20392 -17054
rect 20426 -17122 20464 -17054
rect 20376 -17138 20464 -17122
rect 21264 -17054 21352 -17038
rect 21264 -17122 21302 -17054
rect 21336 -17122 21352 -17054
rect 21264 -17138 21352 -17122
rect 20376 -17212 20464 -17196
rect 20376 -17280 20392 -17212
rect 20426 -17280 20464 -17212
rect 20376 -17296 20464 -17280
rect 21264 -17212 21352 -17196
rect 21264 -17280 21302 -17212
rect 21336 -17280 21352 -17212
rect 21264 -17296 21352 -17280
rect 20376 -17370 20464 -17354
rect 20376 -17438 20392 -17370
rect 20426 -17438 20464 -17370
rect 20376 -17454 20464 -17438
rect 21264 -17370 21352 -17354
rect 21264 -17438 21302 -17370
rect 21336 -17438 21352 -17370
rect 21264 -17454 21352 -17438
rect 20376 -17528 20464 -17512
rect 20376 -17596 20392 -17528
rect 20426 -17596 20464 -17528
rect 20376 -17612 20464 -17596
rect 21264 -17528 21352 -17512
rect 21264 -17596 21302 -17528
rect 21336 -17596 21352 -17528
rect 21264 -17612 21352 -17596
rect 20376 -17686 20464 -17670
rect 20376 -17754 20392 -17686
rect 20426 -17754 20464 -17686
rect 20376 -17770 20464 -17754
rect 21264 -17686 21352 -17670
rect 21264 -17754 21302 -17686
rect 21336 -17754 21352 -17686
rect 21264 -17770 21352 -17754
rect 20376 -17844 20464 -17828
rect 20376 -17912 20392 -17844
rect 20426 -17912 20464 -17844
rect 20376 -17928 20464 -17912
rect 21264 -17844 21352 -17828
rect 21264 -17912 21302 -17844
rect 21336 -17912 21352 -17844
rect 21264 -17928 21352 -17912
rect 22504 -12770 22601 -12754
rect 22504 -13138 22520 -12770
rect 22554 -13138 22601 -12770
rect 22504 -13154 22601 -13138
rect 23401 -12770 23529 -12754
rect 23401 -13138 23448 -12770
rect 23482 -13138 23529 -12770
rect 23401 -13154 23529 -13138
rect 24329 -12770 24426 -12754
rect 24329 -13138 24376 -12770
rect 24410 -13138 24426 -12770
rect 24329 -13154 24426 -13138
rect 22504 -13348 22601 -13332
rect 22504 -13716 22520 -13348
rect 22554 -13716 22601 -13348
rect 22504 -13732 22601 -13716
rect 23401 -13348 23529 -13332
rect 23401 -13716 23448 -13348
rect 23482 -13716 23529 -13348
rect 23401 -13732 23529 -13716
rect 24329 -13348 24426 -13332
rect 24329 -13716 24376 -13348
rect 24410 -13716 24426 -13348
rect 24329 -13732 24426 -13716
rect 22504 -13926 22601 -13910
rect 22504 -14294 22520 -13926
rect 22554 -14294 22601 -13926
rect 22504 -14310 22601 -14294
rect 23401 -13926 23529 -13910
rect 23401 -14294 23448 -13926
rect 23482 -14294 23529 -13926
rect 23401 -14310 23529 -14294
rect 24329 -13926 24426 -13910
rect 24329 -14294 24376 -13926
rect 24410 -14294 24426 -13926
rect 24329 -14310 24426 -14294
rect 22504 -14504 22601 -14488
rect 22504 -14872 22520 -14504
rect 22554 -14872 22601 -14504
rect 22504 -14888 22601 -14872
rect 23401 -14504 23529 -14488
rect 23401 -14872 23448 -14504
rect 23482 -14872 23529 -14504
rect 23401 -14888 23529 -14872
rect 24329 -14504 24426 -14488
rect 24329 -14872 24376 -14504
rect 24410 -14872 24426 -14504
rect 24329 -14888 24426 -14872
rect 22504 -15082 22601 -15066
rect 22504 -15450 22520 -15082
rect 22554 -15450 22601 -15082
rect 22504 -15466 22601 -15450
rect 23401 -15082 23529 -15066
rect 23401 -15450 23448 -15082
rect 23482 -15450 23529 -15082
rect 23401 -15466 23529 -15450
rect 24329 -15082 24426 -15066
rect 24329 -15450 24376 -15082
rect 24410 -15450 24426 -15082
rect 24329 -15466 24426 -15450
rect 22504 -15660 22601 -15644
rect 22504 -16028 22520 -15660
rect 22554 -16028 22601 -15660
rect 22504 -16044 22601 -16028
rect 23401 -15660 23529 -15644
rect 23401 -16028 23448 -15660
rect 23482 -16028 23529 -15660
rect 23401 -16044 23529 -16028
rect 24329 -15660 24426 -15644
rect 24329 -16028 24376 -15660
rect 24410 -16028 24426 -15660
rect 24329 -16044 24426 -16028
rect 22504 -16238 22601 -16222
rect 22504 -16606 22520 -16238
rect 22554 -16606 22601 -16238
rect 22504 -16622 22601 -16606
rect 23401 -16238 23529 -16222
rect 23401 -16606 23448 -16238
rect 23482 -16606 23529 -16238
rect 23401 -16622 23529 -16606
rect 24329 -16238 24426 -16222
rect 24329 -16606 24376 -16238
rect 24410 -16606 24426 -16238
rect 24329 -16622 24426 -16606
rect 22504 -16816 22601 -16800
rect 22504 -17184 22520 -16816
rect 22554 -17184 22601 -16816
rect 22504 -17200 22601 -17184
rect 23401 -16816 23529 -16800
rect 23401 -17184 23448 -16816
rect 23482 -17184 23529 -16816
rect 23401 -17200 23529 -17184
rect 24329 -16816 24426 -16800
rect 24329 -17184 24376 -16816
rect 24410 -17184 24426 -16816
rect 24329 -17200 24426 -17184
rect 22504 -17394 22601 -17378
rect 22504 -17762 22520 -17394
rect 22554 -17762 22601 -17394
rect 22504 -17778 22601 -17762
rect 23401 -17394 23529 -17378
rect 23401 -17762 23448 -17394
rect 23482 -17762 23529 -17394
rect 23401 -17778 23529 -17762
rect 24329 -17394 24426 -17378
rect 24329 -17762 24376 -17394
rect 24410 -17762 24426 -17394
rect 24329 -17778 24426 -17762
<< polycont >>
rect 3165 -1395 3199 -1361
rect 5131 -1395 5165 -1361
rect 3178 -1513 3212 -1479
rect 5118 -1513 5152 -1479
rect 14203 -1822 14237 -1788
rect 2828 -2084 2996 -2050
rect 2828 -2394 2996 -2360
rect 3428 -2076 3596 -2042
rect 3428 -2404 3596 -2370
rect 4740 -2076 4908 -2042
rect 4740 -2404 4908 -2370
rect 5340 -2084 5508 -2050
rect 14203 -1945 14237 -1911
rect 5340 -2394 5508 -2360
rect 7538 -2140 7606 -2106
rect 7696 -2140 7764 -2106
rect 7854 -2140 7922 -2106
rect 8012 -2140 8080 -2106
rect 8170 -2140 8238 -2106
rect 8328 -2140 8396 -2106
rect 8486 -2140 8554 -2106
rect 8644 -2140 8712 -2106
rect 8802 -2140 8870 -2106
rect 8960 -2140 9028 -2106
rect 7538 -3068 7606 -3034
rect 7696 -3068 7764 -3034
rect 7854 -3068 7922 -3034
rect 8012 -3068 8080 -3034
rect 8170 -3068 8238 -3034
rect 8328 -3068 8396 -3034
rect 8486 -3068 8554 -3034
rect 8644 -3068 8712 -3034
rect 8802 -3068 8870 -3034
rect 8960 -3068 9028 -3034
rect 9464 -2154 9532 -2120
rect 9622 -2154 9690 -2120
rect 9780 -2154 9848 -2120
rect 9938 -2154 10006 -2120
rect 10096 -2154 10164 -2120
rect 10254 -2154 10322 -2120
rect 10412 -2154 10480 -2120
rect 10570 -2154 10638 -2120
rect 10728 -2154 10796 -2120
rect 10886 -2154 10954 -2120
rect 9464 -3064 9532 -3030
rect 9622 -3064 9690 -3030
rect 9780 -3064 9848 -3030
rect 9938 -3064 10006 -3030
rect 10096 -3064 10164 -3030
rect 10254 -3064 10322 -3030
rect 10412 -3064 10480 -3030
rect 10570 -3064 10638 -3030
rect 10728 -3064 10796 -3030
rect 10886 -3064 10954 -3030
rect 11496 -2122 11564 -2088
rect 11496 -3050 11564 -3016
rect 14203 -2045 14237 -2011
rect 15012 -2042 15046 -2008
rect 12702 -3036 12736 -2268
rect 12912 -3036 12946 -2268
rect 14203 -2194 14237 -2160
rect 15012 -2110 15046 -2076
rect 15266 -1953 15300 -1919
rect 15164 -2003 15198 -1969
rect 15266 -2021 15300 -1987
rect 15544 -1999 15578 -1965
rect 15164 -2071 15198 -2037
rect 15646 -2014 15680 -1980
rect 16012 -1953 16046 -1919
rect 16114 -1947 16148 -1913
rect 15853 -2060 15887 -2026
rect 14203 -2301 14237 -2267
rect 16034 -2115 16068 -2081
rect 16369 -1953 16403 -1919
rect 16613 -1941 16647 -1907
rect 16283 -2089 16317 -2055
rect 16465 -2001 16499 -1967
rect 16709 -1989 16743 -1955
rect 16853 -1963 16887 -1929
rect 16748 -2115 16782 -2081
rect 16949 -1991 16983 -1957
rect 17149 -1999 17183 -1965
rect 17489 -1999 17523 -1965
rect 17752 -1999 17786 -1965
rect 17026 -2099 17060 -2065
rect 17854 -2014 17888 -1980
rect 18220 -1953 18254 -1919
rect 18322 -1947 18356 -1913
rect 18061 -2060 18095 -2026
rect 18242 -2115 18276 -2081
rect 18577 -1953 18611 -1919
rect 18821 -1941 18855 -1907
rect 18491 -2089 18525 -2055
rect 18673 -2001 18707 -1967
rect 18917 -1989 18951 -1955
rect 19061 -1963 19095 -1929
rect 18956 -2115 18990 -2081
rect 19157 -1991 19191 -1957
rect 19357 -1999 19391 -1965
rect 19697 -1999 19731 -1965
rect 19960 -1999 19994 -1965
rect 19234 -2099 19268 -2065
rect 20062 -2014 20096 -1980
rect 20428 -1953 20462 -1919
rect 20530 -1947 20564 -1913
rect 20269 -2060 20303 -2026
rect 20450 -2115 20484 -2081
rect 20785 -1953 20819 -1919
rect 21029 -1941 21063 -1907
rect 20699 -2089 20733 -2055
rect 20881 -2001 20915 -1967
rect 21125 -1989 21159 -1955
rect 21269 -1963 21303 -1929
rect 21164 -2115 21198 -2081
rect 21365 -1991 21399 -1957
rect 21565 -1999 21599 -1965
rect 21905 -1999 21939 -1965
rect 21442 -2099 21476 -2065
rect 14203 -2397 14237 -2363
rect 14203 -2588 14237 -2554
rect 15012 -2512 15046 -2478
rect 15012 -2580 15046 -2546
rect 14203 -2684 14237 -2650
rect 15164 -2551 15198 -2517
rect 15164 -2619 15198 -2585
rect 15266 -2601 15300 -2567
rect 15266 -2669 15300 -2635
rect 15544 -2623 15578 -2589
rect 15646 -2608 15680 -2574
rect 16034 -2507 16068 -2473
rect 15853 -2562 15887 -2528
rect 16283 -2533 16317 -2499
rect 14203 -2820 14237 -2786
rect 16012 -2669 16046 -2635
rect 16114 -2675 16148 -2641
rect 16369 -2669 16403 -2635
rect 16465 -2621 16499 -2587
rect 16748 -2507 16782 -2473
rect 16613 -2681 16647 -2647
rect 16709 -2633 16743 -2599
rect 17026 -2523 17060 -2489
rect 16853 -2659 16887 -2625
rect 16949 -2631 16983 -2597
rect 17149 -2623 17183 -2589
rect 17489 -2623 17523 -2589
rect 17752 -2623 17786 -2589
rect 17854 -2608 17888 -2574
rect 18242 -2507 18276 -2473
rect 18061 -2562 18095 -2528
rect 18491 -2533 18525 -2499
rect 18220 -2669 18254 -2635
rect 18322 -2675 18356 -2641
rect 18577 -2669 18611 -2635
rect 18673 -2621 18707 -2587
rect 18956 -2507 18990 -2473
rect 18821 -2681 18855 -2647
rect 18917 -2633 18951 -2599
rect 19234 -2523 19268 -2489
rect 19061 -2659 19095 -2625
rect 19157 -2631 19191 -2597
rect 19357 -2623 19391 -2589
rect 19697 -2623 19731 -2589
rect 19960 -2623 19994 -2589
rect 20062 -2608 20096 -2574
rect 20450 -2507 20484 -2473
rect 20269 -2562 20303 -2528
rect 20699 -2533 20733 -2499
rect 20428 -2669 20462 -2635
rect 20530 -2675 20564 -2641
rect 20785 -2669 20819 -2635
rect 20881 -2621 20915 -2587
rect 21164 -2507 21198 -2473
rect 21029 -2681 21063 -2647
rect 21125 -2633 21159 -2599
rect 21442 -2523 21476 -2489
rect 21269 -2659 21303 -2625
rect 21365 -2631 21399 -2597
rect 21565 -2623 21599 -2589
rect 21905 -2623 21939 -2589
rect 15172 -3128 15940 -3094
rect 15172 -3338 15940 -3304
rect 2744 -4088 2812 -4054
rect 2902 -4088 2970 -4054
rect 2744 -4798 2812 -4764
rect 2902 -4798 2970 -4764
rect 3450 -4088 3518 -4054
rect 3608 -4088 3676 -4054
rect 3450 -4798 3518 -4764
rect 3608 -4798 3676 -4764
rect 4660 -4088 4728 -4054
rect 4818 -4088 4886 -4054
rect 4660 -4798 4728 -4764
rect 4818 -4798 4886 -4764
rect 5366 -4088 5434 -4054
rect 5524 -4088 5592 -4054
rect 5366 -4798 5434 -4764
rect 5524 -4798 5592 -4764
rect 2826 -5382 3594 -5348
rect 2826 -5710 3594 -5676
rect 2826 -5986 3594 -5952
rect 2826 -6314 3594 -6280
rect 4742 -5382 5510 -5348
rect 4742 -5710 5510 -5676
rect 4742 -5986 5510 -5952
rect 4742 -6314 5510 -6280
rect 2513 -7215 2581 -7181
rect 2671 -7215 2739 -7181
rect 2829 -7215 2897 -7181
rect 2987 -7215 3055 -7181
rect 3145 -7215 3213 -7181
rect 2513 -8125 2581 -8091
rect 2671 -8125 2739 -8091
rect 2829 -8125 2897 -8091
rect 2987 -8125 3055 -8091
rect 3145 -8125 3213 -8091
rect 3888 -7208 3956 -7174
rect 4046 -7208 4114 -7174
rect 4204 -7208 4272 -7174
rect 4362 -7208 4430 -7174
rect 4520 -7208 4588 -7174
rect 3888 -8136 3956 -8102
rect 4046 -8136 4114 -8102
rect 4204 -8136 4272 -8102
rect 4362 -8136 4430 -8102
rect 4520 -8136 4588 -8102
rect 10674 -4920 11042 -4886
rect 11252 -4920 11620 -4886
rect 11830 -4920 12198 -4886
rect 12408 -4920 12776 -4886
rect 12986 -4920 13354 -4886
rect 13564 -4920 13932 -4886
rect 14142 -4920 14510 -4886
rect 14720 -4920 15088 -4886
rect 10674 -5430 11042 -5396
rect 11252 -5430 11620 -5396
rect 11830 -5430 12198 -5396
rect 12408 -5430 12776 -5396
rect 12986 -5430 13354 -5396
rect 13564 -5430 13932 -5396
rect 14142 -5430 14510 -5396
rect 14720 -5430 15088 -5396
rect 16276 -4700 16644 -4666
rect 16734 -4700 17102 -4666
rect 17192 -4700 17560 -4666
rect 17650 -4700 18018 -4666
rect 16276 -5610 16644 -5576
rect 16734 -5610 17102 -5576
rect 17192 -5610 17560 -5576
rect 17650 -5610 18018 -5576
rect 18964 -5496 20532 -5462
rect 18964 -5706 20532 -5672
rect 21428 -5368 21596 -5334
rect 21686 -5368 21854 -5334
rect 21428 -5578 21596 -5544
rect 21686 -5578 21854 -5544
rect 10698 -5942 11066 -5908
rect 11270 -5942 11638 -5908
rect 11842 -5942 12210 -5908
rect 12414 -5942 12782 -5908
rect 12986 -5942 13354 -5908
rect 13558 -5942 13926 -5908
rect 14130 -5942 14498 -5908
rect 14702 -5942 15070 -5908
rect 21428 -5788 21596 -5754
rect 21686 -5788 21854 -5754
rect 23362 -5632 23396 -5464
rect 23622 -5632 23656 -5464
rect 10698 -6470 11066 -6436
rect 11270 -6470 11638 -6436
rect 11842 -6470 12210 -6436
rect 12414 -6470 12782 -6436
rect 12986 -6470 13354 -6436
rect 13558 -6470 13926 -6436
rect 14130 -6470 14498 -6436
rect 14702 -6470 15070 -6436
rect 10698 -6998 11066 -6964
rect 11270 -6998 11638 -6964
rect 11842 -6998 12210 -6964
rect 12414 -6998 12782 -6964
rect 12986 -6998 13354 -6964
rect 13558 -6998 13926 -6964
rect 14130 -6998 14498 -6964
rect 14702 -6998 15070 -6964
rect 16276 -6050 16644 -6016
rect 16734 -6050 17102 -6016
rect 17192 -6050 17560 -6016
rect 17650 -6050 18018 -6016
rect 16276 -6978 16644 -6944
rect 16734 -6978 17102 -6944
rect 17192 -6978 17560 -6944
rect 17650 -6978 18018 -6944
rect 18944 -6500 20512 -6466
rect 18944 -6728 20512 -6694
rect 21428 -6364 21596 -6330
rect 21686 -6364 21854 -6330
rect 21428 -6592 21596 -6558
rect 21686 -6592 21854 -6558
rect 21428 -6820 21596 -6786
rect 21686 -6820 21854 -6786
rect 23050 -6634 23084 -6466
rect 23978 -6634 24012 -6466
rect 9136 -9330 9170 -7762
rect 9346 -9330 9380 -7762
rect 9716 -9064 9750 -7496
rect 9944 -9064 9978 -7496
rect 7342 -12212 7510 -12178
rect 7342 -12522 7510 -12488
rect 8284 -12272 9852 -12238
rect 9942 -12272 11510 -12238
rect 11600 -12272 13168 -12238
rect 8284 -12466 9852 -12432
rect 9942 -12466 11510 -12432
rect 11600 -12466 13168 -12432
rect 19926 -13130 19960 -12762
rect 20836 -13130 20870 -12762
rect 21746 -13130 21780 -12762
rect 19926 -13708 19960 -13340
rect 20836 -13708 20870 -13340
rect 21746 -13708 21780 -13340
rect 19926 -14286 19960 -13918
rect 20836 -14286 20870 -13918
rect 21746 -14286 21780 -13918
rect 19926 -14864 19960 -14496
rect 20836 -14864 20870 -14496
rect 21746 -14864 21780 -14496
rect 19926 -15442 19960 -15074
rect 20836 -15442 20870 -15074
rect 21746 -15442 21780 -15074
rect 20392 -16174 20426 -16106
rect 21302 -16174 21336 -16106
rect 20392 -16332 20426 -16264
rect 21302 -16332 21336 -16264
rect 20392 -16490 20426 -16422
rect 21302 -16490 21336 -16422
rect 20392 -16648 20426 -16580
rect 21302 -16648 21336 -16580
rect 20392 -16806 20426 -16738
rect 21302 -16806 21336 -16738
rect 20392 -16964 20426 -16896
rect 21302 -16964 21336 -16896
rect 20392 -17122 20426 -17054
rect 21302 -17122 21336 -17054
rect 20392 -17280 20426 -17212
rect 21302 -17280 21336 -17212
rect 20392 -17438 20426 -17370
rect 21302 -17438 21336 -17370
rect 20392 -17596 20426 -17528
rect 21302 -17596 21336 -17528
rect 20392 -17754 20426 -17686
rect 21302 -17754 21336 -17686
rect 20392 -17912 20426 -17844
rect 21302 -17912 21336 -17844
rect 22520 -13138 22554 -12770
rect 23448 -13138 23482 -12770
rect 24376 -13138 24410 -12770
rect 22520 -13716 22554 -13348
rect 23448 -13716 23482 -13348
rect 24376 -13716 24410 -13348
rect 22520 -14294 22554 -13926
rect 23448 -14294 23482 -13926
rect 24376 -14294 24410 -13926
rect 22520 -14872 22554 -14504
rect 23448 -14872 23482 -14504
rect 24376 -14872 24410 -14504
rect 22520 -15450 22554 -15082
rect 23448 -15450 23482 -15082
rect 24376 -15450 24410 -15082
rect 22520 -16028 22554 -15660
rect 23448 -16028 23482 -15660
rect 24376 -16028 24410 -15660
rect 22520 -16606 22554 -16238
rect 23448 -16606 23482 -16238
rect 24376 -16606 24410 -16238
rect 22520 -17184 22554 -16816
rect 23448 -17184 23482 -16816
rect 24376 -17184 24410 -16816
rect 22520 -17762 22554 -17394
rect 23448 -17762 23482 -17394
rect 24376 -17762 24410 -17394
<< xpolycontact >>
rect 10620 -7508 11052 -7438
rect 24220 -7508 24652 -7438
rect 10620 -7674 11052 -7604
rect 24220 -7674 24652 -7604
rect 10620 -7840 11052 -7770
rect 24220 -7840 24652 -7770
rect 10620 -8006 11052 -7936
rect 24220 -8006 24652 -7936
rect 10620 -8172 11052 -8102
rect 24220 -8172 24652 -8102
rect 10620 -8338 11052 -8268
rect 24220 -8338 24652 -8268
rect 10620 -8504 11052 -8434
rect 24220 -8504 24652 -8434
rect 10620 -8670 11052 -8600
rect 24220 -8670 24652 -8600
rect 10620 -8836 11052 -8766
rect 24220 -8836 24652 -8766
rect 10620 -9002 11052 -8932
rect 24220 -9002 24652 -8932
rect 10620 -9168 11052 -9098
rect 24220 -9168 24652 -9098
rect 10620 -9334 11052 -9264
rect 24220 -9334 24652 -9264
rect 10620 -9500 11052 -9430
rect 24220 -9500 24652 -9430
rect 10620 -9666 11052 -9596
rect 24220 -9666 24652 -9596
rect 10620 -9832 11052 -9762
rect 24220 -9832 24652 -9762
rect 3134 -12992 3566 -12922
rect 18534 -12992 18966 -12922
rect 3134 -13158 3566 -13088
rect 18534 -13158 18966 -13088
rect 3134 -13324 3566 -13254
rect 18534 -13324 18966 -13254
rect 3134 -13490 3566 -13420
rect 18534 -13490 18966 -13420
rect 2132 -13930 2564 -13860
rect 18932 -13930 19364 -13860
rect 2132 -14096 2564 -14026
rect 18932 -14096 19364 -14026
rect 2132 -14262 2564 -14192
rect 18932 -14262 19364 -14192
rect 2132 -14428 2564 -14358
rect 18932 -14428 19364 -14358
rect 2132 -14594 2564 -14524
rect 18932 -14594 19364 -14524
rect 2132 -14760 2564 -14690
rect 18932 -14760 19364 -14690
rect 2132 -14926 2564 -14856
rect 18932 -14926 19364 -14856
rect 2132 -15092 2564 -15022
rect 18932 -15092 19364 -15022
rect 2132 -15258 2564 -15188
rect 18932 -15258 19364 -15188
rect 2132 -15424 2564 -15354
rect 18932 -15424 19364 -15354
rect 2132 -15590 2564 -15520
rect 18932 -15590 19364 -15520
rect 2132 -15756 2564 -15686
rect 18932 -15756 19364 -15686
rect 2132 -15922 2564 -15852
rect 18932 -15922 19364 -15852
rect 2132 -16088 2564 -16018
rect 18932 -16088 19364 -16018
rect 2132 -16254 2564 -16184
rect 18932 -16254 19364 -16184
rect 2132 -16420 2564 -16350
rect 18932 -16420 19364 -16350
rect 2132 -16586 2564 -16516
rect 18932 -16586 19364 -16516
rect 2132 -16752 2564 -16682
rect 18932 -16752 19364 -16682
rect 2132 -16918 2564 -16848
rect 18932 -16918 19364 -16848
rect 2132 -17084 2564 -17014
rect 18932 -17084 19364 -17014
rect 2132 -17250 2564 -17180
rect 18932 -17250 19364 -17180
rect 2132 -17416 2564 -17346
rect 18932 -17416 19364 -17346
rect 2132 -17582 2564 -17512
rect 18932 -17582 19364 -17512
rect 2132 -17748 2564 -17678
rect 18932 -17748 19364 -17678
rect 2132 -17914 2564 -17844
rect 18932 -17914 19364 -17844
rect 2132 -18080 2564 -18010
rect 18932 -18080 19364 -18010
rect 2130 -18520 2562 -18450
rect 24530 -18520 24962 -18450
rect 2130 -18686 2562 -18616
rect 24530 -18686 24962 -18616
rect 2130 -18852 2562 -18782
rect 24530 -18852 24962 -18782
rect 2130 -19018 2562 -18948
rect 24530 -19018 24962 -18948
rect 2130 -19184 2562 -19114
rect 24530 -19184 24962 -19114
rect 2130 -19350 2562 -19280
rect 24530 -19350 24962 -19280
rect 2130 -19516 2562 -19446
rect 24530 -19516 24962 -19446
rect 2130 -19682 2562 -19612
rect 24530 -19682 24962 -19612
rect 2130 -19848 2562 -19778
rect 24530 -19848 24962 -19778
rect 2130 -20014 2562 -19944
rect 24530 -20014 24962 -19944
rect 2130 -20180 2562 -20110
rect 24530 -20180 24962 -20110
rect 2130 -20346 2562 -20276
rect 24530 -20346 24962 -20276
rect 2130 -20512 2562 -20442
rect 24530 -20512 24962 -20442
rect 2130 -20678 2562 -20608
rect 24530 -20678 24962 -20608
rect 2130 -20844 2562 -20774
rect 24530 -20844 24962 -20774
rect 2130 -21010 2562 -20940
rect 24530 -21010 24962 -20940
rect 2130 -21176 2562 -21106
rect 24530 -21176 24962 -21106
rect 2130 -21342 2562 -21272
rect 24530 -21342 24962 -21272
rect 2130 -21508 2562 -21438
rect 24530 -21508 24962 -21438
rect 2130 -21674 2562 -21604
rect 24530 -21674 24962 -21604
rect 2130 -21840 2562 -21770
rect 24530 -21840 24962 -21770
rect 2130 -22006 2562 -21936
rect 24530 -22006 24962 -21936
rect 2130 -22172 2562 -22102
rect 24530 -22172 24962 -22102
rect 2130 -22338 2562 -22268
rect 24530 -22338 24962 -22268
rect 2130 -22504 2562 -22434
rect 24530 -22504 24962 -22434
<< xpolyres >>
rect 11052 -7508 24220 -7438
rect 11052 -7674 24220 -7604
rect 11052 -7840 24220 -7770
rect 11052 -8006 24220 -7936
rect 11052 -8172 24220 -8102
rect 11052 -8338 24220 -8268
rect 11052 -8504 24220 -8434
rect 11052 -8670 24220 -8600
rect 11052 -8836 24220 -8766
rect 11052 -9002 24220 -8932
rect 11052 -9168 24220 -9098
rect 11052 -9334 24220 -9264
rect 11052 -9500 24220 -9430
rect 11052 -9666 24220 -9596
rect 11052 -9832 24220 -9762
rect 3566 -12992 18534 -12922
rect 3566 -13158 18534 -13088
rect 3566 -13324 18534 -13254
rect 3566 -13490 18534 -13420
rect 2564 -13930 18932 -13860
rect 2564 -14096 18932 -14026
rect 2564 -14262 18932 -14192
rect 2564 -14428 18932 -14358
rect 2564 -14594 18932 -14524
rect 2564 -14760 18932 -14690
rect 2564 -14926 18932 -14856
rect 2564 -15092 18932 -15022
rect 2564 -15258 18932 -15188
rect 2564 -15424 18932 -15354
rect 2564 -15590 18932 -15520
rect 2564 -15756 18932 -15686
rect 2564 -15922 18932 -15852
rect 2564 -16088 18932 -16018
rect 2564 -16254 18932 -16184
rect 2564 -16420 18932 -16350
rect 2564 -16586 18932 -16516
rect 2564 -16752 18932 -16682
rect 2564 -16918 18932 -16848
rect 2564 -17084 18932 -17014
rect 2564 -17250 18932 -17180
rect 2564 -17416 18932 -17346
rect 2564 -17582 18932 -17512
rect 2564 -17748 18932 -17678
rect 2564 -17914 18932 -17844
rect 2564 -18080 18932 -18010
rect 2562 -18520 24530 -18450
rect 2562 -18686 24530 -18616
rect 2562 -18852 24530 -18782
rect 2562 -19018 24530 -18948
rect 2562 -19184 24530 -19114
rect 2562 -19350 24530 -19280
rect 2562 -19516 24530 -19446
rect 2562 -19682 24530 -19612
rect 2562 -19848 24530 -19778
rect 2562 -20014 24530 -19944
rect 2562 -20180 24530 -20110
rect 2562 -20346 24530 -20276
rect 2562 -20512 24530 -20442
rect 2562 -20678 24530 -20608
rect 2562 -20844 24530 -20774
rect 2562 -21010 24530 -20940
rect 2562 -21176 24530 -21106
rect 2562 -21342 24530 -21272
rect 2562 -21508 24530 -21438
rect 2562 -21674 24530 -21604
rect 2562 -21840 24530 -21770
rect 2562 -22006 24530 -21936
rect 2562 -22172 24530 -22102
rect 2562 -22338 24530 -22268
rect 2562 -22504 24530 -22434
<< pdiode >>
rect 21316 -22942 21406 -22930
rect 21316 -23008 21328 -22942
rect 21394 -23008 21406 -22942
rect 21316 -23020 21406 -23008
rect 22742 -22944 22832 -22932
rect 22742 -23010 22754 -22944
rect 22820 -23010 22832 -22944
rect 22742 -23022 22832 -23010
<< ndiode >>
rect 2888 -964 2978 -952
rect 2888 -1030 2900 -964
rect 2966 -1030 2978 -964
rect 2888 -1042 2978 -1030
rect 5358 -964 5448 -952
rect 5358 -1030 5370 -964
rect 5436 -1030 5448 -964
rect 5358 -1042 5448 -1030
rect 20460 -22952 20550 -22940
rect 20460 -23018 20472 -22952
rect 20538 -23018 20550 -22952
rect 20460 -23030 20550 -23018
rect 23568 -22954 23658 -22942
rect 23568 -23020 23580 -22954
rect 23646 -23020 23658 -22954
rect 23568 -23032 23658 -23020
<< pdiodec >>
rect 21328 -23008 21394 -22942
rect 22754 -23010 22820 -22944
<< ndiodec >>
rect 2900 -1030 2966 -964
rect 5370 -1030 5436 -964
rect 20472 -23018 20538 -22952
rect 23580 -23020 23646 -22954
<< locali >>
rect 2748 -864 2882 -850
rect 2806 -884 2882 -864
rect 2984 -884 3080 -850
rect 2806 -946 2820 -884
rect 3046 -946 3080 -884
rect 5256 -884 5352 -850
rect 5454 -884 5586 -850
rect 5256 -946 5290 -884
rect 2884 -1030 2900 -964
rect 2966 -1030 2982 -964
rect 2806 -1110 2820 -1048
rect 3046 -1110 3080 -1048
rect 2806 -1128 2882 -1110
rect 2984 -1128 3080 -1110
rect 3018 -1144 3080 -1128
rect 3146 -956 3246 -946
rect 3018 -1182 3046 -1144
rect 3146 -1180 3156 -956
rect 3236 -1180 3246 -956
rect 3146 -1194 3246 -1180
rect 5086 -958 5186 -948
rect 5086 -1180 5096 -958
rect 5176 -1180 5186 -958
rect 5516 -946 5530 -884
rect 5354 -1030 5370 -964
rect 5436 -1030 5452 -964
rect 5256 -1110 5290 -1048
rect 5516 -1110 5530 -1048
rect 5256 -1126 5352 -1110
rect 5454 -1126 5530 -1110
rect 5256 -1144 5316 -1126
rect 5290 -1180 5316 -1144
rect 5086 -1192 5186 -1180
rect 2933 -1249 2967 -1232
rect 2933 -1261 3112 -1249
rect 2967 -1295 3061 -1261
rect 3095 -1295 3112 -1261
rect 2933 -1307 3112 -1295
rect 2933 -1353 2967 -1307
rect 3146 -1345 3210 -1194
rect 3477 -1249 3511 -1232
rect 3244 -1261 3511 -1249
rect 3244 -1295 3279 -1261
rect 3313 -1295 3372 -1261
rect 3406 -1295 3477 -1261
rect 3244 -1307 3511 -1295
rect 3146 -1358 3221 -1345
rect 3477 -1353 3511 -1307
rect 2933 -1429 2967 -1387
rect 3001 -1393 3022 -1359
rect 3056 -1393 3111 -1359
rect 2933 -1445 3043 -1429
rect 2967 -1479 3009 -1445
rect 2933 -1495 3043 -1479
rect 3077 -1458 3111 -1393
rect 3147 -1361 3221 -1358
rect 3147 -1395 3165 -1361
rect 3199 -1395 3221 -1361
rect 3147 -1413 3221 -1395
rect 3257 -1359 3443 -1357
rect 3257 -1393 3325 -1359
rect 3359 -1393 3393 -1359
rect 3427 -1393 3443 -1359
rect 3257 -1458 3291 -1393
rect 3477 -1429 3511 -1387
rect 3077 -1479 3291 -1458
rect 3077 -1492 3178 -1479
rect 2933 -1537 2967 -1495
rect 3162 -1513 3178 -1492
rect 3212 -1492 3291 -1479
rect 3325 -1445 3511 -1429
rect 3359 -1479 3393 -1445
rect 3427 -1479 3477 -1445
rect 3212 -1513 3228 -1492
rect 3325 -1495 3511 -1479
rect 3262 -1531 3443 -1529
rect 2933 -1600 2967 -1571
rect 3001 -1565 3039 -1531
rect 3073 -1547 3102 -1531
rect 3262 -1547 3312 -1531
rect 3073 -1565 3312 -1547
rect 3346 -1565 3393 -1531
rect 3427 -1565 3443 -1531
rect 3001 -1583 3443 -1565
rect 3477 -1537 3511 -1495
rect 3038 -1694 3426 -1583
rect 3477 -1600 3511 -1571
rect 4819 -1249 4853 -1232
rect 4819 -1261 5086 -1249
rect 4853 -1295 4924 -1261
rect 4958 -1295 5017 -1261
rect 5051 -1295 5086 -1261
rect 4819 -1307 5086 -1295
rect 4819 -1353 4853 -1307
rect 5120 -1345 5184 -1192
rect 5363 -1249 5397 -1232
rect 5218 -1261 5397 -1249
rect 5218 -1295 5235 -1261
rect 5269 -1295 5363 -1261
rect 5218 -1307 5397 -1295
rect 5109 -1350 5184 -1345
rect 4819 -1429 4853 -1387
rect 4887 -1359 5073 -1357
rect 4887 -1393 4903 -1359
rect 4937 -1393 4971 -1359
rect 5005 -1393 5073 -1359
rect 4819 -1445 5005 -1429
rect 4853 -1479 4903 -1445
rect 4937 -1479 4971 -1445
rect 4819 -1495 5005 -1479
rect 5039 -1458 5073 -1393
rect 5109 -1361 5183 -1350
rect 5363 -1353 5397 -1307
rect 5109 -1395 5131 -1361
rect 5165 -1395 5183 -1361
rect 5109 -1413 5183 -1395
rect 5219 -1393 5274 -1359
rect 5308 -1393 5329 -1359
rect 5219 -1458 5253 -1393
rect 5363 -1429 5397 -1387
rect 5039 -1479 5253 -1458
rect 5039 -1492 5118 -1479
rect 4819 -1537 4853 -1495
rect 5102 -1513 5118 -1492
rect 5152 -1492 5253 -1479
rect 5287 -1445 5397 -1429
rect 5321 -1479 5363 -1445
rect 5152 -1513 5168 -1492
rect 5287 -1495 5397 -1479
rect 4819 -1600 4853 -1571
rect 4887 -1531 5068 -1529
rect 4887 -1565 4903 -1531
rect 4937 -1565 4984 -1531
rect 5018 -1547 5068 -1531
rect 5228 -1547 5257 -1531
rect 5018 -1565 5257 -1547
rect 5291 -1565 5329 -1531
rect 4887 -1583 5329 -1565
rect 5363 -1537 5397 -1495
rect 3038 -1768 3050 -1694
rect 3412 -1768 3426 -1694
rect 3038 -1780 3426 -1768
rect 4904 -1686 5292 -1583
rect 5363 -1600 5397 -1571
rect 13662 -1580 14244 -1566
rect 4904 -1760 4916 -1686
rect 5278 -1760 5292 -1686
rect 4904 -1772 5292 -1760
rect 13662 -1752 13676 -1580
rect 13848 -1616 14244 -1580
rect 13848 -1752 13862 -1616
rect 13662 -1766 13862 -1752
rect 13971 -1675 14005 -1658
rect 13971 -1687 14150 -1675
rect 14005 -1721 14099 -1687
rect 14133 -1721 14150 -1687
rect 13971 -1733 14150 -1721
rect 13971 -1779 14005 -1733
rect 14204 -1768 14244 -1616
rect 14515 -1675 14549 -1658
rect 14282 -1687 14549 -1675
rect 14282 -1721 14317 -1687
rect 14351 -1721 14410 -1687
rect 14444 -1721 14515 -1687
rect 14282 -1733 14549 -1721
rect 13971 -1853 14005 -1813
rect 14039 -1819 14083 -1785
rect 14117 -1819 14169 -1785
rect 13971 -1869 14101 -1853
rect 13971 -1871 14059 -1869
rect 14005 -1903 14059 -1871
rect 14093 -1903 14101 -1869
rect 14005 -1905 14101 -1903
rect 13971 -1919 14101 -1905
rect 3076 -1982 3172 -1948
rect 3138 -2044 3172 -1982
rect 2812 -2084 2828 -2050
rect 2996 -2084 3012 -2050
rect 2766 -2134 2800 -2118
rect 2766 -2326 2800 -2310
rect 3024 -2134 3058 -2118
rect 3024 -2326 3058 -2310
rect 2812 -2394 2828 -2360
rect 2996 -2394 3012 -2360
rect 3138 -2462 3172 -2400
rect 3076 -2496 3172 -2462
rect 3252 -1974 3348 -1940
rect 3252 -2036 3286 -1974
rect 3412 -2076 3428 -2042
rect 3596 -2076 3612 -2042
rect 3366 -2135 3400 -2119
rect 3366 -2327 3400 -2311
rect 3624 -2135 3658 -2119
rect 3624 -2327 3658 -2311
rect 3412 -2404 3428 -2370
rect 3596 -2404 3612 -2370
rect 3252 -2472 3286 -2410
rect 3252 -2506 3348 -2472
rect 4988 -1974 5084 -1940
rect 5050 -2036 5084 -1974
rect 4724 -2076 4740 -2042
rect 4908 -2076 4924 -2042
rect 4678 -2135 4712 -2119
rect 4678 -2327 4712 -2311
rect 4936 -2135 4970 -2119
rect 4936 -2327 4970 -2311
rect 4724 -2404 4740 -2370
rect 4908 -2404 4924 -2370
rect 5050 -2472 5084 -2410
rect 4988 -2506 5084 -2472
rect 5164 -1982 5260 -1948
rect 5164 -2044 5198 -1982
rect 11300 -1984 11396 -1950
rect 11664 -1984 11760 -1950
rect 5324 -2084 5340 -2050
rect 5508 -2084 5524 -2050
rect 5278 -2134 5312 -2118
rect 5278 -2326 5312 -2310
rect 5536 -2134 5570 -2118
rect 5536 -2326 5570 -2310
rect 5324 -2394 5340 -2360
rect 5508 -2394 5524 -2360
rect 5164 -2462 5198 -2400
rect 5164 -2496 5260 -2462
rect 7362 -2038 7458 -2004
rect 9108 -2038 9204 -2004
rect 7362 -2100 7396 -2038
rect 7506 -2082 9044 -2072
rect 7506 -2128 7514 -2082
rect 9032 -2128 9044 -2082
rect 7506 -2140 7538 -2128
rect 7606 -2140 7696 -2128
rect 7764 -2140 7854 -2128
rect 7922 -2140 8012 -2128
rect 8080 -2140 8170 -2128
rect 8238 -2140 8328 -2128
rect 8396 -2140 8486 -2128
rect 8554 -2140 8644 -2128
rect 8712 -2140 8802 -2128
rect 8870 -2140 8960 -2128
rect 9028 -2140 9044 -2128
rect 9170 -2100 9204 -2038
rect 7476 -2184 7510 -2183
rect 7396 -2188 7510 -2184
rect 7634 -2188 7668 -2183
rect 7792 -2188 7826 -2183
rect 7950 -2188 7984 -2183
rect 8108 -2188 8142 -2183
rect 8266 -2186 8300 -2183
rect 7396 -2198 7552 -2188
rect 7396 -2976 7444 -2198
rect 7540 -2976 7552 -2198
rect 7396 -2988 7552 -2976
rect 7592 -2198 7712 -2188
rect 7592 -2976 7604 -2198
rect 7700 -2976 7712 -2198
rect 7592 -2988 7712 -2976
rect 7750 -2198 7870 -2188
rect 7750 -2976 7762 -2198
rect 7858 -2976 7870 -2198
rect 7750 -2988 7870 -2976
rect 7908 -2198 8028 -2188
rect 7908 -2976 7920 -2198
rect 8016 -2976 8028 -2198
rect 7908 -2988 8028 -2976
rect 8066 -2198 8186 -2188
rect 8066 -2976 8078 -2198
rect 8174 -2976 8186 -2198
rect 8066 -2988 8186 -2976
rect 8222 -2198 8342 -2186
rect 8424 -2188 8458 -2183
rect 8582 -2186 8616 -2183
rect 8222 -2976 8234 -2198
rect 8330 -2976 8342 -2198
rect 8222 -2986 8342 -2976
rect 8380 -2198 8500 -2188
rect 8380 -2976 8392 -2198
rect 8488 -2976 8500 -2198
rect 7476 -2991 7510 -2988
rect 7634 -2991 7668 -2988
rect 7792 -2991 7826 -2988
rect 7950 -2991 7984 -2988
rect 8108 -2991 8142 -2988
rect 8266 -2991 8300 -2986
rect 8380 -2988 8500 -2976
rect 8540 -2198 8660 -2186
rect 8740 -2188 8774 -2183
rect 8898 -2188 8932 -2183
rect 9056 -2186 9090 -2183
rect 9056 -2188 9170 -2186
rect 8540 -2976 8552 -2198
rect 8648 -2976 8660 -2198
rect 8540 -2986 8660 -2976
rect 8696 -2198 8816 -2188
rect 8696 -2976 8708 -2198
rect 8804 -2976 8816 -2198
rect 8424 -2991 8458 -2988
rect 8582 -2991 8616 -2986
rect 8696 -2988 8816 -2976
rect 8854 -2198 8974 -2188
rect 8854 -2976 8866 -2198
rect 8962 -2976 8974 -2198
rect 8854 -2988 8974 -2976
rect 9012 -2198 9170 -2188
rect 9012 -2976 9024 -2198
rect 9120 -2976 9170 -2198
rect 9012 -2988 9170 -2976
rect 8740 -2991 8774 -2988
rect 8898 -2991 8932 -2988
rect 9056 -2990 9170 -2988
rect 9056 -2991 9090 -2990
rect 7362 -3136 7396 -3074
rect 7502 -3046 7538 -3034
rect 7606 -3046 7696 -3034
rect 7764 -3046 7854 -3034
rect 7922 -3046 8012 -3034
rect 8080 -3046 8170 -3034
rect 8238 -3046 8328 -3034
rect 8396 -3046 8486 -3034
rect 8554 -3046 8644 -3034
rect 8712 -3046 8802 -3034
rect 8870 -3046 8960 -3034
rect 9028 -3046 9044 -3034
rect 7502 -3092 7512 -3046
rect 9034 -3092 9044 -3046
rect 7502 -3102 9044 -3092
rect 9170 -3136 9204 -3074
rect 7362 -3170 7458 -3136
rect 9108 -3170 9204 -3136
rect 9288 -2052 9384 -2018
rect 11034 -2052 11130 -2018
rect 9288 -2114 9322 -2052
rect 9428 -2092 10970 -2086
rect 9428 -2140 9438 -2092
rect 10952 -2120 10970 -2092
rect 9428 -2154 9464 -2140
rect 9532 -2154 9622 -2140
rect 9690 -2154 9780 -2140
rect 9848 -2154 9938 -2140
rect 10006 -2154 10096 -2140
rect 10164 -2154 10254 -2140
rect 10322 -2154 10412 -2140
rect 10480 -2154 10570 -2140
rect 10638 -2154 10728 -2140
rect 10796 -2154 10886 -2140
rect 10954 -2154 10970 -2120
rect 11096 -2114 11130 -2052
rect 9402 -2190 9436 -2188
rect 9322 -2192 9436 -2190
rect 9560 -2192 9594 -2188
rect 9718 -2192 9752 -2188
rect 9876 -2192 9910 -2188
rect 10034 -2192 10068 -2188
rect 10192 -2192 10226 -2188
rect 10350 -2192 10384 -2188
rect 10508 -2192 10542 -2188
rect 10666 -2192 10700 -2188
rect 10824 -2192 10858 -2188
rect 10982 -2190 11016 -2188
rect 10982 -2192 11096 -2190
rect 9322 -2202 9478 -2192
rect 9322 -2980 9370 -2202
rect 9466 -2980 9478 -2202
rect 9322 -2992 9478 -2980
rect 9516 -2202 9636 -2192
rect 9516 -2980 9528 -2202
rect 9624 -2980 9636 -2202
rect 9516 -2992 9636 -2980
rect 9676 -2202 9796 -2192
rect 9676 -2980 9688 -2202
rect 9784 -2980 9796 -2202
rect 9676 -2992 9796 -2980
rect 9834 -2202 9954 -2192
rect 9834 -2980 9846 -2202
rect 9942 -2980 9954 -2202
rect 9834 -2992 9954 -2980
rect 9990 -2202 10110 -2192
rect 9990 -2980 10002 -2202
rect 10098 -2980 10110 -2202
rect 9990 -2992 10110 -2980
rect 10150 -2202 10270 -2192
rect 10150 -2980 10162 -2202
rect 10258 -2980 10270 -2202
rect 10150 -2992 10270 -2980
rect 10306 -2202 10426 -2192
rect 10306 -2980 10318 -2202
rect 10414 -2980 10426 -2202
rect 10306 -2992 10426 -2980
rect 10464 -2202 10584 -2192
rect 10464 -2980 10476 -2202
rect 10572 -2980 10584 -2202
rect 10464 -2992 10584 -2980
rect 10624 -2202 10744 -2192
rect 10624 -2980 10636 -2202
rect 10732 -2980 10744 -2202
rect 10624 -2992 10744 -2980
rect 10780 -2202 10900 -2192
rect 10780 -2980 10792 -2202
rect 10888 -2980 10900 -2202
rect 10780 -2992 10900 -2980
rect 10938 -2202 11096 -2192
rect 10938 -2980 10950 -2202
rect 11046 -2980 11096 -2202
rect 10938 -2992 11096 -2980
rect 9322 -2994 9436 -2992
rect 9402 -2996 9436 -2994
rect 9560 -2996 9594 -2992
rect 9718 -2996 9752 -2992
rect 9876 -2996 9910 -2992
rect 10034 -2996 10068 -2992
rect 10192 -2996 10226 -2992
rect 10350 -2996 10384 -2992
rect 10508 -2996 10542 -2992
rect 10666 -2996 10700 -2992
rect 10824 -2996 10858 -2992
rect 10982 -2994 11096 -2992
rect 10982 -2996 11016 -2994
rect 9288 -3132 9322 -3070
rect 9426 -3044 9464 -3030
rect 9532 -3044 9622 -3030
rect 9690 -3044 9780 -3030
rect 9848 -3044 9938 -3030
rect 10006 -3044 10096 -3030
rect 10164 -3044 10254 -3030
rect 10322 -3044 10412 -3030
rect 10480 -3044 10570 -3030
rect 10638 -3044 10728 -3030
rect 10796 -3044 10886 -3030
rect 9426 -3092 9436 -3044
rect 10954 -3064 10970 -3030
rect 10952 -3092 10970 -3064
rect 9426 -3098 10970 -3092
rect 11096 -3132 11130 -3070
rect 9288 -3166 9384 -3132
rect 11034 -3166 11130 -3132
rect 11300 -2046 11334 -1984
rect 11726 -2046 11760 -1984
rect 11480 -2122 11496 -2088
rect 11564 -2122 11580 -2088
rect 11334 -2180 11474 -2164
rect 11468 -2958 11474 -2180
rect 11334 -2974 11474 -2958
rect 11592 -2170 11626 -2165
rect 11592 -2181 11678 -2170
rect 11626 -2182 11678 -2181
rect 11666 -2956 11678 -2182
rect 11626 -2957 11678 -2956
rect 11592 -2968 11678 -2957
rect 11592 -2973 11626 -2968
rect 11480 -3050 11496 -3016
rect 11564 -3050 11580 -3016
rect 11300 -3154 11334 -3092
rect 13971 -1963 14005 -1919
rect 14135 -1964 14169 -1819
rect 14203 -1788 14245 -1768
rect 14515 -1779 14549 -1733
rect 14868 -1767 14897 -1733
rect 14931 -1767 14989 -1733
rect 15023 -1767 15081 -1733
rect 15115 -1767 15173 -1733
rect 15207 -1767 15265 -1733
rect 15299 -1767 15357 -1733
rect 15391 -1767 15449 -1733
rect 15483 -1767 15541 -1733
rect 15575 -1767 15633 -1733
rect 15667 -1767 15725 -1733
rect 15759 -1767 15817 -1733
rect 15851 -1767 15909 -1733
rect 15943 -1767 16001 -1733
rect 16035 -1767 16093 -1733
rect 16127 -1767 16185 -1733
rect 16219 -1767 16277 -1733
rect 16311 -1767 16369 -1733
rect 16403 -1767 16461 -1733
rect 16495 -1767 16553 -1733
rect 16587 -1767 16645 -1733
rect 16679 -1767 16737 -1733
rect 16771 -1767 16829 -1733
rect 16863 -1767 16921 -1733
rect 16955 -1767 17013 -1733
rect 17047 -1767 17105 -1733
rect 17139 -1767 17197 -1733
rect 17231 -1767 17289 -1733
rect 17323 -1767 17381 -1733
rect 17415 -1767 17473 -1733
rect 17507 -1767 17565 -1733
rect 17599 -1767 17657 -1733
rect 17691 -1767 17749 -1733
rect 17783 -1767 17841 -1733
rect 17875 -1767 17933 -1733
rect 17967 -1767 18025 -1733
rect 18059 -1767 18117 -1733
rect 18151 -1767 18209 -1733
rect 18243 -1767 18301 -1733
rect 18335 -1767 18393 -1733
rect 18427 -1767 18485 -1733
rect 18519 -1767 18577 -1733
rect 18611 -1767 18669 -1733
rect 18703 -1767 18761 -1733
rect 18795 -1767 18853 -1733
rect 18887 -1767 18945 -1733
rect 18979 -1767 19037 -1733
rect 19071 -1767 19129 -1733
rect 19163 -1767 19221 -1733
rect 19255 -1767 19313 -1733
rect 19347 -1767 19405 -1733
rect 19439 -1767 19497 -1733
rect 19531 -1767 19589 -1733
rect 19623 -1767 19681 -1733
rect 19715 -1767 19773 -1733
rect 19807 -1767 19865 -1733
rect 19899 -1767 19957 -1733
rect 19991 -1767 20049 -1733
rect 20083 -1767 20141 -1733
rect 20175 -1767 20233 -1733
rect 20267 -1767 20325 -1733
rect 20359 -1767 20417 -1733
rect 20451 -1767 20509 -1733
rect 20543 -1767 20601 -1733
rect 20635 -1767 20693 -1733
rect 20727 -1767 20785 -1733
rect 20819 -1767 20877 -1733
rect 20911 -1767 20969 -1733
rect 21003 -1767 21061 -1733
rect 21095 -1767 21153 -1733
rect 21187 -1767 21245 -1733
rect 21279 -1767 21337 -1733
rect 21371 -1767 21429 -1733
rect 21463 -1767 21521 -1733
rect 21555 -1767 21613 -1733
rect 21647 -1767 21705 -1733
rect 21739 -1767 21797 -1733
rect 21831 -1767 21889 -1733
rect 21923 -1767 21981 -1733
rect 22015 -1767 22073 -1733
rect 22107 -1767 22136 -1733
rect 14237 -1822 14245 -1788
rect 14203 -1838 14245 -1822
rect 14279 -1819 14301 -1785
rect 14335 -1819 14431 -1785
rect 14465 -1819 14481 -1785
rect 14203 -1911 14204 -1872
rect 14203 -1960 14204 -1945
rect 14242 -1960 14243 -1872
rect 14203 -1961 14243 -1960
rect 13971 -2055 14005 -1997
rect 11726 -3154 11760 -3092
rect 11300 -3188 11396 -3154
rect 11664 -3188 11760 -3154
rect 12600 -2126 12696 -2092
rect 12952 -2126 13048 -2092
rect 12600 -2156 13048 -2126
rect 12600 -2188 12634 -2156
rect 12770 -2206 12878 -2156
rect 12770 -2240 12786 -2206
rect 12862 -2240 12878 -2206
rect 13014 -2188 13048 -2156
rect 12702 -2268 12736 -2252
rect 12702 -3052 12736 -3036
rect 12912 -2268 12946 -2252
rect 12912 -3052 12946 -3036
rect 12770 -3098 12786 -3064
rect 12862 -3098 12878 -3064
rect 12600 -3178 12634 -3116
rect 13971 -2147 14005 -2089
rect 13971 -2239 14005 -2181
rect 14039 -1998 14169 -1964
rect 14039 -2037 14089 -1998
rect 14203 -2011 14243 -1995
rect 14039 -2071 14055 -2037
rect 14039 -2141 14089 -2071
rect 14123 -2040 14203 -2034
rect 14123 -2074 14138 -2040
rect 14237 -2045 14243 -2011
rect 14230 -2074 14243 -2045
rect 14123 -2090 14243 -2074
rect 14039 -2175 14055 -2141
rect 14039 -2237 14089 -2175
rect 14123 -2156 14243 -2144
rect 14123 -2190 14136 -2156
rect 14228 -2160 14243 -2156
rect 14123 -2194 14203 -2190
rect 14237 -2194 14243 -2160
rect 14123 -2201 14243 -2194
rect 14203 -2210 14243 -2201
rect 14039 -2271 14169 -2237
rect 13971 -2305 14005 -2273
rect 13971 -2321 14101 -2305
rect 13971 -2331 14051 -2321
rect 14005 -2355 14051 -2331
rect 14085 -2355 14101 -2321
rect 14005 -2365 14101 -2355
rect 13971 -2371 14101 -2365
rect 14135 -2363 14169 -2271
rect 14203 -2250 14243 -2244
rect 14203 -2267 14204 -2250
rect 14203 -2317 14204 -2301
rect 14242 -2317 14243 -2250
rect 14279 -2363 14313 -1819
rect 14347 -1869 14481 -1853
rect 14347 -1903 14363 -1869
rect 14397 -1903 14431 -1869
rect 14465 -1903 14481 -1869
rect 14347 -1919 14481 -1903
rect 14347 -1987 14363 -1953
rect 14397 -1987 14413 -1953
rect 14347 -1999 14413 -1987
rect 14347 -2230 14395 -1999
rect 14447 -2021 14481 -1919
rect 14439 -2037 14481 -2021
rect 14473 -2071 14481 -2037
rect 14439 -2087 14481 -2071
rect 14515 -1871 14549 -1813
rect 14515 -1963 14549 -1905
rect 14885 -1861 14943 -1767
rect 15150 -1805 15238 -1767
rect 14885 -1895 14897 -1861
rect 14931 -1895 14943 -1861
rect 14885 -1912 14943 -1895
rect 14997 -1822 15058 -1806
rect 14997 -1856 15008 -1822
rect 15042 -1856 15058 -1822
rect 15150 -1839 15179 -1805
rect 15213 -1839 15238 -1805
rect 15150 -1855 15238 -1839
rect 15272 -1809 15403 -1801
rect 15272 -1843 15288 -1809
rect 15322 -1843 15403 -1809
rect 15272 -1855 15403 -1843
rect 14997 -1889 15058 -1856
rect 14997 -1919 15316 -1889
rect 14997 -1932 15266 -1919
rect 14997 -1940 15114 -1932
rect 14515 -2055 14549 -1997
rect 14977 -1988 15046 -1987
rect 14515 -2125 14549 -2089
rect 14431 -2141 14549 -2125
rect 14465 -2147 14549 -2141
rect 14465 -2175 14515 -2147
rect 14431 -2181 14515 -2175
rect 14431 -2196 14549 -2181
rect 14347 -2264 14361 -2230
rect 14395 -2264 14431 -2230
rect 14465 -2264 14481 -2230
rect 14347 -2280 14481 -2264
rect 14515 -2239 14549 -2196
rect 14515 -2314 14549 -2273
rect 13971 -2423 14005 -2371
rect 14135 -2397 14203 -2363
rect 14237 -2397 14313 -2363
rect 14363 -2330 14549 -2314
rect 14397 -2364 14431 -2330
rect 14465 -2331 14549 -2330
rect 14465 -2364 14515 -2331
rect 14363 -2365 14515 -2364
rect 14363 -2380 14549 -2365
rect 13048 -2468 13668 -2446
rect 13048 -3026 13052 -2468
rect 13648 -3026 13668 -2468
rect 13971 -2515 14005 -2457
rect 14039 -2448 14055 -2414
rect 14089 -2428 14105 -2414
rect 14089 -2431 14121 -2428
rect 14347 -2431 14363 -2414
rect 14089 -2448 14363 -2431
rect 14397 -2448 14431 -2414
rect 14465 -2448 14481 -2414
rect 14039 -2465 14481 -2448
rect 14515 -2423 14549 -2380
rect 14188 -2472 14332 -2465
rect 14188 -2503 14208 -2472
rect 13971 -2592 14005 -2549
rect 14039 -2524 14153 -2503
rect 14039 -2558 14060 -2524
rect 14094 -2558 14153 -2524
rect 13971 -2607 14085 -2592
rect 14005 -2617 14085 -2607
rect 14005 -2641 14043 -2617
rect 13971 -2651 14043 -2641
rect 14077 -2651 14085 -2617
rect 13971 -2684 14085 -2651
rect 14119 -2650 14153 -2558
rect 14187 -2554 14208 -2503
rect 14308 -2503 14332 -2472
rect 14187 -2588 14203 -2554
rect 14308 -2572 14333 -2503
rect 14237 -2588 14333 -2572
rect 14187 -2616 14333 -2588
rect 14367 -2524 14481 -2503
rect 14367 -2558 14426 -2524
rect 14460 -2558 14481 -2524
rect 14367 -2566 14481 -2558
rect 14515 -2515 14549 -2457
rect 14367 -2650 14401 -2566
rect 14515 -2600 14549 -2549
rect 14119 -2684 14203 -2650
rect 14237 -2684 14401 -2650
rect 14435 -2607 14549 -2600
rect 14435 -2618 14515 -2607
rect 14435 -2652 14443 -2618
rect 14477 -2641 14515 -2618
rect 14477 -2652 14549 -2641
rect 14435 -2684 14549 -2652
rect 13971 -2699 14005 -2684
rect 14515 -2699 14549 -2684
rect 13971 -2738 14005 -2733
rect 13918 -2754 14005 -2738
rect 13978 -2791 14005 -2754
rect 13918 -2825 13971 -2814
rect 13918 -2830 14005 -2825
rect 13971 -2854 14005 -2830
rect 14039 -2752 14481 -2718
rect 14039 -2783 14107 -2752
rect 14039 -2817 14055 -2783
rect 14089 -2817 14107 -2783
rect 14413 -2783 14481 -2752
rect 14039 -2837 14107 -2817
rect 14141 -2820 14203 -2786
rect 14237 -2820 14379 -2786
rect 14141 -2837 14379 -2820
rect 14413 -2817 14431 -2783
rect 14465 -2817 14481 -2783
rect 14413 -2837 14481 -2817
rect 14515 -2791 14549 -2733
rect 14040 -2888 14106 -2837
rect 14040 -2902 14140 -2888
rect 14212 -3016 14312 -2837
rect 14414 -2888 14480 -2837
rect 14515 -2854 14549 -2825
rect 14660 -2026 14826 -2012
rect 14660 -2098 14740 -2026
rect 14812 -2098 14826 -2026
rect 14660 -2112 14826 -2098
rect 14885 -2079 14943 -2044
rect 14660 -2476 14760 -2112
rect 14885 -2113 14897 -2079
rect 14931 -2113 14943 -2079
rect 14885 -2172 14943 -2113
rect 14977 -2140 14980 -1988
rect 15040 -2008 15046 -1988
rect 15040 -2076 15046 -2042
rect 15040 -2140 15046 -2110
rect 14977 -2141 15046 -2140
rect 14885 -2206 14897 -2172
rect 14931 -2206 14943 -2172
rect 15080 -2177 15114 -1940
rect 15250 -1953 15266 -1932
rect 15300 -1953 15316 -1919
rect 15148 -1969 15214 -1966
rect 15148 -1986 15164 -1969
rect 15198 -1986 15214 -1969
rect 15148 -2066 15160 -1986
rect 15200 -2066 15214 -1986
rect 15250 -1987 15316 -1953
rect 15250 -2021 15266 -1987
rect 15300 -2021 15316 -1987
rect 15250 -2037 15316 -2021
rect 15350 -1954 15403 -1855
rect 15437 -1861 15495 -1767
rect 15615 -1809 15681 -1767
rect 15437 -1895 15449 -1861
rect 15483 -1895 15495 -1861
rect 15437 -1912 15495 -1895
rect 15530 -1835 15581 -1819
rect 15530 -1869 15547 -1835
rect 15615 -1843 15631 -1809
rect 15665 -1843 15681 -1809
rect 15821 -1805 15887 -1767
rect 15715 -1835 15749 -1819
rect 15530 -1877 15581 -1869
rect 15821 -1839 15837 -1805
rect 15871 -1839 15887 -1805
rect 16407 -1809 16473 -1767
rect 15530 -1911 15680 -1877
rect 15530 -1954 15600 -1945
rect 15350 -1965 15600 -1954
rect 15350 -1999 15544 -1965
rect 15578 -1999 15600 -1965
rect 15350 -2004 15600 -1999
rect 15148 -2071 15164 -2066
rect 15198 -2071 15214 -2066
rect 15148 -2073 15214 -2071
rect 15350 -2117 15403 -2004
rect 15182 -2133 15284 -2117
rect 15182 -2167 15248 -2133
rect 15282 -2167 15284 -2133
rect 14885 -2277 14943 -2206
rect 14992 -2201 15046 -2185
rect 14992 -2235 15008 -2201
rect 15042 -2235 15046 -2201
rect 14992 -2277 15046 -2235
rect 15080 -2193 15133 -2177
rect 15080 -2227 15096 -2193
rect 15130 -2227 15133 -2193
rect 15080 -2243 15133 -2227
rect 15182 -2201 15284 -2167
rect 15216 -2235 15250 -2201
rect 15182 -2277 15284 -2235
rect 15318 -2133 15403 -2117
rect 15318 -2167 15336 -2133
rect 15370 -2167 15403 -2133
rect 15318 -2201 15403 -2167
rect 15318 -2235 15336 -2201
rect 15370 -2235 15403 -2201
rect 15318 -2243 15403 -2235
rect 15437 -2079 15495 -2044
rect 15530 -2075 15600 -2004
rect 15634 -1971 15680 -1911
rect 15668 -1980 15680 -1971
rect 15634 -2014 15646 -2005
rect 15437 -2113 15449 -2079
rect 15483 -2113 15495 -2079
rect 15634 -2109 15680 -2014
rect 15437 -2172 15495 -2113
rect 15437 -2206 15449 -2172
rect 15483 -2206 15495 -2172
rect 15437 -2277 15495 -2206
rect 15530 -2125 15680 -2109
rect 15530 -2159 15547 -2125
rect 15581 -2143 15680 -2125
rect 15715 -2107 15749 -1869
rect 15921 -1845 15970 -1811
rect 16004 -1845 16020 -1811
rect 16061 -1845 16077 -1811
rect 16111 -1845 16232 -1811
rect 15795 -2026 15887 -1873
rect 15795 -2036 15853 -2026
rect 15795 -2076 15814 -2036
rect 15854 -2076 15887 -2060
rect 15795 -2083 15887 -2076
rect 15530 -2193 15581 -2159
rect 15530 -2227 15547 -2193
rect 15530 -2243 15581 -2227
rect 15615 -2211 15631 -2177
rect 15665 -2211 15681 -2177
rect 15615 -2277 15681 -2211
rect 15715 -2193 15749 -2159
rect 15715 -2243 15749 -2227
rect 15783 -2240 15848 -2083
rect 15921 -2117 15955 -1845
rect 15989 -1919 16059 -1903
rect 15989 -1953 16012 -1919
rect 16046 -1953 16059 -1919
rect 15989 -1971 16059 -1953
rect 15989 -2005 16001 -1971
rect 16035 -2005 16059 -1971
rect 15989 -2027 16059 -2005
rect 16093 -1913 16164 -1903
rect 16093 -1947 16114 -1913
rect 16148 -1947 16164 -1913
rect 16093 -2065 16127 -1947
rect 16198 -1987 16232 -1845
rect 16407 -1843 16423 -1809
rect 16457 -1843 16473 -1809
rect 16407 -1859 16473 -1843
rect 16515 -1839 16535 -1805
rect 16569 -1839 16585 -1805
rect 16629 -1809 16819 -1801
rect 16307 -1937 16345 -1903
rect 16379 -1919 16431 -1903
rect 16515 -1917 16567 -1839
rect 16629 -1843 16645 -1809
rect 16679 -1843 16819 -1809
rect 16629 -1857 16819 -1843
rect 16853 -1805 16891 -1767
rect 16853 -1839 16857 -1805
rect 16853 -1855 16891 -1839
rect 16925 -1825 17139 -1809
rect 16925 -1843 17075 -1825
rect 16273 -1953 16369 -1937
rect 16403 -1953 16431 -1919
rect 16465 -1967 16499 -1951
rect 16034 -2081 16127 -2065
rect 16068 -2107 16127 -2081
rect 16068 -2115 16093 -2107
rect 15921 -2151 16000 -2117
rect 16034 -2141 16093 -2115
rect 16034 -2143 16127 -2141
rect 16161 -2001 16465 -1987
rect 16161 -2021 16499 -2001
rect 15966 -2177 16000 -2151
rect 16161 -2177 16195 -2021
rect 16533 -2055 16567 -1917
rect 16267 -2089 16283 -2055
rect 16317 -2089 16567 -2055
rect 16605 -1907 16647 -1891
rect 16605 -1941 16613 -1907
rect 16605 -2049 16647 -1941
rect 16681 -1955 16751 -1891
rect 16681 -1989 16709 -1955
rect 16743 -1971 16751 -1955
rect 16681 -2005 16717 -1989
rect 16681 -2015 16751 -2005
rect 16785 -2013 16819 -1857
rect 16925 -1889 16959 -1843
rect 17109 -1859 17139 -1825
rect 16853 -1923 16959 -1889
rect 16993 -1903 17041 -1877
rect 16853 -1929 16897 -1923
rect 16887 -1963 16897 -1929
rect 17027 -1937 17041 -1903
rect 16993 -1957 17041 -1937
rect 16853 -1979 16897 -1963
rect 16933 -1966 16949 -1957
rect 16983 -1991 17041 -1957
rect 16967 -2000 17041 -1991
rect 16785 -2047 16866 -2013
rect 16933 -2031 17041 -2000
rect 17075 -1914 17139 -1859
rect 17179 -1848 17213 -1767
rect 17179 -1904 17213 -1882
rect 17247 -1813 17313 -1805
rect 17247 -1847 17263 -1813
rect 17297 -1847 17313 -1813
rect 17247 -1881 17313 -1847
rect 17075 -1949 17140 -1914
rect 17247 -1915 17263 -1881
rect 17297 -1915 17313 -1881
rect 17075 -1965 17199 -1949
rect 17075 -1999 17149 -1965
rect 17183 -1999 17199 -1965
rect 17075 -2009 17199 -1999
rect 17110 -2015 17199 -2009
rect 16605 -2081 16740 -2049
rect 16832 -2065 16866 -2047
rect 16605 -2083 16748 -2081
rect 16533 -2117 16567 -2089
rect 16706 -2107 16748 -2083
rect 15882 -2201 15932 -2185
rect 15882 -2235 15898 -2201
rect 15882 -2277 15932 -2235
rect 15966 -2193 16016 -2177
rect 15966 -2227 15982 -2193
rect 15966 -2243 16016 -2227
rect 16059 -2199 16195 -2177
rect 16059 -2233 16075 -2199
rect 16109 -2233 16195 -2199
rect 16229 -2157 16444 -2123
rect 16533 -2151 16645 -2117
rect 16706 -2141 16717 -2107
rect 16782 -2115 16798 -2081
rect 16751 -2141 16798 -2115
rect 16832 -2099 17026 -2065
rect 17060 -2099 17076 -2065
rect 16229 -2175 16263 -2157
rect 16410 -2175 16444 -2157
rect 16229 -2225 16263 -2209
rect 16310 -2225 16326 -2191
rect 16360 -2225 16376 -2191
rect 16410 -2225 16444 -2209
rect 16503 -2201 16577 -2185
rect 16059 -2243 16195 -2233
rect 16310 -2277 16376 -2225
rect 16503 -2235 16523 -2201
rect 16557 -2235 16577 -2201
rect 16503 -2277 16577 -2235
rect 16611 -2193 16645 -2151
rect 16832 -2175 16866 -2099
rect 17110 -2133 17144 -2015
rect 17247 -2041 17313 -1915
rect 16611 -2243 16645 -2227
rect 16692 -2200 16866 -2175
rect 16984 -2167 17144 -2133
rect 17232 -2057 17313 -2041
rect 17266 -2091 17313 -2057
rect 17232 -2125 17313 -2091
rect 17266 -2159 17313 -2125
rect 16984 -2175 17018 -2167
rect 16692 -2234 16708 -2200
rect 16742 -2234 16866 -2200
rect 16692 -2243 16866 -2234
rect 16900 -2201 16950 -2185
rect 16934 -2235 16950 -2201
rect 17232 -2193 17313 -2159
rect 16984 -2225 17018 -2209
rect 16900 -2277 16950 -2235
rect 17054 -2235 17070 -2201
rect 17104 -2235 17148 -2201
rect 17182 -2235 17198 -2201
rect 17054 -2277 17198 -2235
rect 17266 -2227 17313 -2193
rect 17232 -2243 17313 -2227
rect 17351 -1835 17401 -1819
rect 17351 -1869 17367 -1835
rect 17351 -1949 17401 -1869
rect 17464 -1829 17498 -1767
rect 17464 -1886 17498 -1863
rect 17548 -1859 17599 -1803
rect 17582 -1893 17599 -1859
rect 17548 -1909 17599 -1893
rect 17351 -1965 17523 -1949
rect 17351 -1999 17489 -1965
rect 17351 -2015 17523 -1999
rect 17557 -1954 17599 -1909
rect 17645 -1861 17703 -1767
rect 17823 -1809 17889 -1767
rect 17645 -1895 17657 -1861
rect 17691 -1895 17703 -1861
rect 17645 -1912 17703 -1895
rect 17738 -1835 17789 -1819
rect 17738 -1869 17755 -1835
rect 17823 -1843 17839 -1809
rect 17873 -1843 17889 -1809
rect 18029 -1805 18095 -1767
rect 17923 -1835 17957 -1819
rect 17738 -1877 17789 -1869
rect 18029 -1839 18045 -1805
rect 18079 -1839 18095 -1805
rect 18615 -1809 18681 -1767
rect 17738 -1911 17888 -1877
rect 17738 -1954 17808 -1945
rect 17557 -1965 17808 -1954
rect 17557 -1999 17752 -1965
rect 17786 -1999 17808 -1965
rect 17557 -2004 17808 -1999
rect 17351 -2133 17417 -2015
rect 17557 -2039 17599 -2004
rect 17351 -2167 17367 -2133
rect 17401 -2167 17417 -2133
rect 17351 -2201 17417 -2167
rect 17351 -2235 17367 -2201
rect 17401 -2235 17417 -2201
rect 17464 -2065 17498 -2049
rect 17464 -2133 17498 -2099
rect 17464 -2201 17498 -2167
rect 17548 -2050 17599 -2039
rect 17548 -2088 17556 -2050
rect 17594 -2088 17599 -2050
rect 17548 -2097 17599 -2088
rect 17582 -2131 17599 -2097
rect 17548 -2165 17599 -2131
rect 17582 -2199 17599 -2165
rect 17548 -2215 17599 -2199
rect 17645 -2079 17703 -2044
rect 17738 -2075 17808 -2004
rect 17842 -1971 17888 -1911
rect 17876 -1980 17888 -1971
rect 17842 -2014 17854 -2005
rect 17645 -2113 17657 -2079
rect 17691 -2113 17703 -2079
rect 17842 -2109 17888 -2014
rect 17645 -2172 17703 -2113
rect 17645 -2206 17657 -2172
rect 17691 -2206 17703 -2172
rect 17464 -2277 17498 -2235
rect 17645 -2277 17703 -2206
rect 17738 -2125 17888 -2109
rect 17738 -2159 17755 -2125
rect 17789 -2143 17888 -2125
rect 17923 -2107 17957 -1869
rect 18129 -1845 18178 -1811
rect 18212 -1845 18228 -1811
rect 18269 -1845 18285 -1811
rect 18319 -1845 18440 -1811
rect 18003 -2026 18095 -1873
rect 18003 -2036 18061 -2026
rect 18003 -2076 18022 -2036
rect 18062 -2076 18095 -2060
rect 18003 -2083 18095 -2076
rect 17738 -2193 17789 -2159
rect 17738 -2227 17755 -2193
rect 17738 -2243 17789 -2227
rect 17823 -2211 17839 -2177
rect 17873 -2211 17889 -2177
rect 17823 -2277 17889 -2211
rect 17923 -2193 17957 -2159
rect 17923 -2243 17957 -2227
rect 17991 -2240 18056 -2083
rect 18129 -2117 18163 -1845
rect 18197 -1919 18267 -1903
rect 18197 -1953 18220 -1919
rect 18254 -1953 18267 -1919
rect 18197 -1971 18267 -1953
rect 18197 -2005 18209 -1971
rect 18243 -2005 18267 -1971
rect 18197 -2027 18267 -2005
rect 18301 -1913 18372 -1903
rect 18301 -1947 18322 -1913
rect 18356 -1947 18372 -1913
rect 18301 -2065 18335 -1947
rect 18406 -1987 18440 -1845
rect 18615 -1843 18631 -1809
rect 18665 -1843 18681 -1809
rect 18615 -1859 18681 -1843
rect 18723 -1839 18743 -1805
rect 18777 -1839 18793 -1805
rect 18837 -1809 19027 -1801
rect 18515 -1937 18553 -1903
rect 18587 -1919 18639 -1903
rect 18723 -1917 18775 -1839
rect 18837 -1843 18853 -1809
rect 18887 -1843 19027 -1809
rect 18837 -1857 19027 -1843
rect 19061 -1805 19099 -1767
rect 19061 -1839 19065 -1805
rect 19061 -1855 19099 -1839
rect 19133 -1825 19347 -1809
rect 19133 -1843 19283 -1825
rect 18481 -1953 18577 -1937
rect 18611 -1953 18639 -1919
rect 18673 -1967 18707 -1951
rect 18242 -2081 18335 -2065
rect 18276 -2107 18335 -2081
rect 18276 -2115 18301 -2107
rect 18129 -2151 18208 -2117
rect 18242 -2141 18301 -2115
rect 18242 -2143 18335 -2141
rect 18369 -2001 18673 -1987
rect 18369 -2021 18707 -2001
rect 18174 -2177 18208 -2151
rect 18369 -2177 18403 -2021
rect 18741 -2055 18775 -1917
rect 18475 -2089 18491 -2055
rect 18525 -2089 18775 -2055
rect 18813 -1907 18855 -1891
rect 18813 -1941 18821 -1907
rect 18813 -2049 18855 -1941
rect 18889 -1955 18959 -1891
rect 18889 -1989 18917 -1955
rect 18951 -1971 18959 -1955
rect 18889 -2005 18925 -1989
rect 18889 -2015 18959 -2005
rect 18993 -2013 19027 -1857
rect 19133 -1889 19167 -1843
rect 19317 -1859 19347 -1825
rect 19061 -1923 19167 -1889
rect 19201 -1903 19249 -1877
rect 19061 -1929 19105 -1923
rect 19095 -1963 19105 -1929
rect 19235 -1937 19249 -1903
rect 19201 -1957 19249 -1937
rect 19061 -1979 19105 -1963
rect 19141 -1966 19157 -1957
rect 19191 -1991 19249 -1957
rect 19175 -2000 19249 -1991
rect 18993 -2047 19074 -2013
rect 19141 -2031 19249 -2000
rect 19283 -1914 19347 -1859
rect 19387 -1848 19421 -1767
rect 19387 -1904 19421 -1882
rect 19455 -1813 19521 -1805
rect 19455 -1847 19471 -1813
rect 19505 -1847 19521 -1813
rect 19455 -1881 19521 -1847
rect 19283 -1949 19348 -1914
rect 19455 -1915 19471 -1881
rect 19505 -1915 19521 -1881
rect 19283 -1965 19407 -1949
rect 19283 -1999 19357 -1965
rect 19391 -1999 19407 -1965
rect 19283 -2009 19407 -1999
rect 19318 -2015 19407 -2009
rect 18813 -2081 18948 -2049
rect 19040 -2065 19074 -2047
rect 18813 -2083 18956 -2081
rect 18741 -2117 18775 -2089
rect 18914 -2107 18956 -2083
rect 18090 -2201 18140 -2185
rect 18090 -2235 18106 -2201
rect 18090 -2277 18140 -2235
rect 18174 -2193 18224 -2177
rect 18174 -2227 18190 -2193
rect 18174 -2243 18224 -2227
rect 18267 -2199 18403 -2177
rect 18267 -2233 18283 -2199
rect 18317 -2233 18403 -2199
rect 18437 -2157 18652 -2123
rect 18741 -2151 18853 -2117
rect 18914 -2141 18925 -2107
rect 18990 -2115 19006 -2081
rect 18959 -2141 19006 -2115
rect 19040 -2099 19234 -2065
rect 19268 -2099 19284 -2065
rect 18437 -2175 18471 -2157
rect 18618 -2175 18652 -2157
rect 18437 -2225 18471 -2209
rect 18518 -2225 18534 -2191
rect 18568 -2225 18584 -2191
rect 18618 -2225 18652 -2209
rect 18711 -2201 18785 -2185
rect 18267 -2243 18403 -2233
rect 18518 -2277 18584 -2225
rect 18711 -2235 18731 -2201
rect 18765 -2235 18785 -2201
rect 18711 -2277 18785 -2235
rect 18819 -2193 18853 -2151
rect 19040 -2175 19074 -2099
rect 19318 -2133 19352 -2015
rect 19455 -2041 19521 -1915
rect 18819 -2243 18853 -2227
rect 18900 -2200 19074 -2175
rect 19192 -2167 19352 -2133
rect 19440 -2057 19521 -2041
rect 19474 -2091 19521 -2057
rect 19440 -2125 19521 -2091
rect 19474 -2159 19521 -2125
rect 19192 -2175 19226 -2167
rect 18900 -2234 18916 -2200
rect 18950 -2234 19074 -2200
rect 18900 -2243 19074 -2234
rect 19108 -2201 19158 -2185
rect 19142 -2235 19158 -2201
rect 19440 -2193 19521 -2159
rect 19192 -2225 19226 -2209
rect 19108 -2277 19158 -2235
rect 19262 -2235 19278 -2201
rect 19312 -2235 19356 -2201
rect 19390 -2235 19406 -2201
rect 19262 -2277 19406 -2235
rect 19474 -2227 19521 -2193
rect 19440 -2243 19521 -2227
rect 19559 -1835 19609 -1819
rect 19559 -1869 19575 -1835
rect 19559 -1949 19609 -1869
rect 19672 -1829 19706 -1767
rect 19672 -1886 19706 -1863
rect 19756 -1859 19807 -1803
rect 19790 -1893 19807 -1859
rect 19756 -1909 19807 -1893
rect 19559 -1965 19731 -1949
rect 19559 -1999 19697 -1965
rect 19559 -2015 19731 -1999
rect 19765 -1954 19807 -1909
rect 19853 -1861 19911 -1767
rect 20031 -1809 20097 -1767
rect 19853 -1895 19865 -1861
rect 19899 -1895 19911 -1861
rect 19853 -1912 19911 -1895
rect 19946 -1835 19997 -1819
rect 19946 -1869 19963 -1835
rect 20031 -1843 20047 -1809
rect 20081 -1843 20097 -1809
rect 20237 -1805 20303 -1767
rect 20131 -1835 20165 -1819
rect 19946 -1877 19997 -1869
rect 20237 -1839 20253 -1805
rect 20287 -1839 20303 -1805
rect 20823 -1809 20889 -1767
rect 19946 -1911 20096 -1877
rect 19946 -1954 20016 -1945
rect 19765 -1965 20016 -1954
rect 19765 -1999 19960 -1965
rect 19994 -1999 20016 -1965
rect 19765 -2004 20016 -1999
rect 19559 -2133 19625 -2015
rect 19765 -2039 19807 -2004
rect 19559 -2167 19575 -2133
rect 19609 -2167 19625 -2133
rect 19559 -2201 19625 -2167
rect 19559 -2235 19575 -2201
rect 19609 -2235 19625 -2201
rect 19672 -2065 19706 -2049
rect 19672 -2133 19706 -2099
rect 19672 -2201 19706 -2167
rect 19756 -2050 19807 -2039
rect 19756 -2088 19766 -2050
rect 19804 -2088 19807 -2050
rect 19756 -2097 19807 -2088
rect 19790 -2131 19807 -2097
rect 19756 -2165 19807 -2131
rect 19790 -2199 19807 -2165
rect 19756 -2215 19807 -2199
rect 19853 -2079 19911 -2044
rect 19946 -2075 20016 -2004
rect 20050 -1971 20096 -1911
rect 20084 -1980 20096 -1971
rect 20050 -2014 20062 -2005
rect 19853 -2113 19865 -2079
rect 19899 -2113 19911 -2079
rect 20050 -2109 20096 -2014
rect 19853 -2172 19911 -2113
rect 19853 -2206 19865 -2172
rect 19899 -2206 19911 -2172
rect 19672 -2277 19706 -2235
rect 19853 -2277 19911 -2206
rect 19946 -2125 20096 -2109
rect 19946 -2159 19963 -2125
rect 19997 -2143 20096 -2125
rect 20131 -2107 20165 -1869
rect 20337 -1845 20386 -1811
rect 20420 -1845 20436 -1811
rect 20477 -1845 20493 -1811
rect 20527 -1845 20648 -1811
rect 20211 -2026 20303 -1873
rect 20211 -2036 20269 -2026
rect 20211 -2076 20230 -2036
rect 20270 -2076 20303 -2060
rect 20211 -2083 20303 -2076
rect 19946 -2193 19997 -2159
rect 19946 -2227 19963 -2193
rect 19946 -2243 19997 -2227
rect 20031 -2211 20047 -2177
rect 20081 -2211 20097 -2177
rect 20031 -2277 20097 -2211
rect 20131 -2193 20165 -2159
rect 20131 -2243 20165 -2227
rect 20199 -2240 20264 -2083
rect 20337 -2117 20371 -1845
rect 20405 -1919 20475 -1903
rect 20405 -1953 20428 -1919
rect 20462 -1953 20475 -1919
rect 20405 -1971 20475 -1953
rect 20405 -2005 20417 -1971
rect 20451 -2005 20475 -1971
rect 20405 -2027 20475 -2005
rect 20509 -1913 20580 -1903
rect 20509 -1947 20530 -1913
rect 20564 -1947 20580 -1913
rect 20509 -2065 20543 -1947
rect 20614 -1987 20648 -1845
rect 20823 -1843 20839 -1809
rect 20873 -1843 20889 -1809
rect 20823 -1859 20889 -1843
rect 20931 -1839 20951 -1805
rect 20985 -1839 21001 -1805
rect 21045 -1809 21235 -1801
rect 20723 -1937 20761 -1903
rect 20795 -1919 20847 -1903
rect 20931 -1917 20983 -1839
rect 21045 -1843 21061 -1809
rect 21095 -1843 21235 -1809
rect 21045 -1857 21235 -1843
rect 21269 -1805 21307 -1767
rect 21269 -1839 21273 -1805
rect 21269 -1855 21307 -1839
rect 21341 -1825 21555 -1809
rect 21341 -1843 21491 -1825
rect 20689 -1953 20785 -1937
rect 20819 -1953 20847 -1919
rect 20881 -1967 20915 -1951
rect 20450 -2081 20543 -2065
rect 20484 -2107 20543 -2081
rect 20484 -2115 20509 -2107
rect 20337 -2151 20416 -2117
rect 20450 -2141 20509 -2115
rect 20450 -2143 20543 -2141
rect 20577 -2001 20881 -1987
rect 20577 -2021 20915 -2001
rect 20382 -2177 20416 -2151
rect 20577 -2177 20611 -2021
rect 20949 -2055 20983 -1917
rect 20683 -2089 20699 -2055
rect 20733 -2089 20983 -2055
rect 21021 -1907 21063 -1891
rect 21021 -1941 21029 -1907
rect 21021 -2049 21063 -1941
rect 21097 -1955 21167 -1891
rect 21097 -1989 21125 -1955
rect 21159 -1971 21167 -1955
rect 21097 -2005 21133 -1989
rect 21097 -2015 21167 -2005
rect 21201 -2013 21235 -1857
rect 21341 -1889 21375 -1843
rect 21525 -1859 21555 -1825
rect 21269 -1923 21375 -1889
rect 21409 -1903 21457 -1877
rect 21269 -1929 21313 -1923
rect 21303 -1963 21313 -1929
rect 21443 -1937 21457 -1903
rect 21409 -1957 21457 -1937
rect 21269 -1979 21313 -1963
rect 21349 -1966 21365 -1957
rect 21399 -1991 21457 -1957
rect 21383 -2000 21457 -1991
rect 21201 -2047 21282 -2013
rect 21349 -2031 21457 -2000
rect 21491 -1914 21555 -1859
rect 21595 -1848 21629 -1767
rect 21595 -1904 21629 -1882
rect 21663 -1813 21729 -1805
rect 21663 -1847 21679 -1813
rect 21713 -1847 21729 -1813
rect 21663 -1881 21729 -1847
rect 21491 -1949 21556 -1914
rect 21663 -1915 21679 -1881
rect 21713 -1915 21729 -1881
rect 21491 -1965 21615 -1949
rect 21491 -1999 21565 -1965
rect 21599 -1999 21615 -1965
rect 21491 -2009 21615 -1999
rect 21526 -2015 21615 -2009
rect 21021 -2081 21156 -2049
rect 21248 -2065 21282 -2047
rect 21021 -2083 21164 -2081
rect 20949 -2117 20983 -2089
rect 21122 -2107 21164 -2083
rect 20298 -2201 20348 -2185
rect 20298 -2235 20314 -2201
rect 20298 -2277 20348 -2235
rect 20382 -2193 20432 -2177
rect 20382 -2227 20398 -2193
rect 20382 -2243 20432 -2227
rect 20475 -2199 20611 -2177
rect 20475 -2233 20491 -2199
rect 20525 -2233 20611 -2199
rect 20645 -2157 20860 -2123
rect 20949 -2151 21061 -2117
rect 21122 -2141 21133 -2107
rect 21198 -2115 21214 -2081
rect 21167 -2141 21214 -2115
rect 21248 -2099 21442 -2065
rect 21476 -2099 21492 -2065
rect 20645 -2175 20679 -2157
rect 20826 -2175 20860 -2157
rect 20645 -2225 20679 -2209
rect 20726 -2225 20742 -2191
rect 20776 -2225 20792 -2191
rect 20826 -2225 20860 -2209
rect 20919 -2201 20993 -2185
rect 20475 -2243 20611 -2233
rect 20726 -2277 20792 -2225
rect 20919 -2235 20939 -2201
rect 20973 -2235 20993 -2201
rect 20919 -2277 20993 -2235
rect 21027 -2193 21061 -2151
rect 21248 -2175 21282 -2099
rect 21526 -2133 21560 -2015
rect 21663 -2041 21729 -1915
rect 21027 -2243 21061 -2227
rect 21108 -2200 21282 -2175
rect 21400 -2167 21560 -2133
rect 21648 -2057 21729 -2041
rect 21682 -2091 21729 -2057
rect 21648 -2125 21729 -2091
rect 21682 -2159 21729 -2125
rect 21400 -2175 21434 -2167
rect 21108 -2234 21124 -2200
rect 21158 -2234 21282 -2200
rect 21108 -2243 21282 -2234
rect 21316 -2201 21366 -2185
rect 21350 -2235 21366 -2201
rect 21648 -2193 21729 -2159
rect 21400 -2225 21434 -2209
rect 21316 -2277 21366 -2235
rect 21470 -2235 21486 -2201
rect 21520 -2235 21564 -2201
rect 21598 -2235 21614 -2201
rect 21470 -2277 21614 -2235
rect 21682 -2227 21729 -2193
rect 21648 -2243 21729 -2227
rect 21767 -1835 21817 -1819
rect 21767 -1869 21783 -1835
rect 21767 -1949 21817 -1869
rect 21880 -1829 21914 -1767
rect 21880 -1886 21914 -1863
rect 21964 -1859 22015 -1803
rect 21998 -1893 22015 -1859
rect 21964 -1909 22015 -1893
rect 21767 -1965 21939 -1949
rect 21767 -1999 21905 -1965
rect 21767 -2015 21939 -1999
rect 21973 -1966 22015 -1909
rect 22061 -1861 22119 -1767
rect 22061 -1895 22073 -1861
rect 22107 -1895 22119 -1861
rect 22061 -1912 22119 -1895
rect 21767 -2133 21833 -2015
rect 21973 -2039 21974 -1966
rect 21767 -2167 21783 -2133
rect 21817 -2167 21833 -2133
rect 21767 -2201 21833 -2167
rect 21767 -2235 21783 -2201
rect 21817 -2235 21833 -2201
rect 21880 -2065 21914 -2049
rect 21880 -2133 21914 -2099
rect 21880 -2201 21914 -2167
rect 21964 -2097 21974 -2039
rect 21964 -2160 21974 -2131
rect 22014 -2160 22015 -1966
rect 21964 -2165 22015 -2160
rect 21998 -2199 22015 -2165
rect 21964 -2215 22015 -2199
rect 22061 -2079 22119 -2044
rect 22061 -2113 22073 -2079
rect 22107 -2113 22119 -2079
rect 22061 -2172 22119 -2113
rect 22061 -2206 22073 -2172
rect 22107 -2206 22119 -2172
rect 21880 -2277 21914 -2235
rect 22061 -2277 22119 -2206
rect 14868 -2311 14897 -2277
rect 14931 -2311 14989 -2277
rect 15023 -2311 15081 -2277
rect 15115 -2311 15173 -2277
rect 15207 -2311 15265 -2277
rect 15299 -2311 15357 -2277
rect 15391 -2311 15449 -2277
rect 15483 -2311 15541 -2277
rect 15575 -2311 15633 -2277
rect 15667 -2311 15725 -2277
rect 15759 -2311 15817 -2277
rect 15851 -2311 15909 -2277
rect 15943 -2311 16001 -2277
rect 16035 -2311 16093 -2277
rect 16127 -2311 16185 -2277
rect 16219 -2311 16277 -2277
rect 16311 -2311 16369 -2277
rect 16403 -2311 16461 -2277
rect 16495 -2311 16553 -2277
rect 16587 -2311 16645 -2277
rect 16679 -2311 16737 -2277
rect 16771 -2311 16829 -2277
rect 16863 -2311 16921 -2277
rect 16955 -2311 17013 -2277
rect 17047 -2311 17105 -2277
rect 17139 -2311 17197 -2277
rect 17231 -2311 17289 -2277
rect 17323 -2311 17381 -2277
rect 17415 -2311 17473 -2277
rect 17507 -2311 17565 -2277
rect 17599 -2311 17657 -2277
rect 17691 -2311 17749 -2277
rect 17783 -2311 17841 -2277
rect 17875 -2311 17933 -2277
rect 17967 -2311 18025 -2277
rect 18059 -2311 18117 -2277
rect 18151 -2311 18209 -2277
rect 18243 -2311 18301 -2277
rect 18335 -2311 18393 -2277
rect 18427 -2311 18485 -2277
rect 18519 -2311 18577 -2277
rect 18611 -2311 18669 -2277
rect 18703 -2311 18761 -2277
rect 18795 -2311 18853 -2277
rect 18887 -2311 18945 -2277
rect 18979 -2311 19037 -2277
rect 19071 -2311 19129 -2277
rect 19163 -2311 19221 -2277
rect 19255 -2311 19313 -2277
rect 19347 -2311 19405 -2277
rect 19439 -2311 19497 -2277
rect 19531 -2311 19589 -2277
rect 19623 -2311 19681 -2277
rect 19715 -2311 19773 -2277
rect 19807 -2311 19865 -2277
rect 19899 -2311 19957 -2277
rect 19991 -2311 20049 -2277
rect 20083 -2311 20141 -2277
rect 20175 -2311 20233 -2277
rect 20267 -2311 20325 -2277
rect 20359 -2311 20417 -2277
rect 20451 -2311 20509 -2277
rect 20543 -2311 20601 -2277
rect 20635 -2311 20693 -2277
rect 20727 -2311 20785 -2277
rect 20819 -2311 20877 -2277
rect 20911 -2311 20969 -2277
rect 21003 -2311 21061 -2277
rect 21095 -2311 21153 -2277
rect 21187 -2311 21245 -2277
rect 21279 -2311 21337 -2277
rect 21371 -2311 21429 -2277
rect 21463 -2311 21521 -2277
rect 21555 -2311 21613 -2277
rect 21647 -2311 21705 -2277
rect 21739 -2311 21797 -2277
rect 21831 -2311 21889 -2277
rect 21923 -2311 21981 -2277
rect 22015 -2311 22073 -2277
rect 22107 -2311 22136 -2277
rect 14885 -2382 14943 -2311
rect 14885 -2416 14897 -2382
rect 14931 -2416 14943 -2382
rect 14992 -2353 15046 -2311
rect 14992 -2387 15008 -2353
rect 15042 -2387 15046 -2353
rect 14992 -2403 15046 -2387
rect 15080 -2361 15133 -2345
rect 15080 -2395 15096 -2361
rect 15130 -2395 15133 -2361
rect 14885 -2475 14943 -2416
rect 15080 -2411 15133 -2395
rect 15182 -2353 15284 -2311
rect 15216 -2387 15250 -2353
rect 14660 -2490 14826 -2476
rect 14660 -2562 14740 -2490
rect 14812 -2562 14826 -2490
rect 14885 -2509 14897 -2475
rect 14931 -2509 14943 -2475
rect 14885 -2544 14943 -2509
rect 14977 -2448 15046 -2447
rect 14660 -2576 14826 -2562
rect 14414 -2902 14514 -2888
rect 14660 -3016 14760 -2576
rect 14977 -2600 14980 -2448
rect 15040 -2478 15046 -2448
rect 15040 -2546 15046 -2512
rect 15040 -2600 15046 -2580
rect 14977 -2601 15046 -2600
rect 15080 -2648 15114 -2411
rect 15182 -2421 15284 -2387
rect 15182 -2455 15248 -2421
rect 15282 -2455 15284 -2421
rect 15182 -2471 15284 -2455
rect 15318 -2353 15403 -2345
rect 15318 -2387 15336 -2353
rect 15370 -2387 15403 -2353
rect 15318 -2421 15403 -2387
rect 15318 -2455 15336 -2421
rect 15370 -2455 15403 -2421
rect 15318 -2471 15403 -2455
rect 15148 -2517 15214 -2515
rect 15148 -2522 15164 -2517
rect 15198 -2522 15214 -2517
rect 15148 -2602 15160 -2522
rect 15200 -2602 15214 -2522
rect 15148 -2619 15164 -2602
rect 15198 -2619 15214 -2602
rect 15148 -2622 15214 -2619
rect 15250 -2567 15316 -2551
rect 15250 -2601 15266 -2567
rect 15300 -2601 15316 -2567
rect 14997 -2656 15114 -2648
rect 15250 -2635 15316 -2601
rect 15250 -2656 15266 -2635
rect 14997 -2669 15266 -2656
rect 15300 -2669 15316 -2635
rect 14885 -2693 14943 -2676
rect 14885 -2727 14897 -2693
rect 14931 -2727 14943 -2693
rect 14885 -2821 14943 -2727
rect 14997 -2699 15316 -2669
rect 15350 -2584 15403 -2471
rect 15437 -2382 15495 -2311
rect 15437 -2416 15449 -2382
rect 15483 -2416 15495 -2382
rect 15437 -2475 15495 -2416
rect 15437 -2509 15449 -2475
rect 15483 -2509 15495 -2475
rect 15530 -2361 15581 -2345
rect 15530 -2395 15547 -2361
rect 15530 -2429 15581 -2395
rect 15615 -2377 15681 -2311
rect 15615 -2411 15631 -2377
rect 15665 -2411 15681 -2377
rect 15715 -2361 15749 -2345
rect 15530 -2463 15547 -2429
rect 15715 -2429 15749 -2395
rect 15581 -2463 15680 -2445
rect 15530 -2479 15680 -2463
rect 15437 -2544 15495 -2509
rect 15530 -2584 15600 -2513
rect 15350 -2589 15600 -2584
rect 15350 -2623 15544 -2589
rect 15578 -2623 15600 -2589
rect 15350 -2634 15600 -2623
rect 14997 -2732 15058 -2699
rect 14997 -2766 15008 -2732
rect 15042 -2766 15058 -2732
rect 15350 -2733 15403 -2634
rect 15530 -2643 15600 -2634
rect 15634 -2574 15680 -2479
rect 15634 -2583 15646 -2574
rect 15668 -2617 15680 -2608
rect 14997 -2782 15058 -2766
rect 15150 -2749 15238 -2733
rect 15150 -2783 15179 -2749
rect 15213 -2783 15238 -2749
rect 15150 -2821 15238 -2783
rect 15272 -2745 15403 -2733
rect 15272 -2779 15288 -2745
rect 15322 -2779 15403 -2745
rect 15272 -2787 15403 -2779
rect 15437 -2693 15495 -2676
rect 15634 -2677 15680 -2617
rect 15437 -2727 15449 -2693
rect 15483 -2727 15495 -2693
rect 15437 -2821 15495 -2727
rect 15530 -2711 15680 -2677
rect 15530 -2719 15581 -2711
rect 15530 -2753 15547 -2719
rect 15715 -2719 15749 -2481
rect 15783 -2505 15848 -2348
rect 15882 -2353 15932 -2311
rect 15882 -2387 15898 -2353
rect 15882 -2403 15932 -2387
rect 15966 -2361 16016 -2345
rect 15966 -2395 15982 -2361
rect 15966 -2411 16016 -2395
rect 16059 -2355 16195 -2345
rect 16059 -2389 16075 -2355
rect 16109 -2389 16195 -2355
rect 16310 -2363 16376 -2311
rect 16503 -2353 16577 -2311
rect 16059 -2411 16195 -2389
rect 15966 -2437 16000 -2411
rect 15921 -2471 16000 -2437
rect 16034 -2447 16127 -2445
rect 15795 -2512 15887 -2505
rect 15795 -2552 15814 -2512
rect 15854 -2528 15887 -2512
rect 15795 -2562 15853 -2552
rect 15795 -2715 15887 -2562
rect 15530 -2769 15581 -2753
rect 15615 -2779 15631 -2745
rect 15665 -2779 15681 -2745
rect 15921 -2743 15955 -2471
rect 16034 -2473 16093 -2447
rect 16068 -2481 16093 -2473
rect 16068 -2507 16127 -2481
rect 16034 -2523 16127 -2507
rect 15989 -2583 16059 -2561
rect 15989 -2617 16001 -2583
rect 16035 -2617 16059 -2583
rect 15989 -2635 16059 -2617
rect 15989 -2669 16012 -2635
rect 16046 -2669 16059 -2635
rect 15989 -2685 16059 -2669
rect 16093 -2641 16127 -2523
rect 16161 -2567 16195 -2411
rect 16229 -2379 16263 -2363
rect 16310 -2397 16326 -2363
rect 16360 -2397 16376 -2363
rect 16410 -2379 16444 -2363
rect 16229 -2431 16263 -2413
rect 16503 -2387 16523 -2353
rect 16557 -2387 16577 -2353
rect 16503 -2403 16577 -2387
rect 16611 -2361 16645 -2345
rect 16410 -2431 16444 -2413
rect 16229 -2465 16444 -2431
rect 16611 -2437 16645 -2395
rect 16692 -2354 16866 -2345
rect 16692 -2388 16708 -2354
rect 16742 -2388 16866 -2354
rect 16692 -2413 16866 -2388
rect 16900 -2353 16950 -2311
rect 16934 -2387 16950 -2353
rect 17054 -2353 17198 -2311
rect 16900 -2403 16950 -2387
rect 16984 -2379 17018 -2363
rect 16533 -2471 16645 -2437
rect 16533 -2499 16567 -2471
rect 16267 -2533 16283 -2499
rect 16317 -2533 16567 -2499
rect 16706 -2481 16717 -2447
rect 16751 -2473 16798 -2447
rect 16706 -2505 16748 -2481
rect 16161 -2587 16499 -2567
rect 16161 -2601 16465 -2587
rect 16093 -2675 16114 -2641
rect 16148 -2675 16164 -2641
rect 16093 -2685 16164 -2675
rect 16198 -2743 16232 -2601
rect 16273 -2651 16369 -2635
rect 16307 -2685 16345 -2651
rect 16403 -2669 16431 -2635
rect 16465 -2637 16499 -2621
rect 16379 -2685 16431 -2669
rect 16533 -2671 16567 -2533
rect 15715 -2769 15749 -2753
rect 15615 -2821 15681 -2779
rect 15821 -2783 15837 -2749
rect 15871 -2783 15887 -2749
rect 15921 -2777 15970 -2743
rect 16004 -2777 16020 -2743
rect 16061 -2777 16077 -2743
rect 16111 -2777 16232 -2743
rect 16407 -2745 16473 -2729
rect 15821 -2821 15887 -2783
rect 16407 -2779 16423 -2745
rect 16457 -2779 16473 -2745
rect 16407 -2821 16473 -2779
rect 16515 -2749 16567 -2671
rect 16605 -2507 16748 -2505
rect 16782 -2507 16798 -2473
rect 16832 -2489 16866 -2413
rect 17054 -2387 17070 -2353
rect 17104 -2387 17148 -2353
rect 17182 -2387 17198 -2353
rect 17232 -2361 17313 -2345
rect 17464 -2353 17498 -2311
rect 16984 -2421 17018 -2413
rect 17266 -2395 17313 -2361
rect 16984 -2455 17144 -2421
rect 16605 -2539 16740 -2507
rect 16832 -2523 17026 -2489
rect 17060 -2523 17076 -2489
rect 16605 -2647 16647 -2539
rect 16832 -2541 16866 -2523
rect 16605 -2681 16613 -2647
rect 16605 -2697 16647 -2681
rect 16681 -2583 16751 -2573
rect 16681 -2599 16717 -2583
rect 16681 -2633 16709 -2599
rect 16743 -2633 16751 -2617
rect 16681 -2697 16751 -2633
rect 16785 -2575 16866 -2541
rect 16785 -2731 16819 -2575
rect 16933 -2588 17041 -2557
rect 17110 -2573 17144 -2455
rect 17232 -2429 17313 -2395
rect 17266 -2463 17313 -2429
rect 17232 -2497 17313 -2463
rect 17266 -2531 17313 -2497
rect 17232 -2547 17313 -2531
rect 17110 -2579 17199 -2573
rect 16967 -2597 17041 -2588
rect 16853 -2625 16897 -2609
rect 16887 -2659 16897 -2625
rect 16933 -2631 16949 -2622
rect 16983 -2631 17041 -2597
rect 16853 -2665 16897 -2659
rect 16993 -2651 17041 -2631
rect 16853 -2699 16959 -2665
rect 16629 -2745 16819 -2731
rect 16515 -2783 16535 -2749
rect 16569 -2783 16585 -2749
rect 16629 -2779 16645 -2745
rect 16679 -2779 16819 -2745
rect 16629 -2787 16819 -2779
rect 16853 -2749 16891 -2733
rect 16853 -2783 16857 -2749
rect 16925 -2745 16959 -2699
rect 17027 -2685 17041 -2651
rect 16993 -2711 17041 -2685
rect 17075 -2589 17199 -2579
rect 17075 -2623 17149 -2589
rect 17183 -2623 17199 -2589
rect 17075 -2639 17199 -2623
rect 17075 -2674 17140 -2639
rect 17247 -2673 17313 -2547
rect 17075 -2729 17139 -2674
rect 16925 -2763 17075 -2745
rect 17109 -2763 17139 -2729
rect 16925 -2779 17139 -2763
rect 17179 -2706 17213 -2684
rect 16853 -2821 16891 -2783
rect 17179 -2821 17213 -2740
rect 17247 -2707 17263 -2673
rect 17297 -2707 17313 -2673
rect 17247 -2741 17313 -2707
rect 17247 -2775 17263 -2741
rect 17297 -2775 17313 -2741
rect 17351 -2387 17367 -2353
rect 17401 -2387 17417 -2353
rect 17351 -2421 17417 -2387
rect 17351 -2455 17367 -2421
rect 17401 -2455 17417 -2421
rect 17351 -2573 17417 -2455
rect 17464 -2421 17498 -2387
rect 17464 -2489 17498 -2455
rect 17464 -2539 17498 -2523
rect 17548 -2389 17599 -2373
rect 17582 -2423 17599 -2389
rect 17548 -2457 17599 -2423
rect 17582 -2491 17599 -2457
rect 17548 -2500 17599 -2491
rect 17548 -2538 17556 -2500
rect 17594 -2538 17599 -2500
rect 17548 -2549 17599 -2538
rect 17645 -2382 17703 -2311
rect 17645 -2416 17657 -2382
rect 17691 -2416 17703 -2382
rect 17645 -2475 17703 -2416
rect 17645 -2509 17657 -2475
rect 17691 -2509 17703 -2475
rect 17738 -2361 17789 -2345
rect 17738 -2395 17755 -2361
rect 17738 -2429 17789 -2395
rect 17823 -2377 17889 -2311
rect 17823 -2411 17839 -2377
rect 17873 -2411 17889 -2377
rect 17923 -2361 17957 -2345
rect 17738 -2463 17755 -2429
rect 17923 -2429 17957 -2395
rect 17789 -2463 17888 -2445
rect 17738 -2479 17888 -2463
rect 17645 -2544 17703 -2509
rect 17351 -2589 17523 -2573
rect 17351 -2623 17489 -2589
rect 17351 -2639 17523 -2623
rect 17557 -2584 17599 -2549
rect 17738 -2584 17808 -2513
rect 17557 -2589 17808 -2584
rect 17557 -2623 17752 -2589
rect 17786 -2623 17808 -2589
rect 17557 -2634 17808 -2623
rect 17351 -2719 17401 -2639
rect 17557 -2679 17599 -2634
rect 17738 -2643 17808 -2634
rect 17842 -2574 17888 -2479
rect 17842 -2583 17854 -2574
rect 17876 -2617 17888 -2608
rect 17548 -2695 17599 -2679
rect 17351 -2753 17367 -2719
rect 17351 -2769 17401 -2753
rect 17464 -2725 17498 -2702
rect 17247 -2783 17313 -2775
rect 17464 -2821 17498 -2759
rect 17582 -2729 17599 -2695
rect 17548 -2785 17599 -2729
rect 17645 -2693 17703 -2676
rect 17842 -2677 17888 -2617
rect 17645 -2727 17657 -2693
rect 17691 -2727 17703 -2693
rect 17645 -2821 17703 -2727
rect 17738 -2711 17888 -2677
rect 17738 -2719 17789 -2711
rect 17738 -2753 17755 -2719
rect 17923 -2719 17957 -2481
rect 17991 -2505 18056 -2348
rect 18090 -2353 18140 -2311
rect 18090 -2387 18106 -2353
rect 18090 -2403 18140 -2387
rect 18174 -2361 18224 -2345
rect 18174 -2395 18190 -2361
rect 18174 -2411 18224 -2395
rect 18267 -2355 18403 -2345
rect 18267 -2389 18283 -2355
rect 18317 -2389 18403 -2355
rect 18518 -2363 18584 -2311
rect 18711 -2353 18785 -2311
rect 18267 -2411 18403 -2389
rect 18174 -2437 18208 -2411
rect 18129 -2471 18208 -2437
rect 18242 -2447 18335 -2445
rect 18003 -2512 18095 -2505
rect 18003 -2552 18022 -2512
rect 18062 -2528 18095 -2512
rect 18003 -2562 18061 -2552
rect 18003 -2715 18095 -2562
rect 17738 -2769 17789 -2753
rect 17823 -2779 17839 -2745
rect 17873 -2779 17889 -2745
rect 18129 -2743 18163 -2471
rect 18242 -2473 18301 -2447
rect 18276 -2481 18301 -2473
rect 18276 -2507 18335 -2481
rect 18242 -2523 18335 -2507
rect 18197 -2583 18267 -2561
rect 18197 -2617 18209 -2583
rect 18243 -2617 18267 -2583
rect 18197 -2635 18267 -2617
rect 18197 -2669 18220 -2635
rect 18254 -2669 18267 -2635
rect 18197 -2685 18267 -2669
rect 18301 -2641 18335 -2523
rect 18369 -2567 18403 -2411
rect 18437 -2379 18471 -2363
rect 18518 -2397 18534 -2363
rect 18568 -2397 18584 -2363
rect 18618 -2379 18652 -2363
rect 18437 -2431 18471 -2413
rect 18711 -2387 18731 -2353
rect 18765 -2387 18785 -2353
rect 18711 -2403 18785 -2387
rect 18819 -2361 18853 -2345
rect 18618 -2431 18652 -2413
rect 18437 -2465 18652 -2431
rect 18819 -2437 18853 -2395
rect 18900 -2354 19074 -2345
rect 18900 -2388 18916 -2354
rect 18950 -2388 19074 -2354
rect 18900 -2413 19074 -2388
rect 19108 -2353 19158 -2311
rect 19142 -2387 19158 -2353
rect 19262 -2353 19406 -2311
rect 19108 -2403 19158 -2387
rect 19192 -2379 19226 -2363
rect 18741 -2471 18853 -2437
rect 18741 -2499 18775 -2471
rect 18475 -2533 18491 -2499
rect 18525 -2533 18775 -2499
rect 18914 -2481 18925 -2447
rect 18959 -2473 19006 -2447
rect 18914 -2505 18956 -2481
rect 18369 -2587 18707 -2567
rect 18369 -2601 18673 -2587
rect 18301 -2675 18322 -2641
rect 18356 -2675 18372 -2641
rect 18301 -2685 18372 -2675
rect 18406 -2743 18440 -2601
rect 18481 -2651 18577 -2635
rect 18515 -2685 18553 -2651
rect 18611 -2669 18639 -2635
rect 18673 -2637 18707 -2621
rect 18587 -2685 18639 -2669
rect 18741 -2671 18775 -2533
rect 17923 -2769 17957 -2753
rect 17823 -2821 17889 -2779
rect 18029 -2783 18045 -2749
rect 18079 -2783 18095 -2749
rect 18129 -2777 18178 -2743
rect 18212 -2777 18228 -2743
rect 18269 -2777 18285 -2743
rect 18319 -2777 18440 -2743
rect 18615 -2745 18681 -2729
rect 18029 -2821 18095 -2783
rect 18615 -2779 18631 -2745
rect 18665 -2779 18681 -2745
rect 18615 -2821 18681 -2779
rect 18723 -2749 18775 -2671
rect 18813 -2507 18956 -2505
rect 18990 -2507 19006 -2473
rect 19040 -2489 19074 -2413
rect 19262 -2387 19278 -2353
rect 19312 -2387 19356 -2353
rect 19390 -2387 19406 -2353
rect 19440 -2361 19521 -2345
rect 19672 -2353 19706 -2311
rect 19192 -2421 19226 -2413
rect 19474 -2395 19521 -2361
rect 19192 -2455 19352 -2421
rect 18813 -2539 18948 -2507
rect 19040 -2523 19234 -2489
rect 19268 -2523 19284 -2489
rect 18813 -2647 18855 -2539
rect 19040 -2541 19074 -2523
rect 18813 -2681 18821 -2647
rect 18813 -2697 18855 -2681
rect 18889 -2583 18959 -2573
rect 18889 -2599 18925 -2583
rect 18889 -2633 18917 -2599
rect 18951 -2633 18959 -2617
rect 18889 -2697 18959 -2633
rect 18993 -2575 19074 -2541
rect 18993 -2731 19027 -2575
rect 19141 -2588 19249 -2557
rect 19318 -2573 19352 -2455
rect 19440 -2429 19521 -2395
rect 19474 -2463 19521 -2429
rect 19440 -2497 19521 -2463
rect 19474 -2531 19521 -2497
rect 19440 -2547 19521 -2531
rect 19318 -2579 19407 -2573
rect 19175 -2597 19249 -2588
rect 19061 -2625 19105 -2609
rect 19095 -2659 19105 -2625
rect 19141 -2631 19157 -2622
rect 19191 -2631 19249 -2597
rect 19061 -2665 19105 -2659
rect 19201 -2651 19249 -2631
rect 19061 -2699 19167 -2665
rect 18837 -2745 19027 -2731
rect 18723 -2783 18743 -2749
rect 18777 -2783 18793 -2749
rect 18837 -2779 18853 -2745
rect 18887 -2779 19027 -2745
rect 18837 -2787 19027 -2779
rect 19061 -2749 19099 -2733
rect 19061 -2783 19065 -2749
rect 19133 -2745 19167 -2699
rect 19235 -2685 19249 -2651
rect 19201 -2711 19249 -2685
rect 19283 -2589 19407 -2579
rect 19283 -2623 19357 -2589
rect 19391 -2623 19407 -2589
rect 19283 -2639 19407 -2623
rect 19283 -2674 19348 -2639
rect 19455 -2673 19521 -2547
rect 19283 -2729 19347 -2674
rect 19133 -2763 19283 -2745
rect 19317 -2763 19347 -2729
rect 19133 -2779 19347 -2763
rect 19387 -2706 19421 -2684
rect 19061 -2821 19099 -2783
rect 19387 -2821 19421 -2740
rect 19455 -2707 19471 -2673
rect 19505 -2707 19521 -2673
rect 19455 -2741 19521 -2707
rect 19455 -2775 19471 -2741
rect 19505 -2775 19521 -2741
rect 19559 -2387 19575 -2353
rect 19609 -2387 19625 -2353
rect 19559 -2421 19625 -2387
rect 19559 -2455 19575 -2421
rect 19609 -2455 19625 -2421
rect 19559 -2573 19625 -2455
rect 19672 -2421 19706 -2387
rect 19672 -2489 19706 -2455
rect 19672 -2539 19706 -2523
rect 19756 -2389 19807 -2373
rect 19790 -2423 19807 -2389
rect 19756 -2457 19807 -2423
rect 19790 -2491 19807 -2457
rect 19756 -2500 19807 -2491
rect 19756 -2538 19766 -2500
rect 19804 -2538 19807 -2500
rect 19756 -2549 19807 -2538
rect 19853 -2382 19911 -2311
rect 19853 -2416 19865 -2382
rect 19899 -2416 19911 -2382
rect 19853 -2475 19911 -2416
rect 19853 -2509 19865 -2475
rect 19899 -2509 19911 -2475
rect 19946 -2361 19997 -2345
rect 19946 -2395 19963 -2361
rect 19946 -2429 19997 -2395
rect 20031 -2377 20097 -2311
rect 20031 -2411 20047 -2377
rect 20081 -2411 20097 -2377
rect 20131 -2361 20165 -2345
rect 19946 -2463 19963 -2429
rect 20131 -2429 20165 -2395
rect 19997 -2463 20096 -2445
rect 19946 -2479 20096 -2463
rect 19853 -2544 19911 -2509
rect 19559 -2589 19731 -2573
rect 19559 -2623 19697 -2589
rect 19559 -2639 19731 -2623
rect 19765 -2584 19807 -2549
rect 19946 -2584 20016 -2513
rect 19765 -2589 20016 -2584
rect 19765 -2623 19960 -2589
rect 19994 -2623 20016 -2589
rect 19765 -2634 20016 -2623
rect 19559 -2719 19609 -2639
rect 19765 -2679 19807 -2634
rect 19946 -2643 20016 -2634
rect 20050 -2574 20096 -2479
rect 20050 -2583 20062 -2574
rect 20084 -2617 20096 -2608
rect 19756 -2695 19807 -2679
rect 19559 -2753 19575 -2719
rect 19559 -2769 19609 -2753
rect 19672 -2725 19706 -2702
rect 19455 -2783 19521 -2775
rect 19672 -2821 19706 -2759
rect 19790 -2729 19807 -2695
rect 19756 -2785 19807 -2729
rect 19853 -2693 19911 -2676
rect 20050 -2677 20096 -2617
rect 19853 -2727 19865 -2693
rect 19899 -2727 19911 -2693
rect 19853 -2821 19911 -2727
rect 19946 -2711 20096 -2677
rect 19946 -2719 19997 -2711
rect 19946 -2753 19963 -2719
rect 20131 -2719 20165 -2481
rect 20199 -2505 20264 -2348
rect 20298 -2353 20348 -2311
rect 20298 -2387 20314 -2353
rect 20298 -2403 20348 -2387
rect 20382 -2361 20432 -2345
rect 20382 -2395 20398 -2361
rect 20382 -2411 20432 -2395
rect 20475 -2355 20611 -2345
rect 20475 -2389 20491 -2355
rect 20525 -2389 20611 -2355
rect 20726 -2363 20792 -2311
rect 20919 -2353 20993 -2311
rect 20475 -2411 20611 -2389
rect 20382 -2437 20416 -2411
rect 20337 -2471 20416 -2437
rect 20450 -2447 20543 -2445
rect 20211 -2512 20303 -2505
rect 20211 -2552 20230 -2512
rect 20270 -2528 20303 -2512
rect 20211 -2562 20269 -2552
rect 20211 -2715 20303 -2562
rect 19946 -2769 19997 -2753
rect 20031 -2779 20047 -2745
rect 20081 -2779 20097 -2745
rect 20337 -2743 20371 -2471
rect 20450 -2473 20509 -2447
rect 20484 -2481 20509 -2473
rect 20484 -2507 20543 -2481
rect 20450 -2523 20543 -2507
rect 20405 -2583 20475 -2561
rect 20405 -2617 20417 -2583
rect 20451 -2617 20475 -2583
rect 20405 -2635 20475 -2617
rect 20405 -2669 20428 -2635
rect 20462 -2669 20475 -2635
rect 20405 -2685 20475 -2669
rect 20509 -2641 20543 -2523
rect 20577 -2567 20611 -2411
rect 20645 -2379 20679 -2363
rect 20726 -2397 20742 -2363
rect 20776 -2397 20792 -2363
rect 20826 -2379 20860 -2363
rect 20645 -2431 20679 -2413
rect 20919 -2387 20939 -2353
rect 20973 -2387 20993 -2353
rect 20919 -2403 20993 -2387
rect 21027 -2361 21061 -2345
rect 20826 -2431 20860 -2413
rect 20645 -2465 20860 -2431
rect 21027 -2437 21061 -2395
rect 21108 -2354 21282 -2345
rect 21108 -2388 21124 -2354
rect 21158 -2388 21282 -2354
rect 21108 -2413 21282 -2388
rect 21316 -2353 21366 -2311
rect 21350 -2387 21366 -2353
rect 21470 -2353 21614 -2311
rect 21316 -2403 21366 -2387
rect 21400 -2379 21434 -2363
rect 20949 -2471 21061 -2437
rect 20949 -2499 20983 -2471
rect 20683 -2533 20699 -2499
rect 20733 -2533 20983 -2499
rect 21122 -2481 21133 -2447
rect 21167 -2473 21214 -2447
rect 21122 -2505 21164 -2481
rect 20577 -2587 20915 -2567
rect 20577 -2601 20881 -2587
rect 20509 -2675 20530 -2641
rect 20564 -2675 20580 -2641
rect 20509 -2685 20580 -2675
rect 20614 -2743 20648 -2601
rect 20689 -2651 20785 -2635
rect 20723 -2685 20761 -2651
rect 20819 -2669 20847 -2635
rect 20881 -2637 20915 -2621
rect 20795 -2685 20847 -2669
rect 20949 -2671 20983 -2533
rect 20131 -2769 20165 -2753
rect 20031 -2821 20097 -2779
rect 20237 -2783 20253 -2749
rect 20287 -2783 20303 -2749
rect 20337 -2777 20386 -2743
rect 20420 -2777 20436 -2743
rect 20477 -2777 20493 -2743
rect 20527 -2777 20648 -2743
rect 20823 -2745 20889 -2729
rect 20237 -2821 20303 -2783
rect 20823 -2779 20839 -2745
rect 20873 -2779 20889 -2745
rect 20823 -2821 20889 -2779
rect 20931 -2749 20983 -2671
rect 21021 -2507 21164 -2505
rect 21198 -2507 21214 -2473
rect 21248 -2489 21282 -2413
rect 21470 -2387 21486 -2353
rect 21520 -2387 21564 -2353
rect 21598 -2387 21614 -2353
rect 21648 -2361 21729 -2345
rect 21880 -2353 21914 -2311
rect 21400 -2421 21434 -2413
rect 21682 -2395 21729 -2361
rect 21400 -2455 21560 -2421
rect 21021 -2539 21156 -2507
rect 21248 -2523 21442 -2489
rect 21476 -2523 21492 -2489
rect 21021 -2647 21063 -2539
rect 21248 -2541 21282 -2523
rect 21021 -2681 21029 -2647
rect 21021 -2697 21063 -2681
rect 21097 -2583 21167 -2573
rect 21097 -2599 21133 -2583
rect 21097 -2633 21125 -2599
rect 21159 -2633 21167 -2617
rect 21097 -2697 21167 -2633
rect 21201 -2575 21282 -2541
rect 21201 -2731 21235 -2575
rect 21349 -2588 21457 -2557
rect 21526 -2573 21560 -2455
rect 21648 -2429 21729 -2395
rect 21682 -2463 21729 -2429
rect 21648 -2497 21729 -2463
rect 21682 -2531 21729 -2497
rect 21648 -2547 21729 -2531
rect 21526 -2579 21615 -2573
rect 21383 -2597 21457 -2588
rect 21269 -2625 21313 -2609
rect 21303 -2659 21313 -2625
rect 21349 -2631 21365 -2622
rect 21399 -2631 21457 -2597
rect 21269 -2665 21313 -2659
rect 21409 -2651 21457 -2631
rect 21269 -2699 21375 -2665
rect 21045 -2745 21235 -2731
rect 20931 -2783 20951 -2749
rect 20985 -2783 21001 -2749
rect 21045 -2779 21061 -2745
rect 21095 -2779 21235 -2745
rect 21045 -2787 21235 -2779
rect 21269 -2749 21307 -2733
rect 21269 -2783 21273 -2749
rect 21341 -2745 21375 -2699
rect 21443 -2685 21457 -2651
rect 21409 -2711 21457 -2685
rect 21491 -2589 21615 -2579
rect 21491 -2623 21565 -2589
rect 21599 -2623 21615 -2589
rect 21491 -2639 21615 -2623
rect 21491 -2674 21556 -2639
rect 21663 -2673 21729 -2547
rect 21491 -2729 21555 -2674
rect 21341 -2763 21491 -2745
rect 21525 -2763 21555 -2729
rect 21341 -2779 21555 -2763
rect 21595 -2706 21629 -2684
rect 21269 -2821 21307 -2783
rect 21595 -2821 21629 -2740
rect 21663 -2707 21679 -2673
rect 21713 -2707 21729 -2673
rect 21663 -2741 21729 -2707
rect 21663 -2775 21679 -2741
rect 21713 -2775 21729 -2741
rect 21767 -2387 21783 -2353
rect 21817 -2387 21833 -2353
rect 21767 -2421 21833 -2387
rect 21767 -2455 21783 -2421
rect 21817 -2455 21833 -2421
rect 21767 -2573 21833 -2455
rect 21880 -2421 21914 -2387
rect 21880 -2489 21914 -2455
rect 21880 -2539 21914 -2523
rect 21964 -2389 22015 -2373
rect 21998 -2423 22015 -2389
rect 21964 -2428 22015 -2423
rect 21964 -2457 21974 -2428
rect 21964 -2549 21974 -2491
rect 21767 -2589 21939 -2573
rect 21767 -2623 21905 -2589
rect 21767 -2639 21939 -2623
rect 21973 -2622 21974 -2549
rect 22014 -2622 22015 -2428
rect 22061 -2382 22119 -2311
rect 22061 -2416 22073 -2382
rect 22107 -2416 22119 -2382
rect 22061 -2475 22119 -2416
rect 22061 -2509 22073 -2475
rect 22107 -2509 22119 -2475
rect 22061 -2544 22119 -2509
rect 21767 -2719 21817 -2639
rect 21973 -2679 22015 -2622
rect 21964 -2695 22015 -2679
rect 21767 -2753 21783 -2719
rect 21767 -2769 21817 -2753
rect 21880 -2725 21914 -2702
rect 21663 -2783 21729 -2775
rect 21880 -2821 21914 -2759
rect 21998 -2729 22015 -2695
rect 21964 -2785 22015 -2729
rect 22061 -2693 22119 -2676
rect 22061 -2727 22073 -2693
rect 22107 -2727 22119 -2693
rect 22061 -2821 22119 -2727
rect 14868 -2855 14897 -2821
rect 14931 -2855 14989 -2821
rect 15023 -2855 15081 -2821
rect 15115 -2855 15173 -2821
rect 15207 -2855 15265 -2821
rect 15299 -2855 15357 -2821
rect 15391 -2855 15449 -2821
rect 15483 -2855 15541 -2821
rect 15575 -2855 15633 -2821
rect 15667 -2855 15725 -2821
rect 15759 -2855 15817 -2821
rect 15851 -2855 15909 -2821
rect 15943 -2855 16001 -2821
rect 16035 -2855 16093 -2821
rect 16127 -2855 16185 -2821
rect 16219 -2855 16277 -2821
rect 16311 -2855 16369 -2821
rect 16403 -2855 16461 -2821
rect 16495 -2855 16553 -2821
rect 16587 -2855 16645 -2821
rect 16679 -2855 16737 -2821
rect 16771 -2855 16829 -2821
rect 16863 -2855 16921 -2821
rect 16955 -2855 17013 -2821
rect 17047 -2855 17105 -2821
rect 17139 -2855 17197 -2821
rect 17231 -2855 17289 -2821
rect 17323 -2855 17381 -2821
rect 17415 -2855 17473 -2821
rect 17507 -2855 17565 -2821
rect 17599 -2855 17657 -2821
rect 17691 -2855 17749 -2821
rect 17783 -2855 17841 -2821
rect 17875 -2855 17933 -2821
rect 17967 -2855 18025 -2821
rect 18059 -2855 18117 -2821
rect 18151 -2855 18209 -2821
rect 18243 -2855 18301 -2821
rect 18335 -2855 18393 -2821
rect 18427 -2855 18485 -2821
rect 18519 -2855 18577 -2821
rect 18611 -2855 18669 -2821
rect 18703 -2855 18761 -2821
rect 18795 -2855 18853 -2821
rect 18887 -2855 18945 -2821
rect 18979 -2855 19037 -2821
rect 19071 -2855 19129 -2821
rect 19163 -2855 19221 -2821
rect 19255 -2855 19313 -2821
rect 19347 -2855 19405 -2821
rect 19439 -2855 19497 -2821
rect 19531 -2855 19589 -2821
rect 19623 -2855 19681 -2821
rect 19715 -2855 19773 -2821
rect 19807 -2855 19865 -2821
rect 19899 -2855 19957 -2821
rect 19991 -2855 20049 -2821
rect 20083 -2855 20141 -2821
rect 20175 -2855 20233 -2821
rect 20267 -2855 20325 -2821
rect 20359 -2855 20417 -2821
rect 20451 -2855 20509 -2821
rect 20543 -2855 20601 -2821
rect 20635 -2855 20693 -2821
rect 20727 -2855 20785 -2821
rect 20819 -2855 20877 -2821
rect 20911 -2855 20969 -2821
rect 21003 -2855 21061 -2821
rect 21095 -2855 21153 -2821
rect 21187 -2855 21245 -2821
rect 21279 -2855 21337 -2821
rect 21371 -2855 21429 -2821
rect 21463 -2855 21521 -2821
rect 21555 -2855 21613 -2821
rect 21647 -2855 21705 -2821
rect 21739 -2855 21797 -2821
rect 21831 -2855 21889 -2821
rect 21923 -2855 21981 -2821
rect 22015 -2855 22073 -2821
rect 22107 -2855 22136 -2821
rect 13048 -3116 13668 -3026
rect 13014 -3178 13668 -3116
rect 12600 -3190 12696 -3178
rect 12440 -3212 12696 -3190
rect 12952 -3212 13668 -3178
rect 12440 -3216 13668 -3212
rect 6406 -3417 6446 -3416
rect 1905 -3423 6446 -3417
rect 1903 -3457 1963 -3423
rect 6385 -3452 6446 -3423
rect 6385 -3457 6445 -3452
rect 1903 -3483 1943 -3457
rect 1937 -5100 1943 -3483
rect 6407 -3483 6445 -3457
rect 2548 -3918 2644 -3916
rect 2552 -3950 2644 -3918
rect 3070 -3950 3162 -3916
rect 2552 -4012 2582 -3950
rect 3132 -4012 3162 -3950
rect 3258 -3950 3350 -3916
rect 3776 -3950 3870 -3916
rect 3258 -4012 3288 -3950
rect 2728 -4088 2744 -4054
rect 2812 -4088 2828 -4054
rect 2886 -4088 2902 -4054
rect 2970 -4088 2986 -4054
rect 2682 -4138 2716 -4122
rect 2682 -4730 2716 -4714
rect 2840 -4138 2874 -4122
rect 2840 -4730 2874 -4714
rect 2998 -4138 3032 -4122
rect 2998 -4730 3032 -4714
rect 2728 -4798 2744 -4764
rect 2812 -4798 2828 -4764
rect 2886 -4798 2902 -4764
rect 2970 -4798 2986 -4764
rect 2552 -4902 2582 -4840
rect 3838 -4012 3870 -3950
rect 3434 -4088 3450 -4054
rect 3518 -4088 3534 -4054
rect 3592 -4088 3608 -4054
rect 3676 -4088 3692 -4054
rect 3388 -4138 3422 -4122
rect 3388 -4730 3422 -4714
rect 3546 -4138 3580 -4122
rect 3546 -4730 3580 -4714
rect 3704 -4138 3738 -4122
rect 3704 -4730 3738 -4714
rect 3434 -4798 3450 -4764
rect 3518 -4798 3534 -4764
rect 3592 -4798 3608 -4764
rect 3676 -4798 3692 -4764
rect 3132 -4902 3162 -4840
rect 2552 -4936 2644 -4902
rect 3070 -4934 3162 -4902
rect 3258 -4902 3288 -4840
rect 3838 -4902 3870 -4840
rect 3258 -4934 3350 -4902
rect 3070 -4936 3166 -4934
rect 3254 -4936 3350 -4934
rect 3776 -4934 3870 -4902
rect 4466 -3950 4560 -3916
rect 4986 -3950 5078 -3916
rect 4466 -4012 4498 -3950
rect 5048 -4012 5078 -3950
rect 5174 -3950 5266 -3916
rect 5692 -3918 5788 -3916
rect 5692 -3950 5784 -3918
rect 5174 -4012 5204 -3950
rect 4644 -4088 4660 -4054
rect 4728 -4088 4744 -4054
rect 4802 -4088 4818 -4054
rect 4886 -4088 4902 -4054
rect 4598 -4138 4632 -4122
rect 4598 -4730 4632 -4714
rect 4756 -4138 4790 -4122
rect 4756 -4730 4790 -4714
rect 4914 -4138 4948 -4122
rect 4914 -4730 4948 -4714
rect 4644 -4798 4660 -4764
rect 4728 -4798 4744 -4764
rect 4802 -4798 4818 -4764
rect 4886 -4798 4902 -4764
rect 4466 -4902 4498 -4840
rect 5754 -4012 5784 -3950
rect 5350 -4088 5366 -4054
rect 5434 -4088 5450 -4054
rect 5508 -4088 5524 -4054
rect 5592 -4088 5608 -4054
rect 5304 -4138 5338 -4122
rect 5304 -4730 5338 -4714
rect 5462 -4138 5496 -4122
rect 5462 -4730 5496 -4714
rect 5620 -4138 5654 -4122
rect 5620 -4730 5654 -4714
rect 5350 -4798 5366 -4764
rect 5434 -4798 5450 -4764
rect 5508 -4798 5524 -4764
rect 5592 -4798 5608 -4764
rect 5048 -4902 5078 -4840
rect 4466 -4934 4560 -4902
rect 3776 -4936 3872 -4934
rect 4464 -4936 4560 -4934
rect 4986 -4934 5078 -4902
rect 5174 -4902 5204 -4840
rect 5754 -4902 5784 -4840
rect 5174 -4934 5266 -4902
rect 4986 -4936 5082 -4934
rect 5170 -4936 5266 -4934
rect 5692 -4936 5784 -4902
rect 1937 -5154 2644 -5100
rect 6407 -5104 6411 -3483
rect 1937 -6772 1990 -5154
rect 2476 -5174 2644 -5154
rect 5692 -5156 6411 -5104
rect 5692 -5174 5838 -5156
rect 2476 -5848 2586 -5174
rect 2706 -5244 2726 -5210
rect 3694 -5244 3790 -5210
rect 3756 -5306 3790 -5244
rect 2810 -5382 2826 -5348
rect 3594 -5382 3610 -5348
rect 2764 -5441 2798 -5425
rect 2764 -5633 2798 -5617
rect 3622 -5441 3656 -5425
rect 3622 -5633 3656 -5617
rect 2810 -5710 2826 -5676
rect 3594 -5710 3610 -5676
rect 3756 -5812 3790 -5752
rect 4546 -5244 4642 -5210
rect 5610 -5244 5630 -5210
rect 4546 -5306 4580 -5244
rect 4726 -5382 4742 -5348
rect 5510 -5382 5526 -5348
rect 4680 -5441 4714 -5425
rect 4680 -5633 4714 -5617
rect 5538 -5441 5572 -5425
rect 5538 -5633 5572 -5617
rect 4726 -5710 4742 -5676
rect 5510 -5710 5526 -5676
rect 4546 -5812 4580 -5752
rect 2706 -5848 2726 -5814
rect 3694 -5848 3714 -5814
rect 2476 -5910 2664 -5848
rect 2476 -6356 2630 -5910
rect 2810 -5986 2826 -5952
rect 3594 -5986 3610 -5952
rect 2764 -6045 2798 -6029
rect 2764 -6237 2798 -6221
rect 3622 -6045 3656 -6029
rect 3622 -6237 3656 -6221
rect 2810 -6314 2826 -6280
rect 3594 -6314 3610 -6280
rect 2476 -6418 2664 -6356
rect 2476 -6452 2726 -6418
rect 3694 -6452 3714 -6418
rect 2476 -6772 2644 -6452
rect 3706 -6486 3714 -6452
rect 4622 -5848 4642 -5814
rect 5610 -5848 5630 -5814
rect 5750 -5848 5838 -5174
rect 5672 -5910 5838 -5848
rect 4726 -5986 4742 -5952
rect 5510 -5986 5526 -5952
rect 4680 -6045 4714 -6029
rect 4680 -6237 4714 -6221
rect 5538 -6045 5572 -6029
rect 5538 -6237 5572 -6221
rect 4726 -6314 4742 -6280
rect 5510 -6314 5526 -6280
rect 3834 -6486 4502 -6434
rect 5706 -6356 5838 -5910
rect 5672 -6418 5838 -6356
rect 4622 -6452 4642 -6418
rect 5610 -6452 5838 -6418
rect 4622 -6486 5838 -6452
rect 3706 -6560 5838 -6486
rect 1937 -6822 2644 -6772
rect 3634 -6774 5838 -6560
rect 6324 -6774 6411 -5156
rect 1937 -8969 1943 -6822
rect 2128 -7043 3504 -6958
rect 2128 -7064 2413 -7043
rect 2130 -7077 2413 -7064
rect 3313 -7077 3504 -7043
rect 2130 -7139 2351 -7077
rect 2130 -8167 2317 -7139
rect 2496 -7126 3228 -7116
rect 2496 -7214 2510 -7126
rect 3375 -7139 3504 -7077
rect 2497 -7215 2513 -7214
rect 2581 -7215 2597 -7214
rect 2655 -7215 2671 -7214
rect 2739 -7215 2755 -7214
rect 2813 -7215 2829 -7214
rect 2897 -7215 2913 -7214
rect 2971 -7215 2987 -7214
rect 3055 -7215 3071 -7214
rect 3129 -7215 3145 -7214
rect 3213 -7215 3229 -7214
rect 2451 -7250 2485 -7249
rect 2351 -7254 2485 -7250
rect 2609 -7254 2643 -7249
rect 2767 -7254 2801 -7249
rect 2925 -7254 2959 -7249
rect 3083 -7254 3117 -7249
rect 3241 -7254 3275 -7249
rect 2351 -7265 2526 -7254
rect 2351 -7266 2451 -7265
rect 2485 -7266 2526 -7265
rect 2351 -8042 2420 -7266
rect 2512 -8042 2526 -7266
rect 2351 -8054 2526 -8042
rect 2564 -7265 2684 -7254
rect 2564 -7266 2609 -7265
rect 2643 -7266 2684 -7265
rect 2564 -8042 2578 -7266
rect 2670 -8042 2684 -7266
rect 2564 -8054 2684 -8042
rect 2722 -7265 2842 -7254
rect 2722 -7266 2767 -7265
rect 2801 -7266 2842 -7265
rect 2722 -8042 2736 -7266
rect 2828 -8042 2842 -7266
rect 2722 -8054 2842 -8042
rect 2880 -7265 3000 -7254
rect 2880 -7266 2925 -7265
rect 2959 -7266 3000 -7265
rect 2880 -8042 2894 -7266
rect 2986 -8042 3000 -7266
rect 2880 -8054 3000 -8042
rect 3036 -7265 3156 -7254
rect 3036 -7266 3083 -7265
rect 3117 -7266 3156 -7265
rect 3036 -8042 3050 -7266
rect 3142 -8042 3156 -7266
rect 3036 -8054 3156 -8042
rect 3196 -7265 3316 -7254
rect 3196 -7266 3241 -7265
rect 3275 -7266 3316 -7265
rect 3196 -8042 3210 -7266
rect 3302 -8042 3316 -7266
rect 3196 -8054 3316 -8042
rect 2351 -8057 2485 -8054
rect 2609 -8057 2643 -8054
rect 2767 -8057 2801 -8054
rect 2925 -8057 2959 -8054
rect 3083 -8057 3117 -8054
rect 3241 -8057 3275 -8054
rect 2351 -8058 2482 -8057
rect 2497 -8092 2513 -8091
rect 2581 -8092 2597 -8091
rect 2655 -8092 2671 -8091
rect 2739 -8092 2755 -8091
rect 2813 -8092 2829 -8091
rect 2897 -8092 2913 -8091
rect 2971 -8092 2987 -8091
rect 3055 -8092 3071 -8091
rect 3129 -8092 3145 -8091
rect 2130 -8229 2351 -8167
rect 2496 -8172 2512 -8092
rect 3213 -8125 3229 -8091
rect 3212 -8172 3228 -8125
rect 2496 -8184 3228 -8172
rect 3409 -8167 3504 -7139
rect 3375 -8229 3504 -8167
rect 2130 -8263 2413 -8229
rect 3313 -8263 3504 -8229
rect 2130 -8812 3504 -8263
rect 3634 -7036 6411 -6774
rect 3634 -7070 3788 -7036
rect 4688 -7070 6411 -7036
rect 3634 -7132 3726 -7070
rect 3634 -8178 3692 -7132
rect 3872 -7120 4600 -7110
rect 3872 -7208 3888 -7120
rect 4588 -7174 4600 -7120
rect 4750 -7132 6411 -7070
rect 4588 -7208 4604 -7174
rect 3826 -7254 3860 -7251
rect 3984 -7254 4018 -7251
rect 4142 -7254 4176 -7251
rect 4300 -7254 4334 -7251
rect 4458 -7254 4492 -7251
rect 4616 -7252 4650 -7251
rect 4616 -7254 4750 -7252
rect 3782 -7266 3902 -7254
rect 3782 -8044 3796 -7266
rect 3888 -8044 3902 -7266
rect 3782 -8054 3902 -8044
rect 3940 -7266 4060 -7254
rect 3940 -8044 3954 -7266
rect 4046 -8044 4060 -7266
rect 3940 -8054 4060 -8044
rect 4098 -7266 4218 -7254
rect 4098 -8044 4112 -7266
rect 4204 -8044 4218 -7266
rect 4098 -8054 4218 -8044
rect 4256 -7266 4376 -7254
rect 4256 -8044 4270 -7266
rect 4362 -8044 4376 -7266
rect 4256 -8054 4376 -8044
rect 4414 -7266 4534 -7254
rect 4414 -8044 4428 -7266
rect 4520 -8044 4534 -7266
rect 4414 -8054 4534 -8044
rect 4572 -7266 4750 -7254
rect 4572 -8044 4586 -7266
rect 4678 -8044 4750 -7266
rect 4572 -8054 4750 -8044
rect 3826 -8059 3860 -8054
rect 3984 -8059 4018 -8054
rect 4142 -8059 4176 -8054
rect 4300 -8059 4334 -8054
rect 4458 -8059 4492 -8054
rect 4616 -8060 4750 -8054
rect 3634 -8240 3726 -8178
rect 3872 -8188 3888 -8102
rect 4594 -8188 4608 -8102
rect 3872 -8196 4608 -8188
rect 4784 -8178 6411 -7132
rect 4750 -8240 6411 -8178
rect 3634 -8274 3788 -8240
rect 4688 -8274 6411 -8240
rect 2130 -8814 3468 -8812
rect 1903 -8988 1943 -8969
rect 3634 -8969 6411 -8274
rect 12440 -3630 12462 -3216
rect 12588 -3416 13668 -3216
rect 13646 -3630 13668 -3416
rect 13936 -3116 14760 -3016
rect 14996 -3026 15092 -2992
rect 16020 -3004 16222 -2992
rect 16020 -3026 16120 -3004
rect 14996 -3088 15030 -3026
rect 13936 -3128 14136 -3116
rect 13936 -3460 13950 -3128
rect 14122 -3460 14136 -3128
rect 16082 -3088 16120 -3026
rect 15156 -3128 15172 -3094
rect 15940 -3128 15956 -3094
rect 15110 -3178 15144 -3162
rect 15110 -3270 15144 -3254
rect 15968 -3178 16002 -3162
rect 15968 -3270 16002 -3254
rect 15156 -3338 15172 -3304
rect 15940 -3338 15956 -3304
rect 14996 -3406 15030 -3344
rect 16116 -3344 16120 -3088
rect 16082 -3406 16120 -3344
rect 14996 -3440 15092 -3406
rect 16020 -3440 16120 -3406
rect 13936 -3476 14136 -3460
rect 15008 -3442 16120 -3440
rect 16212 -3438 16222 -3004
rect 15008 -3516 15034 -3442
rect 16212 -3516 16220 -3438
rect 15008 -3534 16220 -3516
rect 12440 -3646 13668 -3630
rect 1902 -8989 1944 -8988
rect 3634 -8989 6445 -8969
rect 1902 -8995 6445 -8989
rect 1902 -9029 1963 -8995
rect 6385 -9029 6445 -8995
rect 8757 -4231 8817 -4197
rect 25211 -4231 25271 -4197
rect 8757 -4257 8791 -4231
rect 1902 -9030 1944 -9029
rect 25237 -4257 25271 -4231
rect 8880 -4316 25158 -4298
rect 8791 -5608 8792 -5450
rect 8880 -5476 8900 -4316
rect 11694 -4734 12058 -4548
rect 10462 -4748 12058 -4734
rect 16094 -4556 16958 -4548
rect 17330 -4556 18192 -4548
rect 16094 -4564 18192 -4556
rect 16094 -4598 16196 -4564
rect 18098 -4598 18192 -4564
rect 16094 -4660 16134 -4598
rect 10462 -4782 10574 -4748
rect 15188 -4782 15282 -4750
rect 10462 -4844 10512 -4782
rect 10462 -4970 10478 -4844
rect 11436 -4886 12014 -4818
rect 12592 -4886 12844 -4816
rect 13748 -4886 14326 -4818
rect 15250 -4844 15282 -4782
rect 10658 -4920 10674 -4886
rect 11042 -4920 11058 -4886
rect 11236 -4920 11252 -4886
rect 11620 -4920 11830 -4886
rect 12198 -4920 12214 -4886
rect 12392 -4920 12408 -4886
rect 12776 -4920 12844 -4886
rect 12970 -4920 12986 -4886
rect 13354 -4920 13370 -4886
rect 13548 -4920 13564 -4886
rect 13932 -4920 14142 -4886
rect 14510 -4920 14526 -4886
rect 14704 -4920 14720 -4886
rect 15088 -4920 15104 -4886
rect 10612 -4958 10646 -4954
rect 11070 -4958 11104 -4954
rect 11190 -4958 11224 -4954
rect 11436 -4958 12014 -4920
rect 12226 -4958 12260 -4954
rect 12346 -4958 12380 -4954
rect 12592 -4958 12844 -4920
rect 12924 -4958 12958 -4954
rect 13382 -4958 13416 -4954
rect 13502 -4958 13536 -4954
rect 13748 -4958 14326 -4920
rect 14538 -4958 14572 -4954
rect 14658 -4958 14692 -4954
rect 15116 -4958 15150 -4954
rect 10512 -4970 11230 -4958
rect 11224 -5346 11230 -4970
rect 10462 -5472 10478 -5346
rect 10512 -5358 11230 -5346
rect 11436 -5354 11452 -4958
rect 11992 -5354 12014 -4958
rect 10612 -5362 10646 -5358
rect 11070 -5362 11104 -5358
rect 11190 -5362 11224 -5358
rect 11436 -5396 12014 -5354
rect 12104 -4970 12504 -4958
rect 12104 -5346 12122 -4970
rect 12488 -5346 12504 -4970
rect 12104 -5358 12504 -5346
rect 12592 -5358 12604 -4958
rect 12826 -4970 12844 -4958
rect 12838 -5346 12844 -4970
rect 12826 -5358 12844 -5346
rect 12918 -4970 13178 -4958
rect 12918 -5346 12924 -4970
rect 13168 -5346 13178 -4970
rect 12918 -5358 13178 -5346
rect 13260 -4970 13660 -4958
rect 13260 -5346 13276 -4970
rect 13642 -5346 13660 -4970
rect 13260 -5358 13660 -5346
rect 13748 -5354 13768 -4958
rect 14308 -5354 14326 -4958
rect 12226 -5362 12260 -5358
rect 12346 -5362 12380 -5358
rect 12592 -5396 12844 -5358
rect 12924 -5362 12958 -5358
rect 13382 -5362 13416 -5358
rect 13502 -5362 13536 -5358
rect 13748 -5396 14326 -5354
rect 14532 -4970 15250 -4958
rect 14532 -5346 14538 -4970
rect 14532 -5358 15250 -5346
rect 14538 -5362 14572 -5358
rect 14658 -5362 14692 -5358
rect 15116 -5362 15150 -5358
rect 10658 -5430 10674 -5396
rect 11042 -5430 11058 -5396
rect 11236 -5430 11252 -5396
rect 11620 -5430 11830 -5396
rect 12198 -5430 12214 -5396
rect 12392 -5430 12408 -5396
rect 12776 -5430 12844 -5396
rect 12970 -5430 12986 -5396
rect 13354 -5430 13370 -5396
rect 13548 -5430 13564 -5396
rect 13932 -5430 14142 -5396
rect 14510 -5430 14526 -5396
rect 14704 -5430 14720 -5396
rect 15088 -5430 15104 -5396
rect 10462 -5476 10512 -5472
rect 8880 -5494 10512 -5476
rect 10478 -5534 10512 -5494
rect 11436 -5500 12014 -5430
rect 12592 -5500 12844 -5430
rect 13748 -5500 14326 -5430
rect 15250 -5530 15282 -5472
rect 16094 -5530 16100 -4660
rect 15250 -5534 16100 -5530
rect 10478 -5568 10574 -5534
rect 15188 -5548 16100 -5534
rect 15188 -5568 15284 -5548
rect 8791 -5636 16060 -5608
rect 8791 -5640 15260 -5636
rect 8791 -7366 8878 -5640
rect 15938 -5752 16060 -5636
rect 16260 -4666 18034 -4640
rect 16260 -4700 16276 -4666
rect 16644 -4700 16734 -4666
rect 17102 -4700 17192 -4666
rect 17560 -4700 17650 -4666
rect 18018 -4700 18034 -4666
rect 18160 -4660 18192 -4598
rect 16648 -4734 16924 -4700
rect 16210 -4744 16924 -4734
rect 16210 -4750 16666 -4744
rect 16210 -5526 16214 -4750
rect 16248 -4794 16666 -4750
rect 16248 -5526 16666 -5484
rect 16210 -5530 16666 -5526
rect 16878 -5530 16924 -4744
rect 16210 -5542 16924 -5530
rect 17026 -4750 17266 -4734
rect 17026 -5526 17044 -4750
rect 17246 -5526 17266 -4750
rect 17026 -5542 17266 -5526
rect 17498 -4750 18082 -4734
rect 17498 -5526 17514 -4750
rect 18080 -5526 18082 -4750
rect 17498 -5542 18082 -5526
rect 16648 -5576 16924 -5542
rect 16100 -5678 16134 -5616
rect 16260 -5610 16276 -5576
rect 16644 -5610 16734 -5576
rect 17102 -5610 17192 -5576
rect 17560 -5610 17650 -5576
rect 18018 -5610 18034 -5576
rect 16260 -5636 18034 -5610
rect 21246 -5232 22086 -5218
rect 21246 -5266 21348 -5232
rect 21934 -5266 22086 -5232
rect 21246 -5328 21286 -5266
rect 18848 -5360 20732 -5352
rect 18848 -5394 18884 -5360
rect 20612 -5394 20732 -5360
rect 18160 -5674 18192 -5616
rect 18848 -5530 18878 -5394
rect 20674 -5456 20732 -5394
rect 18948 -5496 18964 -5462
rect 20532 -5496 20548 -5462
rect 18848 -5546 18936 -5530
rect 18848 -5548 18902 -5546
rect 18160 -5678 18788 -5674
rect 16100 -5712 16196 -5678
rect 18098 -5694 18788 -5678
rect 18098 -5712 18194 -5694
rect 18862 -5622 18902 -5548
rect 18862 -5638 18936 -5622
rect 20560 -5546 20594 -5530
rect 20560 -5638 20594 -5622
rect 15938 -5758 18742 -5752
rect 16602 -5762 18742 -5758
rect 10492 -5806 15260 -5776
rect 10492 -5840 10618 -5806
rect 15150 -5840 15260 -5806
rect 10492 -5902 10556 -5840
rect 10492 -6000 10522 -5902
rect 10682 -5908 15086 -5888
rect 10682 -5942 10698 -5908
rect 11066 -5942 11270 -5908
rect 11638 -5942 11842 -5908
rect 12210 -5942 12414 -5908
rect 12782 -5942 12986 -5908
rect 13354 -5942 13558 -5908
rect 13926 -5942 14130 -5908
rect 14498 -5942 14702 -5908
rect 15070 -5942 15086 -5908
rect 10682 -5948 15086 -5942
rect 15212 -5902 15260 -5840
rect 16602 -5878 16776 -5762
rect 17510 -5878 17700 -5762
rect 18728 -5850 18742 -5762
rect 18788 -5790 18808 -5712
rect 18862 -5774 18904 -5638
rect 18948 -5706 18964 -5672
rect 20532 -5706 20548 -5672
rect 20708 -5712 20732 -5456
rect 21246 -5486 21252 -5328
rect 20674 -5774 20732 -5712
rect 18862 -5790 18884 -5774
rect 18788 -5808 18884 -5790
rect 20612 -5776 20732 -5774
rect 21214 -5776 21252 -5486
rect 20612 -5790 21252 -5776
rect 20612 -5808 20708 -5790
rect 21996 -5328 22086 -5266
rect 21412 -5368 21428 -5334
rect 21596 -5368 21612 -5334
rect 21670 -5368 21686 -5334
rect 21854 -5368 21870 -5334
rect 21286 -5418 21400 -5402
rect 21286 -5494 21366 -5418
rect 21286 -5508 21400 -5494
rect 21366 -5510 21400 -5508
rect 21624 -5418 21658 -5402
rect 21624 -5510 21658 -5494
rect 21882 -5418 21916 -5402
rect 21882 -5510 21916 -5494
rect 21412 -5578 21428 -5544
rect 21596 -5578 21612 -5544
rect 21670 -5578 21686 -5544
rect 21854 -5578 21870 -5544
rect 21366 -5628 21400 -5612
rect 21366 -5720 21400 -5704
rect 21624 -5628 21658 -5612
rect 21624 -5720 21658 -5704
rect 21882 -5628 21916 -5612
rect 21882 -5720 21916 -5704
rect 21412 -5788 21428 -5754
rect 21596 -5788 21612 -5754
rect 21670 -5788 21686 -5754
rect 21854 -5788 21870 -5754
rect 18728 -5864 21204 -5850
rect 20504 -5870 21204 -5864
rect 10636 -5988 10670 -5985
rect 11088 -5988 11248 -5984
rect 10556 -6000 11248 -5988
rect 11242 -6378 11248 -6000
rect 10492 -6528 10522 -6378
rect 10556 -6388 11248 -6378
rect 10636 -6393 10670 -6388
rect 11088 -6394 11248 -6388
rect 11362 -6430 11542 -5948
rect 11588 -6000 11892 -5984
rect 11588 -6378 11602 -6000
rect 11878 -6378 11892 -6000
rect 11588 -6394 11892 -6378
rect 11936 -6430 12116 -5948
rect 12912 -5982 13260 -5948
rect 12164 -6000 12850 -5984
rect 12164 -6378 12176 -6000
rect 12452 -6001 12850 -6000
rect 12452 -6377 12810 -6001
rect 12844 -6377 12850 -6001
rect 12452 -6378 12850 -6377
rect 12164 -6394 12850 -6378
rect 12912 -6392 12924 -5982
rect 13252 -6392 13260 -5982
rect 12912 -6430 13260 -6392
rect 13300 -6000 13604 -5984
rect 13300 -6378 13316 -6000
rect 13592 -6378 13604 -6000
rect 13300 -6394 13604 -6378
rect 13650 -6430 13830 -5948
rect 13874 -6000 14178 -5984
rect 13874 -6378 13886 -6000
rect 14162 -6378 14178 -6000
rect 13874 -6394 14178 -6378
rect 14222 -6430 14402 -5948
rect 14520 -5988 14680 -5984
rect 15098 -5988 15132 -5985
rect 14520 -6000 15212 -5988
rect 15246 -6000 15260 -5902
rect 15938 -5912 16176 -5888
rect 18118 -5912 18330 -5886
rect 15938 -5974 16114 -5912
rect 14520 -6378 14526 -6000
rect 14520 -6388 15212 -6378
rect 14520 -6394 14680 -6388
rect 15098 -6393 15132 -6388
rect 10682 -6436 15086 -6430
rect 10682 -6470 10698 -6436
rect 11066 -6470 11270 -6436
rect 11638 -6470 11842 -6436
rect 12210 -6470 12414 -6436
rect 12782 -6470 12986 -6436
rect 13354 -6470 13558 -6436
rect 13926 -6470 14130 -6436
rect 14498 -6470 14702 -6436
rect 15070 -6470 15086 -6436
rect 10682 -6476 15086 -6470
rect 10636 -6518 10670 -6513
rect 11088 -6518 11248 -6512
rect 10556 -6528 11248 -6518
rect 11242 -6906 11248 -6528
rect 10492 -7004 10522 -6906
rect 10556 -6918 11248 -6906
rect 10636 -6921 10670 -6918
rect 11088 -6922 11248 -6918
rect 11362 -6958 11542 -6476
rect 11586 -6528 11890 -6512
rect 11586 -6906 11602 -6528
rect 11878 -6906 11890 -6528
rect 11586 -6922 11890 -6906
rect 11936 -6958 12116 -6476
rect 12160 -6528 12464 -6512
rect 12160 -6530 12238 -6528
rect 12160 -6908 12174 -6530
rect 12388 -6530 12464 -6528
rect 12450 -6908 12464 -6530
rect 12160 -6922 12464 -6908
rect 12508 -6958 12688 -6476
rect 12730 -6528 13034 -6512
rect 12730 -6906 12742 -6528
rect 13018 -6906 13034 -6528
rect 12730 -6922 13034 -6906
rect 13080 -6958 13260 -6476
rect 13304 -6528 13608 -6512
rect 13304 -6906 13316 -6528
rect 13592 -6906 13608 -6528
rect 13304 -6922 13608 -6906
rect 13650 -6958 13830 -6476
rect 13876 -6528 14180 -6512
rect 13876 -6906 13888 -6528
rect 14164 -6906 14180 -6528
rect 13876 -6922 14180 -6906
rect 14222 -6958 14402 -6476
rect 14522 -6518 14682 -6512
rect 15098 -6518 15132 -6513
rect 14522 -6528 15212 -6518
rect 15246 -6528 15260 -6378
rect 14522 -6906 14526 -6528
rect 14522 -6918 15212 -6906
rect 14522 -6922 14682 -6918
rect 15098 -6921 15132 -6918
rect 10492 -7066 10556 -7004
rect 10682 -6964 15086 -6958
rect 10682 -6998 10698 -6964
rect 11066 -6998 11270 -6964
rect 11638 -6998 11842 -6964
rect 12210 -6998 12414 -6964
rect 12782 -6998 12986 -6964
rect 13354 -6998 13558 -6964
rect 13926 -6998 14130 -6964
rect 14498 -6998 14702 -6964
rect 15070 -6998 15086 -6964
rect 10682 -7018 15086 -6998
rect 15246 -7004 15260 -6906
rect 15212 -7066 15260 -7004
rect 10492 -7100 10618 -7066
rect 15150 -7100 15260 -7066
rect 10492 -7114 15260 -7100
rect 15938 -7020 16080 -5974
rect 16156 -5956 17118 -5950
rect 16156 -5960 16770 -5956
rect 16156 -6050 16162 -5960
rect 16608 -6016 16770 -5960
rect 17066 -6016 17118 -5956
rect 16644 -6050 16734 -6016
rect 17102 -6050 17118 -6016
rect 17176 -5956 18138 -5950
rect 17176 -6016 17228 -5956
rect 17524 -5960 18138 -5956
rect 17524 -6016 17686 -5960
rect 17176 -6050 17192 -6016
rect 17560 -6050 17650 -6016
rect 18132 -6050 18138 -5960
rect 18180 -5974 18330 -5912
rect 16208 -6108 16770 -6092
rect 16208 -6109 16224 -6108
rect 16208 -6885 16214 -6109
rect 16208 -6886 16224 -6885
rect 16758 -6886 16770 -6108
rect 16208 -6902 16770 -6886
rect 16998 -6106 17298 -6092
rect 16998 -6890 17014 -6106
rect 17280 -6890 17298 -6106
rect 16998 -6902 17298 -6890
rect 17520 -6108 18082 -6092
rect 17520 -6886 17532 -6108
rect 18066 -6109 18082 -6108
rect 18080 -6885 18082 -6109
rect 18066 -6886 18082 -6885
rect 17520 -6902 18082 -6886
rect 15938 -7082 16114 -7020
rect 16156 -7034 16162 -6944
rect 17102 -6978 17118 -6944
rect 17078 -7034 17118 -6978
rect 16156 -7044 17118 -7034
rect 17176 -6978 17192 -6944
rect 17176 -7034 17216 -6978
rect 18132 -7034 18138 -6944
rect 17176 -7044 18138 -7034
rect 18214 -7020 18330 -5974
rect 20504 -6354 20736 -5870
rect 18834 -6364 20736 -6354
rect 18834 -6398 18864 -6364
rect 20592 -6398 20736 -6364
rect 18834 -6543 18892 -6398
rect 20654 -6460 20736 -6398
rect 18928 -6500 18944 -6466
rect 20512 -6500 20528 -6466
rect 18834 -6559 18916 -6543
rect 18834 -6635 18882 -6559
rect 18834 -6651 18916 -6635
rect 20540 -6559 20574 -6543
rect 20540 -6651 20574 -6635
rect 18834 -6796 18892 -6651
rect 18928 -6728 18944 -6694
rect 20512 -6728 20528 -6694
rect 20688 -6734 20736 -6460
rect 21184 -5924 21204 -5870
rect 21252 -5856 21286 -5794
rect 22030 -5794 22086 -5328
rect 23274 -5322 23356 -5298
rect 23662 -5322 23778 -5298
rect 23274 -5384 23294 -5322
rect 23376 -5402 23642 -5322
rect 23376 -5404 23446 -5402
rect 22816 -5712 23260 -5406
rect 23430 -5436 23446 -5404
rect 23572 -5404 23642 -5402
rect 23724 -5384 23778 -5322
rect 23572 -5436 23588 -5404
rect 23362 -5464 23396 -5448
rect 23362 -5648 23396 -5632
rect 23622 -5464 23656 -5448
rect 23622 -5648 23656 -5632
rect 23430 -5694 23446 -5660
rect 23572 -5694 23588 -5660
rect 22816 -5758 23294 -5712
rect 21996 -5852 22086 -5794
rect 22638 -5774 23294 -5758
rect 23758 -5712 23778 -5384
rect 23724 -5774 23778 -5712
rect 22638 -5808 23356 -5774
rect 23662 -5808 23778 -5774
rect 22638 -5834 23778 -5808
rect 25134 -5834 25158 -4316
rect 22638 -5852 25158 -5834
rect 21996 -5856 25158 -5852
rect 21252 -5890 21348 -5856
rect 21934 -5872 25158 -5856
rect 21934 -5890 22030 -5872
rect 23754 -5874 25158 -5872
rect 21184 -5946 25237 -5924
rect 21184 -5948 24312 -5946
rect 21184 -6224 22398 -5948
rect 21184 -6228 22118 -6224
rect 21184 -6262 21348 -6228
rect 21934 -6262 22118 -6228
rect 21184 -6324 21286 -6262
rect 21184 -6580 21252 -6324
rect 20654 -6796 20736 -6734
rect 18834 -6830 18864 -6796
rect 20592 -6830 20736 -6796
rect 18834 -6844 20736 -6830
rect 21202 -6826 21252 -6580
rect 21996 -6324 22118 -6262
rect 21412 -6364 21428 -6330
rect 21596 -6364 21612 -6330
rect 21670 -6364 21686 -6330
rect 21854 -6364 21870 -6330
rect 21366 -6423 21400 -6407
rect 21366 -6515 21400 -6499
rect 21624 -6423 21658 -6407
rect 21624 -6515 21658 -6499
rect 21882 -6423 21916 -6407
rect 21882 -6515 21916 -6499
rect 21412 -6592 21428 -6558
rect 21596 -6592 21612 -6558
rect 21670 -6592 21686 -6558
rect 21854 -6592 21870 -6558
rect 21366 -6636 21400 -6635
rect 21286 -6651 21400 -6636
rect 21286 -6727 21366 -6651
rect 21286 -6742 21400 -6727
rect 21366 -6743 21400 -6742
rect 21624 -6651 21658 -6635
rect 21624 -6743 21658 -6727
rect 21882 -6651 21916 -6635
rect 21882 -6743 21916 -6727
rect 21412 -6820 21428 -6786
rect 21596 -6820 21612 -6786
rect 21670 -6820 21686 -6786
rect 21854 -6820 21870 -6786
rect 21202 -6888 21286 -6826
rect 22030 -6826 22118 -6324
rect 22620 -6246 24312 -5948
rect 22620 -6290 24114 -6246
rect 22620 -6324 23044 -6290
rect 24018 -6324 24114 -6290
rect 22620 -6386 22982 -6324
rect 22620 -6694 22948 -6386
rect 22930 -6714 22948 -6694
rect 24080 -6386 24114 -6324
rect 23127 -6438 23143 -6404
rect 23919 -6438 23935 -6404
rect 23050 -6466 23084 -6450
rect 23050 -6650 23084 -6634
rect 23978 -6466 24012 -6450
rect 23978 -6650 24012 -6634
rect 23127 -6696 23143 -6662
rect 23919 -6696 23935 -6662
rect 22930 -6776 22982 -6714
rect 23332 -6774 23730 -6696
rect 24080 -6774 24114 -6714
rect 23332 -6776 24114 -6774
rect 22930 -6802 23044 -6776
rect 24018 -6802 24114 -6776
rect 25178 -6802 25237 -5946
rect 21996 -6888 22118 -6826
rect 21202 -6922 21348 -6888
rect 21934 -6922 22118 -6888
rect 21202 -6930 22118 -6922
rect 18180 -7082 18330 -7020
rect 15938 -7114 16176 -7082
rect 18118 -7114 18330 -7082
rect 25180 -7248 25237 -6802
rect 21202 -7250 25237 -7248
rect 10008 -7270 25237 -7250
rect 10008 -7320 10078 -7270
rect 10008 -7366 10080 -7320
rect 8791 -7416 10080 -7366
rect 10490 -7342 10586 -7308
rect 24686 -7342 24782 -7308
rect 10490 -7380 10524 -7342
rect 8791 -7454 9614 -7416
rect 8920 -7608 9130 -7586
rect 8920 -10142 8940 -7608
rect 9046 -7620 9130 -7608
rect 9386 -7620 9482 -7586
rect 9046 -7682 9068 -7620
rect 9448 -7682 9482 -7620
rect 9150 -7700 9366 -7684
rect 9150 -7734 9220 -7700
rect 9296 -7734 9366 -7700
rect 9150 -7746 9366 -7734
rect 9136 -7762 9380 -7746
rect 9170 -7774 9346 -7762
rect 9170 -9240 9208 -7774
rect 9304 -9240 9346 -7774
rect 9170 -9268 9346 -9240
rect 9136 -9346 9170 -9330
rect 9346 -9346 9380 -9330
rect 9046 -9422 9068 -9410
rect 9204 -9392 9220 -9358
rect 9296 -9392 9312 -9358
rect 9204 -9422 9312 -9392
rect 9648 -7434 10046 -7416
rect 9648 -7438 9809 -7434
rect 9792 -7454 9809 -7438
rect 9793 -7468 9809 -7454
rect 9885 -7438 10046 -7434
rect 9885 -7454 9902 -7438
rect 9885 -7468 9901 -7454
rect 9716 -7496 9750 -7480
rect 9944 -7496 9978 -7480
rect 9750 -7570 9944 -7552
rect 9750 -9050 9788 -7570
rect 9904 -9050 9944 -7570
rect 9750 -9064 9944 -9050
rect 9716 -9080 9978 -9064
rect 9736 -9092 9952 -9080
rect 9736 -9126 9809 -9092
rect 9885 -9126 9952 -9092
rect 9736 -9136 9952 -9126
rect 9614 -9206 9648 -9144
rect 10046 -9206 10080 -9144
rect 9614 -9240 9710 -9206
rect 9984 -9240 10080 -9206
rect 10146 -7404 10524 -7380
rect 10146 -9088 10490 -7404
rect 10146 -9386 10162 -9088
rect 9482 -9408 10162 -9386
rect 9448 -9422 9466 -9410
rect 9046 -9442 9466 -9422
rect 10362 -9866 10490 -9088
rect 24748 -7368 24782 -7342
rect 24748 -7404 25152 -7368
rect 10618 -7508 10620 -7438
rect 10618 -7604 11048 -7508
rect 10618 -7674 10620 -7604
rect 24220 -7770 24650 -7674
rect 10620 -7936 11050 -7840
rect 24220 -8102 24650 -8006
rect 10620 -8268 11050 -8172
rect 24220 -8268 24650 -8266
rect 24220 -8434 24650 -8338
rect 10620 -8600 11050 -8504
rect 24220 -8600 24650 -8598
rect 24220 -8766 24650 -8670
rect 10620 -8932 11050 -8836
rect 24220 -8932 24650 -8930
rect 24220 -9098 24650 -9002
rect 10620 -9264 11050 -9168
rect 10620 -9430 11050 -9428
rect 24220 -9430 24650 -9334
rect 10620 -9596 11050 -9500
rect 24220 -9762 24650 -9666
rect 10362 -9928 10524 -9866
rect 24782 -9866 24788 -7404
rect 24748 -9928 24788 -9866
rect 10362 -9960 10586 -9928
rect 24686 -9960 24788 -9928
rect 25116 -10142 25152 -7404
rect 8920 -10176 25152 -10142
rect 8757 -10301 8791 -10275
rect 25237 -10301 25271 -10275
rect 8757 -10335 8817 -10301
rect 25211 -10335 25271 -10301
rect 1683 -11629 1743 -11595
rect 25453 -11629 25513 -11595
rect 1683 -11655 1717 -11629
rect 22120 -11655 25513 -11629
rect 22120 -11668 25479 -11655
rect 1844 -11798 21916 -11756
rect 1844 -11824 7814 -11798
rect 1844 -13814 1996 -11824
rect 7070 -12034 7814 -11824
rect 7070 -12040 13436 -12034
rect 7070 -12074 7242 -12040
rect 7610 -12074 13436 -12040
rect 7070 -12136 7180 -12074
rect 7070 -12564 7146 -12136
rect 7672 -12100 13436 -12074
rect 7672 -12134 8184 -12100
rect 13268 -12134 13436 -12100
rect 7672 -12136 8232 -12134
rect 7326 -12212 7342 -12178
rect 7510 -12212 7526 -12178
rect 7180 -12262 7314 -12246
rect 7180 -12438 7280 -12262
rect 7180 -12454 7314 -12438
rect 7538 -12262 7572 -12246
rect 7538 -12454 7572 -12438
rect 7326 -12522 7342 -12488
rect 7510 -12522 7526 -12488
rect 7070 -12626 7180 -12564
rect 7706 -12196 8232 -12136
rect 7706 -12508 8088 -12196
rect 8122 -12304 8232 -12196
rect 13330 -12194 13436 -12134
rect 13330 -12196 20656 -12194
rect 8268 -12272 8284 -12238
rect 9852 -12264 9868 -12238
rect 9852 -12272 9886 -12264
rect 9926 -12272 9942 -12238
rect 11510 -12272 11526 -12238
rect 11584 -12272 11600 -12238
rect 13168 -12272 13184 -12238
rect 8122 -12322 8256 -12304
rect 8122 -12382 8222 -12322
rect 8122 -12400 8256 -12382
rect 8336 -12306 9886 -12272
rect 8336 -12322 9914 -12306
rect 8336 -12382 8348 -12322
rect 9840 -12382 9880 -12322
rect 8336 -12398 9914 -12382
rect 11538 -12322 11572 -12306
rect 11538 -12398 11572 -12382
rect 13196 -12322 13230 -12306
rect 13196 -12398 13230 -12382
rect 8122 -12508 8232 -12400
rect 8336 -12432 9886 -12398
rect 8268 -12466 8284 -12432
rect 9852 -12442 9886 -12432
rect 9852 -12466 9868 -12442
rect 9926 -12466 9942 -12432
rect 11510 -12466 11526 -12432
rect 11584 -12466 11600 -12432
rect 13168 -12466 13184 -12432
rect 7706 -12564 8232 -12508
rect 7672 -12570 8232 -12564
rect 13364 -12508 20656 -12196
rect 13330 -12510 20656 -12508
rect 13330 -12570 13436 -12510
rect 20150 -12566 20656 -12510
rect 21870 -12566 21916 -11798
rect 22120 -12538 22152 -11668
rect 25426 -11672 25479 -11668
rect 7672 -12604 8184 -12570
rect 13268 -12604 13436 -12570
rect 7672 -12626 13436 -12604
rect 7070 -12660 7242 -12626
rect 7610 -12660 13436 -12626
rect 7070 -12680 13436 -12660
rect 20150 -12646 20656 -12600
rect 21870 -12646 21918 -12566
rect 20150 -12662 21918 -12646
rect 7070 -12792 7778 -12680
rect 20150 -12700 21884 -12662
rect 20786 -12734 20920 -12700
rect 21696 -12734 21884 -12700
rect 20150 -12752 21884 -12734
rect 7070 -12862 7778 -12826
rect 2982 -12888 7778 -12862
rect 2982 -13524 3004 -12888
rect 3038 -12898 7778 -12888
rect 3038 -12922 19062 -12898
rect 3038 -12988 3134 -12922
rect 3566 -12988 18534 -12922
rect 18502 -12992 18534 -12988
rect 18966 -12992 19062 -12922
rect 18502 -13088 19062 -12992
rect 18502 -13154 18534 -13088
rect 18966 -13154 19062 -13088
rect 19822 -12762 21884 -12752
rect 3134 -13254 3566 -13158
rect 3038 -13490 3134 -13422
rect 3566 -13490 18534 -13422
rect 18966 -13490 19062 -13422
rect 3038 -13524 19062 -13490
rect 19096 -13524 19788 -13098
rect 2982 -13538 19788 -13524
rect 19328 -13730 19788 -13538
rect 19398 -13764 19788 -13730
rect 19328 -13814 19788 -13764
rect 1844 -13826 19788 -13814
rect 1844 -18114 2002 -13826
rect 2036 -13860 19460 -13826
rect 2036 -13926 2132 -13860
rect 2564 -13926 18932 -13860
rect 19364 -13926 19460 -13860
rect 2132 -14192 2564 -14096
rect 18932 -14358 19364 -14262
rect 2564 -14428 2566 -14368
rect 2134 -14524 2566 -14428
rect 2564 -14584 2566 -14524
rect 18932 -14690 19364 -14594
rect 2132 -14856 2564 -14760
rect 18932 -15022 19364 -14926
rect 2132 -15188 2564 -15092
rect 18932 -15354 19364 -15258
rect 2130 -15424 2132 -15362
rect 2130 -15520 2562 -15424
rect 2130 -15578 2132 -15520
rect 18932 -15686 19364 -15590
rect 2132 -15852 2564 -15756
rect 18932 -16018 19364 -15922
rect 2132 -16184 2564 -16088
rect 18932 -16350 19364 -16254
rect 2132 -16516 2564 -16420
rect 18932 -16682 19364 -16586
rect 2130 -16752 2132 -16692
rect 2130 -16848 2562 -16752
rect 2130 -16908 2132 -16848
rect 18932 -17014 19364 -16918
rect 2130 -17084 2132 -17024
rect 2130 -17180 2562 -17084
rect 2130 -17240 2132 -17180
rect 18932 -17346 19364 -17250
rect 2132 -17512 2564 -17416
rect 18932 -17678 19364 -17582
rect 2132 -17844 2564 -17748
rect 2036 -18080 2132 -18014
rect 2564 -18080 18932 -18014
rect 19364 -18080 19460 -18014
rect 2036 -18114 19460 -18080
rect 19494 -15542 19788 -13826
rect 19822 -13130 19926 -12762
rect 19960 -13130 20836 -12762
rect 20870 -13130 21746 -12762
rect 21780 -13130 21884 -12762
rect 19822 -13158 21884 -13130
rect 19822 -13190 20010 -13158
rect 19822 -15014 19874 -13190
rect 19994 -13192 20010 -13190
rect 20786 -13190 20920 -13158
rect 20786 -13192 20802 -13190
rect 20904 -13192 20920 -13190
rect 21696 -13190 21884 -13158
rect 21696 -13192 21712 -13190
rect 19994 -13242 21712 -13228
rect 19994 -13244 20918 -13242
rect 19926 -13340 19960 -13324
rect 19994 -13352 20008 -13244
rect 20788 -13286 20918 -13244
rect 20788 -13352 20802 -13286
rect 19994 -13368 20802 -13352
rect 20836 -13340 20870 -13324
rect 19924 -13626 19926 -13426
rect 20904 -13350 20918 -13286
rect 21698 -13350 21712 -13242
rect 20904 -13368 21712 -13350
rect 21746 -13340 21780 -13324
rect 19960 -13452 20836 -13426
rect 19960 -13600 19998 -13452
rect 20798 -13600 20836 -13452
rect 19960 -13626 20836 -13600
rect 20870 -13452 21746 -13426
rect 20870 -13600 20908 -13452
rect 21708 -13600 21746 -13452
rect 20870 -13626 21746 -13600
rect 19926 -13724 19960 -13708
rect 19994 -13702 20802 -13680
rect 19994 -13890 20010 -13702
rect 20786 -13760 20802 -13702
rect 20836 -13724 20870 -13708
rect 20904 -13700 21712 -13680
rect 20904 -13760 20920 -13700
rect 20786 -13800 20920 -13760
rect 21696 -13800 21712 -13700
rect 21746 -13724 21780 -13708
rect 20786 -13820 21712 -13800
rect 21816 -13758 21884 -13190
rect 22120 -12574 24616 -12538
rect 22120 -12608 22478 -12574
rect 24452 -12608 24616 -12574
rect 22120 -12670 24616 -12608
rect 21918 -13758 21956 -13746
rect 20786 -13890 20802 -13820
rect 19994 -13896 20204 -13890
rect 19926 -13918 19960 -13902
rect 19926 -14302 19960 -14286
rect 20174 -14308 20204 -13896
rect 19994 -14314 20204 -14308
rect 20622 -13896 20802 -13890
rect 20622 -14308 20654 -13896
rect 20836 -13918 20870 -13902
rect 20904 -13952 20920 -13856
rect 21696 -13952 21712 -13856
rect 21816 -13874 21828 -13758
rect 21944 -13874 21956 -13758
rect 20904 -13966 21712 -13952
rect 21746 -13918 21780 -13902
rect 20870 -14052 21746 -14008
rect 20870 -14286 20916 -14052
rect 20836 -14302 20916 -14286
rect 20854 -14308 20916 -14302
rect 21698 -14286 21746 -14052
rect 21698 -14302 21780 -14286
rect 21698 -14308 21764 -14302
rect 20622 -14314 20802 -14308
rect 19926 -14496 19960 -14480
rect 19994 -14500 20010 -14314
rect 20786 -14384 20802 -14314
rect 20854 -14314 21764 -14308
rect 20854 -14330 20920 -14314
rect 20904 -14348 20920 -14330
rect 21696 -14330 21764 -14314
rect 21696 -14348 21712 -14330
rect 20786 -14404 21712 -14384
rect 20786 -14444 20920 -14404
rect 20786 -14500 20802 -14444
rect 19994 -14524 20802 -14500
rect 20836 -14496 20870 -14480
rect 20904 -14504 20920 -14444
rect 21696 -14504 21712 -14404
rect 20904 -14524 21712 -14504
rect 21746 -14496 21780 -14480
rect 19960 -14602 20836 -14576
rect 19960 -14750 19998 -14602
rect 20798 -14750 20836 -14602
rect 19960 -14776 20836 -14750
rect 20870 -14600 21746 -14576
rect 20870 -14748 20908 -14600
rect 21708 -14748 21746 -14600
rect 20870 -14776 21746 -14748
rect 19926 -14880 19960 -14864
rect 19994 -14854 20802 -14838
rect 19994 -14962 20008 -14854
rect 20788 -14920 20802 -14854
rect 21780 -14776 21782 -14576
rect 20836 -14880 20870 -14864
rect 20904 -14854 21712 -14838
rect 20904 -14920 20920 -14854
rect 20788 -14962 20920 -14920
rect 21700 -14962 21712 -14854
rect 21746 -14880 21780 -14864
rect 19994 -14978 21712 -14962
rect 19994 -15014 20010 -15012
rect 19822 -15046 20010 -15014
rect 20786 -15014 20802 -15012
rect 20904 -15014 20920 -15012
rect 20786 -15046 20920 -15014
rect 21696 -15014 21712 -15012
rect 21816 -15014 21884 -13874
rect 21696 -15046 21884 -15014
rect 19822 -15074 21884 -15046
rect 19822 -15442 19926 -15074
rect 19960 -15442 20836 -15074
rect 20870 -15442 21746 -15074
rect 21780 -15442 21884 -15074
rect 19822 -15470 21884 -15442
rect 19822 -15504 20010 -15470
rect 20786 -15504 20920 -15470
rect 21696 -15504 21884 -15470
rect 19822 -15542 21884 -15504
rect 21918 -13886 21956 -13874
rect 19494 -15548 21918 -15542
rect 19494 -18114 19534 -15548
rect 21862 -15638 21918 -15548
rect 20220 -15910 21532 -15878
rect 20220 -15944 20350 -15910
rect 21378 -15944 21532 -15910
rect 20220 -16006 20288 -15944
rect 20220 -16020 20254 -16006
rect 20222 -17992 20254 -16020
rect 1844 -18128 19534 -18114
rect 20220 -18012 20254 -17992
rect 20462 -16008 21266 -15944
rect 20462 -16044 20474 -16008
rect 21252 -16044 21266 -16008
rect 21440 -16006 21532 -15944
rect 20460 -16078 20474 -16044
rect 21252 -16078 21268 -16044
rect 20392 -16106 20426 -16090
rect 20392 -16190 20426 -16174
rect 20462 -16202 20474 -16078
rect 21252 -16202 21266 -16078
rect 21302 -16106 21336 -16090
rect 21302 -16190 21336 -16174
rect 20460 -16236 20474 -16202
rect 21252 -16236 21268 -16202
rect 20392 -16264 20426 -16248
rect 20462 -16268 20474 -16236
rect 21252 -16268 21266 -16236
rect 20462 -16284 21266 -16268
rect 21302 -16264 21336 -16248
rect 20392 -16348 20426 -16332
rect 20464 -16332 21264 -16318
rect 20464 -16360 20476 -16332
rect 21252 -16360 21264 -16332
rect 21302 -16348 21336 -16332
rect 20460 -16394 20476 -16360
rect 21252 -16394 21268 -16360
rect 20392 -16422 20426 -16406
rect 20464 -16424 20476 -16394
rect 21252 -16424 21264 -16394
rect 20464 -16436 21264 -16424
rect 21302 -16422 21336 -16406
rect 20392 -16506 20426 -16490
rect 20464 -16490 21264 -16476
rect 20464 -16518 20476 -16490
rect 21252 -16518 21264 -16490
rect 21302 -16506 21336 -16490
rect 20460 -16552 20476 -16518
rect 21252 -16552 21268 -16518
rect 20392 -16580 20426 -16564
rect 20464 -16582 20476 -16552
rect 21252 -16582 21264 -16552
rect 20464 -16594 21264 -16582
rect 21302 -16580 21336 -16564
rect 20392 -16664 20426 -16648
rect 20464 -16648 21264 -16634
rect 20464 -16676 20476 -16648
rect 21252 -16676 21264 -16648
rect 21302 -16664 21336 -16648
rect 20460 -16710 20476 -16676
rect 21252 -16710 21268 -16676
rect 20392 -16738 20426 -16722
rect 20464 -16740 20476 -16710
rect 21252 -16740 21264 -16710
rect 20464 -16752 21264 -16740
rect 21302 -16738 21336 -16722
rect 20392 -16822 20426 -16806
rect 20464 -16806 21264 -16792
rect 20464 -16834 20476 -16806
rect 21252 -16834 21264 -16806
rect 21302 -16822 21336 -16806
rect 20460 -16868 20476 -16834
rect 21252 -16868 21268 -16834
rect 20392 -16896 20426 -16880
rect 20464 -16898 20476 -16868
rect 21252 -16898 21264 -16868
rect 20464 -16910 21264 -16898
rect 21302 -16896 21336 -16880
rect 20392 -16980 20426 -16964
rect 20464 -16964 21264 -16950
rect 20464 -16992 20476 -16964
rect 21252 -16992 21264 -16964
rect 21302 -16980 21336 -16964
rect 20460 -17026 20476 -16992
rect 21252 -17026 21268 -16992
rect 20392 -17054 20426 -17038
rect 20464 -17056 20476 -17026
rect 21252 -17056 21264 -17026
rect 20464 -17068 21264 -17056
rect 21302 -17054 21336 -17038
rect 20392 -17138 20426 -17122
rect 20464 -17122 21264 -17108
rect 20464 -17150 20476 -17122
rect 21252 -17150 21264 -17122
rect 21302 -17138 21336 -17122
rect 20460 -17184 20476 -17150
rect 21252 -17184 21268 -17150
rect 20392 -17212 20426 -17196
rect 20464 -17214 20476 -17184
rect 21252 -17214 21264 -17184
rect 20464 -17226 21264 -17214
rect 21302 -17212 21336 -17196
rect 20392 -17296 20426 -17280
rect 20464 -17280 21264 -17266
rect 20464 -17308 20476 -17280
rect 21252 -17308 21264 -17280
rect 21302 -17296 21336 -17280
rect 20460 -17342 20476 -17308
rect 21252 -17342 21268 -17308
rect 20392 -17370 20426 -17354
rect 20464 -17372 20476 -17342
rect 21252 -17372 21264 -17342
rect 20464 -17384 21264 -17372
rect 21302 -17370 21336 -17354
rect 20392 -17454 20426 -17438
rect 20464 -17438 21264 -17424
rect 20464 -17466 20476 -17438
rect 21252 -17466 21264 -17438
rect 21302 -17454 21336 -17438
rect 20460 -17500 20476 -17466
rect 21252 -17500 21268 -17466
rect 20392 -17528 20426 -17512
rect 20464 -17530 20476 -17500
rect 21252 -17530 21264 -17500
rect 20464 -17542 21264 -17530
rect 21302 -17528 21336 -17512
rect 20392 -17612 20426 -17596
rect 20464 -17596 21264 -17582
rect 20464 -17624 20476 -17596
rect 21252 -17624 21264 -17596
rect 21302 -17612 21336 -17596
rect 20460 -17658 20476 -17624
rect 21252 -17658 21268 -17624
rect 20392 -17686 20426 -17670
rect 20464 -17688 20476 -17658
rect 21252 -17688 21264 -17658
rect 20464 -17700 21264 -17688
rect 21302 -17686 21336 -17670
rect 20392 -17770 20426 -17754
rect 20462 -17756 21266 -17734
rect 20462 -17782 20472 -17756
rect 21252 -17782 21266 -17756
rect 21302 -17770 21336 -17754
rect 20460 -17816 20472 -17782
rect 21252 -17816 21268 -17782
rect 20392 -17844 20426 -17828
rect 20392 -17928 20426 -17912
rect 20462 -17940 20472 -17816
rect 21252 -17940 21266 -17816
rect 21302 -17844 21336 -17828
rect 21302 -17928 21336 -17912
rect 20460 -17974 20472 -17940
rect 21252 -17974 21268 -17940
rect 20462 -17996 20472 -17974
rect 20462 -18010 20474 -17996
rect 21252 -18010 21266 -17974
rect 20462 -18012 21266 -18010
rect 21474 -16254 21532 -16006
rect 21862 -16254 21914 -15638
rect 21474 -18012 21914 -16254
rect 22120 -17862 22382 -12670
rect 22416 -12708 24514 -12670
rect 22416 -12714 22613 -12708
rect 22596 -12742 22613 -12714
rect 23389 -12714 23541 -12708
rect 23389 -12742 23405 -12714
rect 23524 -12742 23541 -12714
rect 24317 -12714 24514 -12708
rect 24317 -12742 24333 -12714
rect 22520 -12770 22554 -12754
rect 22452 -13138 22520 -12794
rect 22452 -13348 22554 -13138
rect 22452 -13716 22520 -13348
rect 22596 -13092 23404 -12742
rect 22596 -13392 22608 -13092
rect 23388 -13138 23404 -13092
rect 23390 -13166 23404 -13138
rect 23448 -12770 23482 -12754
rect 23390 -13200 23405 -13166
rect 23390 -13286 23404 -13200
rect 23390 -13320 23405 -13286
rect 23390 -13344 23404 -13320
rect 23388 -13392 23404 -13344
rect 22596 -13402 23404 -13392
rect 23448 -13348 23482 -13138
rect 22554 -13586 23448 -13486
rect 22452 -13926 22554 -13716
rect 22452 -14294 22520 -13926
rect 22594 -13668 23402 -13656
rect 22594 -13968 22610 -13668
rect 23390 -13702 23402 -13668
rect 23524 -13090 24332 -12742
rect 23524 -13390 23538 -13090
rect 24318 -13166 24332 -13090
rect 24376 -12770 24410 -12754
rect 24410 -13138 24478 -12794
rect 24318 -13200 24333 -13166
rect 24318 -13286 24332 -13200
rect 24318 -13320 24333 -13286
rect 24318 -13390 24332 -13320
rect 23524 -13402 24332 -13390
rect 24376 -13348 24478 -13138
rect 23482 -13586 24376 -13486
rect 23390 -13744 23404 -13702
rect 23390 -13778 23405 -13744
rect 23390 -13864 23404 -13778
rect 23390 -13898 23405 -13864
rect 23390 -13942 23404 -13898
rect 23448 -13926 23482 -13716
rect 23390 -13968 23402 -13942
rect 22594 -13980 23402 -13968
rect 22554 -14156 23448 -14056
rect 22452 -14504 22554 -14294
rect 22452 -14872 22520 -14504
rect 22596 -14242 23404 -14230
rect 22596 -14542 22608 -14242
rect 23388 -14298 23404 -14242
rect 23390 -14322 23404 -14298
rect 23520 -13666 24328 -13656
rect 23520 -13966 23536 -13666
rect 24316 -13702 24328 -13666
rect 24316 -13716 24330 -13702
rect 24318 -13744 24330 -13716
rect 24410 -13716 24478 -13348
rect 24318 -13778 24333 -13744
rect 24318 -13864 24332 -13778
rect 24318 -13898 24333 -13864
rect 24318 -13922 24330 -13898
rect 24316 -13942 24330 -13922
rect 24376 -13926 24478 -13716
rect 24316 -13966 24328 -13942
rect 23520 -13980 24328 -13966
rect 23482 -14156 24376 -14056
rect 23390 -14356 23405 -14322
rect 23390 -14442 23404 -14356
rect 23390 -14476 23405 -14442
rect 23390 -14504 23404 -14476
rect 23388 -14542 23404 -14504
rect 22596 -14554 23404 -14542
rect 23448 -14504 23482 -14294
rect 22554 -14732 23448 -14632
rect 22452 -15082 22554 -14872
rect 22596 -14814 23404 -14802
rect 22596 -14976 22610 -14814
rect 23390 -14900 23404 -14814
rect 23524 -14238 24332 -14230
rect 23524 -14538 23538 -14238
rect 24318 -14322 24332 -14238
rect 24410 -14294 24478 -13926
rect 24318 -14356 24333 -14322
rect 24318 -14442 24332 -14356
rect 24318 -14476 24333 -14442
rect 24318 -14538 24332 -14476
rect 23524 -14554 24332 -14538
rect 24376 -14504 24478 -14294
rect 23482 -14732 24376 -14632
rect 23390 -14934 23405 -14900
rect 23390 -14976 23404 -14934
rect 22596 -14982 23404 -14976
rect 22597 -15054 22613 -15020
rect 23389 -15054 23405 -15020
rect 22452 -15450 22520 -15082
rect 22452 -15560 22554 -15450
rect 22598 -15478 23404 -15054
rect 23448 -15082 23482 -14872
rect 24410 -14872 24478 -14504
rect 22597 -15512 22613 -15478
rect 23389 -15512 23405 -15478
rect 23448 -15560 23482 -15450
rect 22452 -15598 23482 -15560
rect 22452 -15642 22612 -15598
rect 23390 -15642 23482 -15598
rect 23524 -14900 24332 -14894
rect 23524 -14934 23541 -14900
rect 24317 -14934 24333 -14900
rect 23524 -15020 23570 -14934
rect 24284 -15020 24332 -14934
rect 23524 -15054 23541 -15020
rect 24317 -15054 24333 -15020
rect 23524 -15478 23570 -15054
rect 24284 -15478 24332 -15054
rect 24376 -15082 24478 -14872
rect 24410 -15450 24478 -15082
rect 23524 -15512 23541 -15478
rect 24317 -15512 24333 -15478
rect 23524 -15598 23570 -15512
rect 24284 -15598 24332 -15512
rect 23524 -15632 23541 -15598
rect 24317 -15632 24333 -15598
rect 23524 -15638 24332 -15632
rect 22452 -15660 22610 -15642
rect 22452 -16028 22520 -15660
rect 22554 -15914 22610 -15660
rect 23392 -15660 23482 -15642
rect 23392 -15914 23448 -15660
rect 22554 -15940 23448 -15914
rect 22452 -16238 22554 -16028
rect 22452 -16606 22520 -16238
rect 22596 -15988 23404 -15978
rect 22596 -16288 22610 -15988
rect 23390 -16056 23404 -15988
rect 24376 -15660 24478 -15450
rect 23482 -15888 24376 -15788
rect 23390 -16090 23405 -16056
rect 23390 -16176 23404 -16090
rect 23390 -16210 23405 -16176
rect 23390 -16288 23404 -16210
rect 22596 -16302 23404 -16288
rect 23448 -16238 23482 -16028
rect 22554 -16466 23448 -16366
rect 22452 -16816 22554 -16606
rect 22452 -17184 22520 -16816
rect 22596 -16552 23404 -16540
rect 22596 -16852 22610 -16552
rect 23390 -16634 23404 -16552
rect 23522 -15988 24330 -15978
rect 23522 -16288 23538 -15988
rect 24318 -16056 24330 -15988
rect 24410 -16028 24478 -15660
rect 24318 -16090 24333 -16056
rect 24318 -16176 24332 -16090
rect 24318 -16210 24333 -16176
rect 24318 -16288 24330 -16210
rect 23522 -16302 24330 -16288
rect 24376 -16238 24478 -16028
rect 23482 -16466 24376 -16366
rect 23390 -16668 23405 -16634
rect 23390 -16754 23404 -16668
rect 23390 -16788 23405 -16754
rect 23390 -16852 23404 -16788
rect 22596 -16864 23404 -16852
rect 23448 -16816 23482 -16606
rect 22554 -17040 23448 -16940
rect 22452 -17394 22554 -17184
rect 22452 -17736 22520 -17394
rect 22520 -17778 22554 -17762
rect 22596 -17138 23404 -17126
rect 22596 -17438 22610 -17138
rect 23390 -17212 23404 -17138
rect 23524 -16552 24332 -16540
rect 23524 -16852 23536 -16552
rect 24316 -16606 24332 -16552
rect 24318 -16634 24332 -16606
rect 24410 -16606 24478 -16238
rect 24318 -16668 24333 -16634
rect 24318 -16754 24332 -16668
rect 24318 -16788 24333 -16754
rect 24318 -16812 24332 -16788
rect 24316 -16852 24332 -16812
rect 23524 -16864 24332 -16852
rect 24376 -16816 24478 -16606
rect 23482 -17040 24376 -16940
rect 23390 -17246 23405 -17212
rect 23390 -17332 23404 -17246
rect 23390 -17366 23405 -17332
rect 23390 -17438 23404 -17366
rect 22596 -17790 23404 -17438
rect 23448 -17394 23482 -17184
rect 23448 -17778 23482 -17762
rect 23524 -17136 24332 -17126
rect 23524 -17436 23538 -17136
rect 24318 -17212 24332 -17136
rect 24410 -17184 24478 -16816
rect 24318 -17246 24333 -17212
rect 24318 -17332 24332 -17246
rect 24318 -17366 24333 -17332
rect 24318 -17436 24332 -17366
rect 23524 -17790 24332 -17436
rect 24376 -17394 24478 -17184
rect 24410 -17736 24478 -17394
rect 24376 -17778 24410 -17762
rect 22596 -17820 22613 -17790
rect 22416 -17824 22613 -17820
rect 23389 -17820 23405 -17790
rect 23524 -17820 23541 -17790
rect 23389 -17824 23541 -17820
rect 24317 -17820 24333 -17790
rect 24317 -17824 24514 -17820
rect 22416 -17862 24514 -17824
rect 24548 -17862 24616 -12670
rect 22120 -17924 24616 -17862
rect 25428 -17924 25479 -11672
rect 22120 -17958 22478 -17924
rect 24452 -17958 25479 -17924
rect 22120 -17984 25479 -17958
rect 20220 -18074 21914 -18012
rect 20220 -18108 20350 -18074
rect 21378 -18108 21914 -18074
rect 1844 -18408 1996 -18128
rect 18346 -18176 18856 -18128
rect 20220 -18184 21914 -18108
rect 18346 -18320 18856 -18210
rect 20220 -18320 24962 -18184
rect 24996 -18354 25092 -18320
rect 18346 -18408 18856 -18354
rect 1844 -18416 19534 -18408
rect 1844 -22538 2000 -18416
rect 2034 -18450 19534 -18416
rect 2034 -18516 2130 -18450
rect 2562 -18466 19534 -18450
rect 20220 -18416 25092 -18354
rect 20220 -18450 25058 -18416
rect 20220 -18466 24530 -18450
rect 2562 -18516 24530 -18466
rect 2562 -18518 2564 -18516
rect 24528 -18520 24530 -18516
rect 24962 -18516 25058 -18450
rect 2562 -18686 2564 -18616
rect 2130 -18782 2564 -18686
rect 2562 -18850 2564 -18782
rect 24962 -18852 24964 -18782
rect 24530 -18948 24964 -18852
rect 2562 -19018 2564 -18950
rect 24962 -19016 24964 -18948
rect 2130 -19114 2564 -19018
rect 2562 -19184 2564 -19114
rect 24962 -19184 24964 -19114
rect 24530 -19280 24964 -19184
rect 2562 -19350 2564 -19280
rect 24962 -19348 24964 -19280
rect 2130 -19446 2564 -19350
rect 2562 -19514 2564 -19446
rect 24962 -19516 24964 -19446
rect 24530 -19612 24964 -19516
rect 2562 -19682 2564 -19612
rect 24962 -19680 24964 -19612
rect 2130 -19778 2564 -19682
rect 2562 -19846 2564 -19778
rect 24962 -19848 24964 -19778
rect 24530 -19944 24964 -19848
rect 2562 -20014 2564 -19946
rect 24962 -20012 24964 -19944
rect 2130 -20110 2564 -20014
rect 2562 -20180 2564 -20110
rect 24962 -20180 24964 -20110
rect 24530 -20276 24964 -20180
rect 2562 -20346 2564 -20276
rect 24962 -20344 24964 -20276
rect 2130 -20442 2564 -20346
rect 2562 -20510 2564 -20442
rect 24962 -20512 24964 -20442
rect 24530 -20608 24964 -20512
rect 2562 -20678 2564 -20608
rect 24962 -20676 24964 -20608
rect 2130 -20774 2564 -20678
rect 2562 -20842 2564 -20774
rect 24962 -20844 24964 -20774
rect 24530 -20940 24964 -20844
rect 2128 -21010 2130 -20940
rect 24962 -21008 24964 -20940
rect 2128 -21106 2562 -21010
rect 2128 -21174 2130 -21106
rect 24528 -21176 24530 -21108
rect 24528 -21272 24962 -21176
rect 2562 -21342 2564 -21272
rect 24528 -21342 24530 -21272
rect 2130 -21438 2564 -21342
rect 2562 -21506 2564 -21438
rect 24962 -21508 24964 -21438
rect 24530 -21604 24964 -21508
rect 2562 -21674 2564 -21604
rect 24962 -21672 24964 -21604
rect 2130 -21770 2564 -21674
rect 2562 -21838 2564 -21770
rect 24528 -21840 24530 -21770
rect 24528 -21936 24962 -21840
rect 2128 -22006 2130 -21936
rect 24528 -22004 24530 -21936
rect 2128 -22102 2562 -22006
rect 2128 -22170 2130 -22102
rect 24528 -22172 24530 -22104
rect 24528 -22268 24962 -22172
rect 24528 -22338 24530 -22268
rect 2562 -22504 2564 -22444
rect 2130 -22518 2564 -22504
rect 24962 -22504 24964 -22442
rect 24530 -22518 24964 -22504
rect 2034 -22538 25058 -22518
rect 1844 -22600 25092 -22538
rect 1844 -22634 2096 -22600
rect 24996 -22634 25092 -22600
rect 1844 -22690 23876 -22634
rect 1844 -22710 21172 -22690
rect 1844 -23440 1890 -22710
rect 20268 -22724 21172 -22710
rect 21550 -22692 23876 -22690
rect 21550 -22724 22598 -22692
rect 20268 -22786 21110 -22724
rect 20268 -22838 21076 -22786
rect 20268 -22872 20454 -22838
rect 20556 -22872 21076 -22838
rect 20268 -22934 20392 -22872
rect 20268 -23036 20358 -22934
rect 20618 -22934 21076 -22872
rect 20456 -23018 20472 -22952
rect 20538 -23018 20554 -22952
rect 20268 -23098 20392 -23036
rect 20652 -23036 21076 -22934
rect 20618 -23098 21076 -23036
rect 20268 -23132 20454 -23098
rect 20556 -23132 21076 -23098
rect 20268 -23164 21076 -23132
rect 21612 -22726 22598 -22724
rect 22976 -22726 23876 -22692
rect 25198 -22706 25479 -17984
rect 21612 -22786 22536 -22726
rect 21214 -22862 21310 -22828
rect 21412 -22862 21482 -22828
rect 21214 -22924 21248 -22862
rect 21474 -22924 21482 -22862
rect 21312 -23008 21328 -22942
rect 21394 -23008 21410 -22942
rect 21214 -23088 21248 -23026
rect 21474 -23088 21482 -23026
rect 21214 -23096 21310 -23088
rect 21412 -23096 21482 -23088
rect 21214 -23158 21226 -23096
rect 20268 -23226 21110 -23164
rect 21646 -22788 22536 -22786
rect 21646 -22982 22502 -22788
rect 21612 -23226 21646 -23164
rect 20268 -23260 21172 -23226
rect 21550 -23260 21646 -23226
rect 21744 -23090 22390 -23068
rect 20268 -23440 21092 -23260
rect 21744 -23348 21764 -23090
rect 1844 -23486 21092 -23440
rect 1683 -23613 1717 -23587
rect 21288 -23598 21764 -23348
rect 22366 -23348 22390 -23090
rect 23038 -22788 23876 -22726
rect 22666 -22864 22736 -22830
rect 22838 -22864 22934 -22830
rect 22666 -22926 22674 -22864
rect 22900 -22926 22934 -22864
rect 22738 -23010 22754 -22944
rect 22820 -23010 22836 -22944
rect 22666 -23090 22674 -23028
rect 22900 -23090 22934 -23028
rect 22666 -23098 22736 -23090
rect 22838 -23098 22934 -23090
rect 22922 -23124 22934 -23098
rect 22922 -23160 22928 -23124
rect 22502 -23228 22536 -23166
rect 23072 -22840 23876 -22788
rect 23072 -22874 23562 -22840
rect 23664 -22874 23876 -22840
rect 23072 -22936 23500 -22874
rect 23072 -22982 23466 -22936
rect 23726 -22936 23876 -22874
rect 23564 -23020 23580 -22954
rect 23646 -23020 23662 -22954
rect 23466 -23100 23500 -23038
rect 23760 -22980 23876 -22936
rect 24040 -22730 25479 -22706
rect 23726 -23100 23760 -23038
rect 23466 -23134 23562 -23100
rect 23664 -23134 23760 -23100
rect 23038 -23228 23072 -23166
rect 24040 -23206 24070 -22730
rect 22502 -23262 22598 -23228
rect 22976 -23262 23072 -23228
rect 23168 -23348 24070 -23206
rect 22366 -23568 24070 -23348
rect 25410 -23568 25479 -22730
rect 22366 -23587 25479 -23568
rect 22366 -23598 25513 -23587
rect 21288 -23613 25513 -23598
rect 1683 -23647 1743 -23613
rect 25453 -23647 25513 -23613
<< viali >>
rect 2748 -946 2806 -864
rect 2748 -1048 2786 -946
rect 2786 -1048 2806 -946
rect 2900 -1030 2966 -964
rect 2748 -1128 2806 -1048
rect 2748 -1144 2882 -1128
rect 2882 -1144 2984 -1128
rect 2984 -1144 3018 -1128
rect 2748 -1182 3018 -1144
rect 3156 -1180 3236 -956
rect 5096 -1180 5176 -958
rect 5530 -946 5586 -884
rect 5370 -1030 5436 -964
rect 5530 -1048 5550 -946
rect 5550 -1048 5586 -946
rect 5530 -1126 5586 -1048
rect 5316 -1144 5352 -1126
rect 5352 -1144 5454 -1126
rect 5454 -1144 5586 -1126
rect 5316 -1180 5586 -1144
rect 2933 -1295 2967 -1261
rect 2933 -1387 2967 -1353
rect 3477 -1295 3511 -1261
rect 2933 -1479 2967 -1445
rect 3477 -1387 3511 -1353
rect 3477 -1479 3511 -1445
rect 2933 -1571 2967 -1537
rect 3477 -1571 3511 -1537
rect 4819 -1295 4853 -1261
rect 5363 -1295 5397 -1261
rect 4819 -1387 4853 -1353
rect 4819 -1479 4853 -1445
rect 5363 -1387 5397 -1353
rect 5363 -1479 5397 -1445
rect 4819 -1571 4853 -1537
rect 5363 -1571 5397 -1537
rect 3050 -1768 3412 -1694
rect 4916 -1760 5278 -1686
rect 13676 -1752 13848 -1580
rect 13971 -1721 14005 -1687
rect 14515 -1721 14549 -1687
rect 13971 -1813 14005 -1779
rect 13971 -1905 14005 -1871
rect 2652 -1982 2748 -1948
rect 2652 -2044 2686 -1982
rect 2652 -2400 2686 -2044
rect 2828 -2084 2996 -2050
rect 2766 -2310 2800 -2134
rect 3024 -2310 3058 -2134
rect 2828 -2394 2996 -2360
rect 2652 -2462 2686 -2400
rect 2652 -2496 2748 -2462
rect 3676 -1974 3772 -1940
rect 3738 -2036 3772 -1974
rect 3428 -2076 3596 -2042
rect 3366 -2311 3400 -2135
rect 3624 -2311 3658 -2135
rect 3428 -2404 3596 -2370
rect 3738 -2410 3772 -2036
rect 3738 -2472 3772 -2410
rect 3676 -2506 3772 -2472
rect 4564 -1974 4660 -1940
rect 4564 -2036 4598 -1974
rect 4564 -2410 4598 -2036
rect 4740 -2076 4908 -2042
rect 4678 -2311 4712 -2135
rect 4936 -2311 4970 -2135
rect 4740 -2404 4908 -2370
rect 4564 -2472 4598 -2410
rect 4564 -2506 4660 -2472
rect 5588 -1982 5684 -1948
rect 5650 -2044 5684 -1982
rect 5340 -2084 5508 -2050
rect 5278 -2310 5312 -2134
rect 5536 -2310 5570 -2134
rect 5340 -2394 5508 -2360
rect 5650 -2400 5684 -2044
rect 5650 -2462 5684 -2400
rect 5588 -2496 5684 -2462
rect 7514 -2106 9032 -2082
rect 7514 -2128 7538 -2106
rect 7538 -2128 7606 -2106
rect 7606 -2128 7696 -2106
rect 7696 -2128 7764 -2106
rect 7764 -2128 7854 -2106
rect 7854 -2128 7922 -2106
rect 7922 -2128 8012 -2106
rect 8012 -2128 8080 -2106
rect 8080 -2128 8170 -2106
rect 8170 -2128 8238 -2106
rect 8238 -2128 8328 -2106
rect 8328 -2128 8396 -2106
rect 8396 -2128 8486 -2106
rect 8486 -2128 8554 -2106
rect 8554 -2128 8644 -2106
rect 8644 -2128 8712 -2106
rect 8712 -2128 8802 -2106
rect 8802 -2128 8870 -2106
rect 8870 -2128 8960 -2106
rect 8960 -2128 9028 -2106
rect 9028 -2128 9032 -2106
rect 7444 -2199 7540 -2198
rect 7444 -2975 7476 -2199
rect 7476 -2975 7510 -2199
rect 7510 -2975 7540 -2199
rect 7444 -2976 7540 -2975
rect 7604 -2199 7700 -2198
rect 7604 -2975 7634 -2199
rect 7634 -2975 7668 -2199
rect 7668 -2975 7700 -2199
rect 7604 -2976 7700 -2975
rect 7762 -2199 7858 -2198
rect 7762 -2975 7792 -2199
rect 7792 -2975 7826 -2199
rect 7826 -2975 7858 -2199
rect 7762 -2976 7858 -2975
rect 7920 -2199 8016 -2198
rect 7920 -2975 7950 -2199
rect 7950 -2975 7984 -2199
rect 7984 -2975 8016 -2199
rect 7920 -2976 8016 -2975
rect 8078 -2199 8174 -2198
rect 8078 -2975 8108 -2199
rect 8108 -2975 8142 -2199
rect 8142 -2975 8174 -2199
rect 8078 -2976 8174 -2975
rect 8234 -2199 8330 -2198
rect 8234 -2975 8266 -2199
rect 8266 -2975 8300 -2199
rect 8300 -2975 8330 -2199
rect 8234 -2976 8330 -2975
rect 8392 -2199 8488 -2198
rect 8392 -2975 8424 -2199
rect 8424 -2975 8458 -2199
rect 8458 -2975 8488 -2199
rect 8392 -2976 8488 -2975
rect 8552 -2199 8648 -2198
rect 8552 -2975 8582 -2199
rect 8582 -2975 8616 -2199
rect 8616 -2975 8648 -2199
rect 8552 -2976 8648 -2975
rect 8708 -2199 8804 -2198
rect 8708 -2975 8740 -2199
rect 8740 -2975 8774 -2199
rect 8774 -2975 8804 -2199
rect 8708 -2976 8804 -2975
rect 8866 -2199 8962 -2198
rect 8866 -2975 8898 -2199
rect 8898 -2975 8932 -2199
rect 8932 -2975 8962 -2199
rect 8866 -2976 8962 -2975
rect 9024 -2199 9120 -2198
rect 9024 -2975 9056 -2199
rect 9056 -2975 9090 -2199
rect 9090 -2975 9120 -2199
rect 9024 -2976 9120 -2975
rect 7512 -3068 7538 -3046
rect 7538 -3068 7606 -3046
rect 7606 -3068 7696 -3046
rect 7696 -3068 7764 -3046
rect 7764 -3068 7854 -3046
rect 7854 -3068 7922 -3046
rect 7922 -3068 8012 -3046
rect 8012 -3068 8080 -3046
rect 8080 -3068 8170 -3046
rect 8170 -3068 8238 -3046
rect 8238 -3068 8328 -3046
rect 8328 -3068 8396 -3046
rect 8396 -3068 8486 -3046
rect 8486 -3068 8554 -3046
rect 8554 -3068 8644 -3046
rect 8644 -3068 8712 -3046
rect 8712 -3068 8802 -3046
rect 8802 -3068 8870 -3046
rect 8870 -3068 8960 -3046
rect 8960 -3068 9028 -3046
rect 9028 -3068 9034 -3046
rect 7512 -3092 9034 -3068
rect 9438 -2120 10952 -2092
rect 9438 -2140 9464 -2120
rect 9464 -2140 9532 -2120
rect 9532 -2140 9622 -2120
rect 9622 -2140 9690 -2120
rect 9690 -2140 9780 -2120
rect 9780 -2140 9848 -2120
rect 9848 -2140 9938 -2120
rect 9938 -2140 10006 -2120
rect 10006 -2140 10096 -2120
rect 10096 -2140 10164 -2120
rect 10164 -2140 10254 -2120
rect 10254 -2140 10322 -2120
rect 10322 -2140 10412 -2120
rect 10412 -2140 10480 -2120
rect 10480 -2140 10570 -2120
rect 10570 -2140 10638 -2120
rect 10638 -2140 10728 -2120
rect 10728 -2140 10796 -2120
rect 10796 -2140 10886 -2120
rect 10886 -2140 10952 -2120
rect 9370 -2204 9466 -2202
rect 9370 -2980 9402 -2204
rect 9402 -2980 9436 -2204
rect 9436 -2980 9466 -2204
rect 9528 -2204 9624 -2202
rect 9528 -2980 9560 -2204
rect 9560 -2980 9594 -2204
rect 9594 -2980 9624 -2204
rect 9688 -2204 9784 -2202
rect 9688 -2980 9718 -2204
rect 9718 -2980 9752 -2204
rect 9752 -2980 9784 -2204
rect 9846 -2204 9942 -2202
rect 9846 -2980 9876 -2204
rect 9876 -2980 9910 -2204
rect 9910 -2980 9942 -2204
rect 10002 -2204 10098 -2202
rect 10002 -2980 10034 -2204
rect 10034 -2980 10068 -2204
rect 10068 -2980 10098 -2204
rect 10162 -2204 10258 -2202
rect 10162 -2980 10192 -2204
rect 10192 -2980 10226 -2204
rect 10226 -2980 10258 -2204
rect 10318 -2204 10414 -2202
rect 10318 -2980 10350 -2204
rect 10350 -2980 10384 -2204
rect 10384 -2980 10414 -2204
rect 10476 -2204 10572 -2202
rect 10476 -2980 10508 -2204
rect 10508 -2980 10542 -2204
rect 10542 -2980 10572 -2204
rect 10636 -2204 10732 -2202
rect 10636 -2980 10666 -2204
rect 10666 -2980 10700 -2204
rect 10700 -2980 10732 -2204
rect 10792 -2204 10888 -2202
rect 10792 -2980 10824 -2204
rect 10824 -2980 10858 -2204
rect 10858 -2980 10888 -2204
rect 10950 -2204 11046 -2202
rect 10950 -2980 10982 -2204
rect 10982 -2980 11016 -2204
rect 11016 -2980 11046 -2204
rect 9436 -3064 9464 -3044
rect 9464 -3064 9532 -3044
rect 9532 -3064 9622 -3044
rect 9622 -3064 9690 -3044
rect 9690 -3064 9780 -3044
rect 9780 -3064 9848 -3044
rect 9848 -3064 9938 -3044
rect 9938 -3064 10006 -3044
rect 10006 -3064 10096 -3044
rect 10096 -3064 10164 -3044
rect 10164 -3064 10254 -3044
rect 10254 -3064 10322 -3044
rect 10322 -3064 10412 -3044
rect 10412 -3064 10480 -3044
rect 10480 -3064 10570 -3044
rect 10570 -3064 10638 -3044
rect 10638 -3064 10728 -3044
rect 10728 -3064 10796 -3044
rect 10796 -3064 10886 -3044
rect 10886 -3064 10952 -3044
rect 9436 -3092 10952 -3064
rect 11496 -2122 11564 -2088
rect 11310 -2958 11334 -2180
rect 11334 -2181 11468 -2180
rect 11334 -2957 11434 -2181
rect 11434 -2957 11468 -2181
rect 11334 -2958 11468 -2957
rect 11606 -2956 11626 -2182
rect 11626 -2956 11666 -2182
rect 11496 -3050 11564 -3016
rect 13971 -1997 14005 -1963
rect 14897 -1767 14931 -1733
rect 14989 -1767 15023 -1733
rect 15081 -1767 15115 -1733
rect 15173 -1767 15207 -1733
rect 15265 -1767 15299 -1733
rect 15357 -1767 15391 -1733
rect 15449 -1767 15483 -1733
rect 15541 -1767 15575 -1733
rect 15633 -1767 15667 -1733
rect 15725 -1767 15759 -1733
rect 15817 -1767 15851 -1733
rect 15909 -1767 15943 -1733
rect 16001 -1767 16035 -1733
rect 16093 -1767 16127 -1733
rect 16185 -1767 16219 -1733
rect 16277 -1767 16311 -1733
rect 16369 -1767 16403 -1733
rect 16461 -1767 16495 -1733
rect 16553 -1767 16587 -1733
rect 16645 -1767 16679 -1733
rect 16737 -1767 16771 -1733
rect 16829 -1767 16863 -1733
rect 16921 -1767 16955 -1733
rect 17013 -1767 17047 -1733
rect 17105 -1767 17139 -1733
rect 17197 -1767 17231 -1733
rect 17289 -1767 17323 -1733
rect 17381 -1767 17415 -1733
rect 17473 -1767 17507 -1733
rect 17565 -1767 17599 -1733
rect 17657 -1767 17691 -1733
rect 17749 -1767 17783 -1733
rect 17841 -1767 17875 -1733
rect 17933 -1767 17967 -1733
rect 18025 -1767 18059 -1733
rect 18117 -1767 18151 -1733
rect 18209 -1767 18243 -1733
rect 18301 -1767 18335 -1733
rect 18393 -1767 18427 -1733
rect 18485 -1767 18519 -1733
rect 18577 -1767 18611 -1733
rect 18669 -1767 18703 -1733
rect 18761 -1767 18795 -1733
rect 18853 -1767 18887 -1733
rect 18945 -1767 18979 -1733
rect 19037 -1767 19071 -1733
rect 19129 -1767 19163 -1733
rect 19221 -1767 19255 -1733
rect 19313 -1767 19347 -1733
rect 19405 -1767 19439 -1733
rect 19497 -1767 19531 -1733
rect 19589 -1767 19623 -1733
rect 19681 -1767 19715 -1733
rect 19773 -1767 19807 -1733
rect 19865 -1767 19899 -1733
rect 19957 -1767 19991 -1733
rect 20049 -1767 20083 -1733
rect 20141 -1767 20175 -1733
rect 20233 -1767 20267 -1733
rect 20325 -1767 20359 -1733
rect 20417 -1767 20451 -1733
rect 20509 -1767 20543 -1733
rect 20601 -1767 20635 -1733
rect 20693 -1767 20727 -1733
rect 20785 -1767 20819 -1733
rect 20877 -1767 20911 -1733
rect 20969 -1767 21003 -1733
rect 21061 -1767 21095 -1733
rect 21153 -1767 21187 -1733
rect 21245 -1767 21279 -1733
rect 21337 -1767 21371 -1733
rect 21429 -1767 21463 -1733
rect 21521 -1767 21555 -1733
rect 21613 -1767 21647 -1733
rect 21705 -1767 21739 -1733
rect 21797 -1767 21831 -1733
rect 21889 -1767 21923 -1733
rect 21981 -1767 22015 -1733
rect 22073 -1767 22107 -1733
rect 14515 -1813 14549 -1779
rect 14204 -1911 14242 -1872
rect 14204 -1945 14237 -1911
rect 14237 -1945 14242 -1911
rect 14204 -1960 14242 -1945
rect 13971 -2089 14005 -2055
rect 12786 -2240 12862 -2206
rect 12702 -3036 12736 -2268
rect 12912 -3036 12946 -2268
rect 12786 -3098 12862 -3064
rect 13971 -2181 14005 -2147
rect 13971 -2273 14005 -2239
rect 14138 -2045 14203 -2040
rect 14203 -2045 14230 -2040
rect 14138 -2074 14230 -2045
rect 14136 -2160 14228 -2156
rect 14136 -2190 14203 -2160
rect 14203 -2190 14228 -2160
rect 13971 -2365 14005 -2331
rect 14204 -2267 14242 -2250
rect 14204 -2301 14237 -2267
rect 14237 -2301 14242 -2267
rect 14204 -2328 14242 -2301
rect 14515 -1905 14549 -1871
rect 14515 -1997 14549 -1963
rect 14515 -2089 14549 -2055
rect 14515 -2181 14549 -2147
rect 14515 -2273 14549 -2239
rect 14515 -2365 14549 -2331
rect 13052 -3026 13648 -2468
rect 13971 -2457 14005 -2423
rect 14515 -2457 14549 -2423
rect 13971 -2549 14005 -2515
rect 13971 -2641 14005 -2607
rect 14208 -2554 14308 -2472
rect 14208 -2572 14237 -2554
rect 14237 -2572 14308 -2554
rect 14515 -2549 14549 -2515
rect 14515 -2641 14549 -2607
rect 13971 -2733 14005 -2699
rect 13971 -2814 13978 -2791
rect 13978 -2814 14005 -2791
rect 13971 -2825 14005 -2814
rect 14515 -2733 14549 -2699
rect 14515 -2825 14549 -2791
rect 14040 -2982 14140 -2902
rect 14740 -2098 14812 -2026
rect 14980 -2008 15040 -1988
rect 14980 -2042 15012 -2008
rect 15012 -2042 15040 -2008
rect 14980 -2076 15040 -2042
rect 14980 -2110 15012 -2076
rect 15012 -2110 15040 -2076
rect 14980 -2140 15040 -2110
rect 15160 -2003 15164 -1986
rect 15164 -2003 15198 -1986
rect 15198 -2003 15200 -1986
rect 15160 -2037 15200 -2003
rect 15160 -2066 15164 -2037
rect 15164 -2066 15198 -2037
rect 15198 -2066 15200 -2037
rect 15634 -1980 15668 -1971
rect 15634 -2005 15646 -1980
rect 15646 -2005 15668 -1980
rect 15814 -2060 15853 -2036
rect 15853 -2060 15854 -2036
rect 15814 -2076 15854 -2060
rect 15715 -2125 15749 -2107
rect 15715 -2141 15749 -2125
rect 16001 -2005 16035 -1971
rect 16273 -1937 16307 -1903
rect 16345 -1919 16379 -1903
rect 16345 -1937 16369 -1919
rect 16369 -1937 16379 -1919
rect 16093 -2141 16127 -2107
rect 16717 -1989 16743 -1971
rect 16743 -1989 16751 -1971
rect 16717 -2005 16751 -1989
rect 16993 -1937 17027 -1903
rect 16933 -1991 16949 -1966
rect 16949 -1991 16967 -1966
rect 16933 -2000 16967 -1991
rect 16717 -2115 16748 -2107
rect 16748 -2115 16751 -2107
rect 16717 -2141 16751 -2115
rect 17556 -2088 17594 -2050
rect 17842 -1980 17876 -1971
rect 17842 -2005 17854 -1980
rect 17854 -2005 17876 -1980
rect 18022 -2060 18061 -2036
rect 18061 -2060 18062 -2036
rect 18022 -2076 18062 -2060
rect 17923 -2125 17957 -2107
rect 17923 -2141 17957 -2125
rect 18209 -2005 18243 -1971
rect 18481 -1937 18515 -1903
rect 18553 -1919 18587 -1903
rect 18553 -1937 18577 -1919
rect 18577 -1937 18587 -1919
rect 18301 -2141 18335 -2107
rect 18925 -1989 18951 -1971
rect 18951 -1989 18959 -1971
rect 18925 -2005 18959 -1989
rect 19201 -1937 19235 -1903
rect 19141 -1991 19157 -1966
rect 19157 -1991 19175 -1966
rect 19141 -2000 19175 -1991
rect 18925 -2115 18956 -2107
rect 18956 -2115 18959 -2107
rect 18925 -2141 18959 -2115
rect 19766 -2088 19804 -2050
rect 20050 -1980 20084 -1971
rect 20050 -2005 20062 -1980
rect 20062 -2005 20084 -1980
rect 20230 -2060 20269 -2036
rect 20269 -2060 20270 -2036
rect 20230 -2076 20270 -2060
rect 20131 -2125 20165 -2107
rect 20131 -2141 20165 -2125
rect 20417 -2005 20451 -1971
rect 20689 -1937 20723 -1903
rect 20761 -1919 20795 -1903
rect 20761 -1937 20785 -1919
rect 20785 -1937 20795 -1919
rect 20509 -2141 20543 -2107
rect 21133 -1989 21159 -1971
rect 21159 -1989 21167 -1971
rect 21133 -2005 21167 -1989
rect 21409 -1937 21443 -1903
rect 21349 -1991 21365 -1966
rect 21365 -1991 21383 -1966
rect 21349 -2000 21383 -1991
rect 21133 -2115 21164 -2107
rect 21164 -2115 21167 -2107
rect 21133 -2141 21167 -2115
rect 21974 -2097 22014 -1966
rect 21974 -2131 21998 -2097
rect 21998 -2131 22014 -2097
rect 21974 -2160 22014 -2131
rect 14897 -2311 14931 -2277
rect 14989 -2311 15023 -2277
rect 15081 -2311 15115 -2277
rect 15173 -2311 15207 -2277
rect 15265 -2311 15299 -2277
rect 15357 -2311 15391 -2277
rect 15449 -2311 15483 -2277
rect 15541 -2311 15575 -2277
rect 15633 -2311 15667 -2277
rect 15725 -2311 15759 -2277
rect 15817 -2311 15851 -2277
rect 15909 -2311 15943 -2277
rect 16001 -2311 16035 -2277
rect 16093 -2311 16127 -2277
rect 16185 -2311 16219 -2277
rect 16277 -2311 16311 -2277
rect 16369 -2311 16403 -2277
rect 16461 -2311 16495 -2277
rect 16553 -2311 16587 -2277
rect 16645 -2311 16679 -2277
rect 16737 -2311 16771 -2277
rect 16829 -2311 16863 -2277
rect 16921 -2311 16955 -2277
rect 17013 -2311 17047 -2277
rect 17105 -2311 17139 -2277
rect 17197 -2311 17231 -2277
rect 17289 -2311 17323 -2277
rect 17381 -2311 17415 -2277
rect 17473 -2311 17507 -2277
rect 17565 -2311 17599 -2277
rect 17657 -2311 17691 -2277
rect 17749 -2311 17783 -2277
rect 17841 -2311 17875 -2277
rect 17933 -2311 17967 -2277
rect 18025 -2311 18059 -2277
rect 18117 -2311 18151 -2277
rect 18209 -2311 18243 -2277
rect 18301 -2311 18335 -2277
rect 18393 -2311 18427 -2277
rect 18485 -2311 18519 -2277
rect 18577 -2311 18611 -2277
rect 18669 -2311 18703 -2277
rect 18761 -2311 18795 -2277
rect 18853 -2311 18887 -2277
rect 18945 -2311 18979 -2277
rect 19037 -2311 19071 -2277
rect 19129 -2311 19163 -2277
rect 19221 -2311 19255 -2277
rect 19313 -2311 19347 -2277
rect 19405 -2311 19439 -2277
rect 19497 -2311 19531 -2277
rect 19589 -2311 19623 -2277
rect 19681 -2311 19715 -2277
rect 19773 -2311 19807 -2277
rect 19865 -2311 19899 -2277
rect 19957 -2311 19991 -2277
rect 20049 -2311 20083 -2277
rect 20141 -2311 20175 -2277
rect 20233 -2311 20267 -2277
rect 20325 -2311 20359 -2277
rect 20417 -2311 20451 -2277
rect 20509 -2311 20543 -2277
rect 20601 -2311 20635 -2277
rect 20693 -2311 20727 -2277
rect 20785 -2311 20819 -2277
rect 20877 -2311 20911 -2277
rect 20969 -2311 21003 -2277
rect 21061 -2311 21095 -2277
rect 21153 -2311 21187 -2277
rect 21245 -2311 21279 -2277
rect 21337 -2311 21371 -2277
rect 21429 -2311 21463 -2277
rect 21521 -2311 21555 -2277
rect 21613 -2311 21647 -2277
rect 21705 -2311 21739 -2277
rect 21797 -2311 21831 -2277
rect 21889 -2311 21923 -2277
rect 21981 -2311 22015 -2277
rect 22073 -2311 22107 -2277
rect 14740 -2562 14812 -2490
rect 14414 -2982 14514 -2902
rect 14980 -2478 15040 -2448
rect 14980 -2512 15012 -2478
rect 15012 -2512 15040 -2478
rect 14980 -2546 15040 -2512
rect 14980 -2580 15012 -2546
rect 15012 -2580 15040 -2546
rect 14980 -2600 15040 -2580
rect 15160 -2551 15164 -2522
rect 15164 -2551 15198 -2522
rect 15198 -2551 15200 -2522
rect 15160 -2585 15200 -2551
rect 15160 -2602 15164 -2585
rect 15164 -2602 15198 -2585
rect 15198 -2602 15200 -2585
rect 15634 -2608 15646 -2583
rect 15646 -2608 15668 -2583
rect 15634 -2617 15668 -2608
rect 15715 -2463 15749 -2447
rect 15715 -2481 15749 -2463
rect 15814 -2528 15854 -2512
rect 15814 -2552 15853 -2528
rect 15853 -2552 15854 -2528
rect 16093 -2481 16127 -2447
rect 16001 -2617 16035 -2583
rect 16717 -2473 16751 -2447
rect 16717 -2481 16748 -2473
rect 16748 -2481 16751 -2473
rect 16273 -2685 16307 -2651
rect 16345 -2669 16369 -2651
rect 16369 -2669 16379 -2651
rect 16345 -2685 16379 -2669
rect 16717 -2599 16751 -2583
rect 16717 -2617 16743 -2599
rect 16743 -2617 16751 -2599
rect 16933 -2597 16967 -2588
rect 16933 -2622 16949 -2597
rect 16949 -2622 16967 -2597
rect 16993 -2685 17027 -2651
rect 17556 -2538 17594 -2500
rect 17842 -2608 17854 -2583
rect 17854 -2608 17876 -2583
rect 17842 -2617 17876 -2608
rect 17923 -2463 17957 -2447
rect 17923 -2481 17957 -2463
rect 18022 -2528 18062 -2512
rect 18022 -2552 18061 -2528
rect 18061 -2552 18062 -2528
rect 18301 -2481 18335 -2447
rect 18209 -2617 18243 -2583
rect 18925 -2473 18959 -2447
rect 18925 -2481 18956 -2473
rect 18956 -2481 18959 -2473
rect 18481 -2685 18515 -2651
rect 18553 -2669 18577 -2651
rect 18577 -2669 18587 -2651
rect 18553 -2685 18587 -2669
rect 18925 -2599 18959 -2583
rect 18925 -2617 18951 -2599
rect 18951 -2617 18959 -2599
rect 19141 -2597 19175 -2588
rect 19141 -2622 19157 -2597
rect 19157 -2622 19175 -2597
rect 19201 -2685 19235 -2651
rect 19766 -2538 19804 -2500
rect 20050 -2608 20062 -2583
rect 20062 -2608 20084 -2583
rect 20050 -2617 20084 -2608
rect 20131 -2463 20165 -2447
rect 20131 -2481 20165 -2463
rect 20230 -2528 20270 -2512
rect 20230 -2552 20269 -2528
rect 20269 -2552 20270 -2528
rect 20509 -2481 20543 -2447
rect 20417 -2617 20451 -2583
rect 21133 -2473 21167 -2447
rect 21133 -2481 21164 -2473
rect 21164 -2481 21167 -2473
rect 20689 -2685 20723 -2651
rect 20761 -2669 20785 -2651
rect 20785 -2669 20795 -2651
rect 20761 -2685 20795 -2669
rect 21133 -2599 21167 -2583
rect 21133 -2617 21159 -2599
rect 21159 -2617 21167 -2599
rect 21349 -2597 21383 -2588
rect 21349 -2622 21365 -2597
rect 21365 -2622 21383 -2597
rect 21409 -2685 21443 -2651
rect 21974 -2457 22014 -2428
rect 21974 -2491 21998 -2457
rect 21998 -2491 22014 -2457
rect 21974 -2622 22014 -2491
rect 14897 -2855 14931 -2821
rect 14989 -2855 15023 -2821
rect 15081 -2855 15115 -2821
rect 15173 -2855 15207 -2821
rect 15265 -2855 15299 -2821
rect 15357 -2855 15391 -2821
rect 15449 -2855 15483 -2821
rect 15541 -2855 15575 -2821
rect 15633 -2855 15667 -2821
rect 15725 -2855 15759 -2821
rect 15817 -2855 15851 -2821
rect 15909 -2855 15943 -2821
rect 16001 -2855 16035 -2821
rect 16093 -2855 16127 -2821
rect 16185 -2855 16219 -2821
rect 16277 -2855 16311 -2821
rect 16369 -2855 16403 -2821
rect 16461 -2855 16495 -2821
rect 16553 -2855 16587 -2821
rect 16645 -2855 16679 -2821
rect 16737 -2855 16771 -2821
rect 16829 -2855 16863 -2821
rect 16921 -2855 16955 -2821
rect 17013 -2855 17047 -2821
rect 17105 -2855 17139 -2821
rect 17197 -2855 17231 -2821
rect 17289 -2855 17323 -2821
rect 17381 -2855 17415 -2821
rect 17473 -2855 17507 -2821
rect 17565 -2855 17599 -2821
rect 17657 -2855 17691 -2821
rect 17749 -2855 17783 -2821
rect 17841 -2855 17875 -2821
rect 17933 -2855 17967 -2821
rect 18025 -2855 18059 -2821
rect 18117 -2855 18151 -2821
rect 18209 -2855 18243 -2821
rect 18301 -2855 18335 -2821
rect 18393 -2855 18427 -2821
rect 18485 -2855 18519 -2821
rect 18577 -2855 18611 -2821
rect 18669 -2855 18703 -2821
rect 18761 -2855 18795 -2821
rect 18853 -2855 18887 -2821
rect 18945 -2855 18979 -2821
rect 19037 -2855 19071 -2821
rect 19129 -2855 19163 -2821
rect 19221 -2855 19255 -2821
rect 19313 -2855 19347 -2821
rect 19405 -2855 19439 -2821
rect 19497 -2855 19531 -2821
rect 19589 -2855 19623 -2821
rect 19681 -2855 19715 -2821
rect 19773 -2855 19807 -2821
rect 19865 -2855 19899 -2821
rect 19957 -2855 19991 -2821
rect 20049 -2855 20083 -2821
rect 20141 -2855 20175 -2821
rect 20233 -2855 20267 -2821
rect 20325 -2855 20359 -2821
rect 20417 -2855 20451 -2821
rect 20509 -2855 20543 -2821
rect 20601 -2855 20635 -2821
rect 20693 -2855 20727 -2821
rect 20785 -2855 20819 -2821
rect 20877 -2855 20911 -2821
rect 20969 -2855 21003 -2821
rect 21061 -2855 21095 -2821
rect 21153 -2855 21187 -2821
rect 21245 -2855 21279 -2821
rect 21337 -2855 21371 -2821
rect 21429 -2855 21463 -2821
rect 21521 -2855 21555 -2821
rect 21613 -2855 21647 -2821
rect 21705 -2855 21739 -2821
rect 21797 -2855 21831 -2821
rect 21889 -2855 21923 -2821
rect 21981 -2855 22015 -2821
rect 22073 -2855 22107 -2821
rect 2456 -4012 2552 -3918
rect 2456 -4840 2548 -4012
rect 2548 -4840 2552 -4012
rect 3162 -4012 3258 -3916
rect 2744 -4088 2812 -4054
rect 2902 -4088 2970 -4054
rect 2682 -4714 2716 -4138
rect 2840 -4714 2874 -4138
rect 2998 -4714 3032 -4138
rect 2744 -4798 2812 -4764
rect 2902 -4798 2970 -4764
rect 2456 -4936 2552 -4840
rect 3162 -4840 3166 -4012
rect 3166 -4840 3254 -4012
rect 3254 -4840 3258 -4012
rect 3870 -4012 3966 -3916
rect 3450 -4088 3518 -4054
rect 3608 -4088 3676 -4054
rect 3388 -4714 3422 -4138
rect 3546 -4714 3580 -4138
rect 3704 -4714 3738 -4138
rect 3450 -4798 3518 -4764
rect 3608 -4798 3676 -4764
rect 3162 -4934 3258 -4840
rect 3870 -4840 3872 -4012
rect 3872 -4840 3966 -4012
rect 3870 -4934 3966 -4840
rect 4370 -4012 4466 -3916
rect 4370 -4840 4464 -4012
rect 4464 -4840 4466 -4012
rect 5078 -4012 5174 -3916
rect 4660 -4088 4728 -4054
rect 4818 -4088 4886 -4054
rect 4598 -4714 4632 -4138
rect 4756 -4714 4790 -4138
rect 4914 -4714 4948 -4138
rect 4660 -4798 4728 -4764
rect 4818 -4798 4886 -4764
rect 4370 -4934 4466 -4840
rect 5078 -4840 5082 -4012
rect 5082 -4840 5170 -4012
rect 5170 -4840 5174 -4012
rect 5784 -4012 5880 -3918
rect 5366 -4088 5434 -4054
rect 5524 -4088 5592 -4054
rect 5304 -4714 5338 -4138
rect 5462 -4714 5496 -4138
rect 5620 -4714 5654 -4138
rect 5366 -4798 5434 -4764
rect 5524 -4798 5592 -4764
rect 5078 -4934 5174 -4840
rect 5784 -4840 5788 -4012
rect 5788 -4840 5880 -4012
rect 5784 -4936 5880 -4840
rect 1990 -6772 2476 -5154
rect 2586 -5306 2706 -5174
rect 2586 -5752 2630 -5306
rect 2630 -5752 2664 -5306
rect 2664 -5752 2706 -5306
rect 2826 -5382 3594 -5348
rect 2764 -5617 2798 -5441
rect 3622 -5617 3656 -5441
rect 2826 -5710 3594 -5676
rect 2586 -5848 2706 -5752
rect 5630 -5306 5750 -5174
rect 4742 -5382 5510 -5348
rect 4680 -5617 4714 -5441
rect 5538 -5617 5572 -5441
rect 4742 -5710 5510 -5676
rect 5630 -5752 5672 -5306
rect 5672 -5752 5706 -5306
rect 5706 -5752 5750 -5306
rect 3714 -5910 3834 -5812
rect 2826 -5986 3594 -5952
rect 2764 -6221 2798 -6045
rect 3622 -6221 3656 -6045
rect 2826 -6314 3594 -6280
rect 3714 -6356 3756 -5910
rect 3756 -6356 3790 -5910
rect 3790 -6356 3834 -5910
rect 3714 -6486 3834 -6356
rect 4502 -5910 4622 -5812
rect 5630 -5848 5750 -5752
rect 4502 -6356 4546 -5910
rect 4546 -6356 4580 -5910
rect 4580 -6356 4622 -5910
rect 4742 -5986 5510 -5952
rect 4680 -6221 4714 -6045
rect 5538 -6221 5572 -6045
rect 4742 -6314 5510 -6280
rect 4502 -6486 4622 -6356
rect 5838 -6774 6324 -5156
rect 2510 -7181 3230 -7126
rect 2510 -7214 2513 -7181
rect 2513 -7214 2581 -7181
rect 2581 -7214 2671 -7181
rect 2671 -7214 2739 -7181
rect 2739 -7214 2829 -7181
rect 2829 -7214 2897 -7181
rect 2897 -7214 2987 -7181
rect 2987 -7214 3055 -7181
rect 3055 -7214 3145 -7181
rect 3145 -7214 3213 -7181
rect 3213 -7214 3230 -7181
rect 2420 -8041 2451 -7266
rect 2451 -8041 2485 -7266
rect 2485 -8041 2512 -7266
rect 2420 -8042 2512 -8041
rect 2578 -8041 2609 -7266
rect 2609 -8041 2643 -7266
rect 2643 -8041 2670 -7266
rect 2578 -8042 2670 -8041
rect 2736 -8041 2767 -7266
rect 2767 -8041 2801 -7266
rect 2801 -8041 2828 -7266
rect 2736 -8042 2828 -8041
rect 2894 -8041 2925 -7266
rect 2925 -8041 2959 -7266
rect 2959 -8041 2986 -7266
rect 2894 -8042 2986 -8041
rect 3050 -8041 3083 -7266
rect 3083 -8041 3117 -7266
rect 3117 -8041 3142 -7266
rect 3050 -8042 3142 -8041
rect 3210 -8041 3241 -7266
rect 3241 -8041 3275 -7266
rect 3275 -8041 3302 -7266
rect 3210 -8042 3302 -8041
rect 2512 -8125 2513 -8092
rect 2513 -8125 2581 -8092
rect 2581 -8125 2671 -8092
rect 2671 -8125 2739 -8092
rect 2739 -8125 2829 -8092
rect 2829 -8125 2897 -8092
rect 2897 -8125 2987 -8092
rect 2987 -8125 3055 -8092
rect 3055 -8125 3145 -8092
rect 3145 -8125 3212 -8092
rect 2512 -8172 3212 -8125
rect 3888 -7174 4588 -7120
rect 3888 -7208 3956 -7174
rect 3956 -7208 4046 -7174
rect 4046 -7208 4114 -7174
rect 4114 -7208 4204 -7174
rect 4204 -7208 4272 -7174
rect 4272 -7208 4362 -7174
rect 4362 -7208 4430 -7174
rect 4430 -7208 4520 -7174
rect 4520 -7208 4588 -7174
rect 3796 -7267 3888 -7266
rect 3796 -8043 3826 -7267
rect 3826 -8043 3860 -7267
rect 3860 -8043 3888 -7267
rect 3796 -8044 3888 -8043
rect 3954 -7267 4046 -7266
rect 3954 -8043 3984 -7267
rect 3984 -8043 4018 -7267
rect 4018 -8043 4046 -7267
rect 3954 -8044 4046 -8043
rect 4112 -7267 4204 -7266
rect 4112 -8043 4142 -7267
rect 4142 -8043 4176 -7267
rect 4176 -8043 4204 -7267
rect 4112 -8044 4204 -8043
rect 4270 -7267 4362 -7266
rect 4270 -8043 4300 -7267
rect 4300 -8043 4334 -7267
rect 4334 -8043 4362 -7267
rect 4270 -8044 4362 -8043
rect 4428 -7267 4520 -7266
rect 4428 -8043 4458 -7267
rect 4458 -8043 4492 -7267
rect 4492 -8043 4520 -7267
rect 4428 -8044 4520 -8043
rect 4586 -7267 4678 -7266
rect 4586 -8043 4616 -7267
rect 4616 -8043 4650 -7267
rect 4650 -8043 4678 -7267
rect 4586 -8044 4678 -8043
rect 3888 -8136 3956 -8102
rect 3956 -8136 4046 -8102
rect 4046 -8136 4114 -8102
rect 4114 -8136 4204 -8102
rect 4204 -8136 4272 -8102
rect 4272 -8136 4362 -8102
rect 4362 -8136 4430 -8102
rect 4430 -8136 4520 -8102
rect 4520 -8136 4588 -8102
rect 4588 -8136 4594 -8102
rect 3888 -8188 4594 -8136
rect 12462 -3416 12588 -3216
rect 12462 -3630 13646 -3416
rect 13950 -3460 14122 -3128
rect 15172 -3128 15940 -3094
rect 15110 -3254 15144 -3178
rect 15968 -3254 16002 -3178
rect 15172 -3338 15940 -3304
rect 16120 -3442 16212 -3004
rect 15034 -3516 16212 -3442
rect 8900 -4548 25134 -4316
rect 8900 -4734 11694 -4548
rect 8900 -4970 10462 -4734
rect 12058 -4748 16094 -4548
rect 16958 -4556 17330 -4548
rect 12058 -4750 15188 -4748
rect 15188 -4750 16094 -4748
rect 15282 -4844 16094 -4750
rect 10674 -4920 11042 -4886
rect 11252 -4920 11620 -4886
rect 11830 -4920 12198 -4886
rect 12408 -4920 12776 -4886
rect 12986 -4920 13354 -4886
rect 13564 -4920 13932 -4886
rect 14142 -4920 14510 -4886
rect 14720 -4920 15088 -4886
rect 8900 -5346 10478 -4970
rect 10478 -5346 10512 -4970
rect 10512 -5346 10612 -4970
rect 10612 -5346 10646 -4970
rect 10646 -5346 11070 -4970
rect 11070 -5346 11104 -4970
rect 11104 -5346 11190 -4970
rect 11190 -5346 11224 -4970
rect 8900 -5476 10462 -5346
rect 11452 -4970 11992 -4958
rect 11452 -5346 11648 -4970
rect 11648 -5346 11682 -4970
rect 11682 -5346 11768 -4970
rect 11768 -5346 11802 -4970
rect 11802 -5346 11992 -4970
rect 11452 -5354 11992 -5346
rect 12122 -5346 12226 -4970
rect 12226 -5346 12260 -4970
rect 12260 -5346 12346 -4970
rect 12346 -5346 12380 -4970
rect 12380 -5346 12488 -4970
rect 12604 -4970 12826 -4958
rect 12604 -5346 12804 -4970
rect 12804 -5346 12826 -4970
rect 12604 -5358 12826 -5346
rect 12924 -5346 12958 -4970
rect 12958 -5346 13168 -4970
rect 13276 -5346 13382 -4970
rect 13382 -5346 13416 -4970
rect 13416 -5346 13502 -4970
rect 13502 -5346 13536 -4970
rect 13536 -5346 13642 -4970
rect 13768 -4970 14308 -4958
rect 13768 -5346 13960 -4970
rect 13960 -5346 13994 -4970
rect 13994 -5346 14080 -4970
rect 14080 -5346 14114 -4970
rect 14114 -5346 14308 -4970
rect 13768 -5354 14308 -5346
rect 15282 -4970 15284 -4844
rect 14538 -5346 14572 -4970
rect 14572 -5346 14658 -4970
rect 14658 -5346 14692 -4970
rect 14692 -5346 15116 -4970
rect 15116 -5346 15150 -4970
rect 15150 -5346 15250 -4970
rect 15250 -5346 15284 -4970
rect 10674 -5430 11042 -5396
rect 11252 -5430 11620 -5396
rect 11830 -5430 12198 -5396
rect 12408 -5430 12776 -5396
rect 12986 -5430 13354 -5396
rect 13564 -5430 13932 -5396
rect 14142 -5430 14510 -5396
rect 14720 -5430 15088 -5396
rect 15282 -5472 15284 -5346
rect 15284 -5472 16094 -4844
rect 15282 -5530 16094 -5472
rect 15260 -5640 15938 -5636
rect 8878 -5758 15938 -5640
rect 16313 -4700 16607 -4666
rect 16771 -4700 17065 -4666
rect 17229 -4700 17523 -4666
rect 17687 -4700 17981 -4666
rect 18192 -4660 25134 -4548
rect 16666 -4750 16878 -4744
rect 16666 -4794 16672 -4750
rect 16228 -5484 16248 -4794
rect 16248 -5484 16672 -4794
rect 16666 -5526 16672 -5484
rect 16672 -5526 16706 -4750
rect 16706 -5526 16878 -4750
rect 16666 -5530 16878 -5526
rect 17044 -5526 17130 -4750
rect 17130 -5526 17164 -4750
rect 17164 -5526 17246 -4750
rect 17514 -5526 17588 -4750
rect 17588 -5526 17622 -4750
rect 17622 -5526 18046 -4750
rect 18046 -5526 18064 -4750
rect 16313 -5610 16607 -5576
rect 16771 -5610 17065 -5576
rect 17229 -5610 17523 -5576
rect 17687 -5610 17981 -5576
rect 18192 -5616 18194 -4660
rect 18194 -5218 25134 -4660
rect 18194 -5352 21246 -5218
rect 18194 -5456 18848 -5352
rect 18194 -5616 18788 -5456
rect 18192 -5674 18788 -5616
rect 18788 -5674 18822 -5456
rect 18822 -5548 18848 -5456
rect 18964 -5496 20532 -5462
rect 18808 -5712 18822 -5674
rect 18822 -5712 18862 -5548
rect 18902 -5622 18936 -5546
rect 20560 -5622 20594 -5546
rect 8878 -5776 16602 -5758
rect 8878 -6000 10492 -5776
rect 10735 -5942 11029 -5908
rect 11307 -5942 11601 -5908
rect 11879 -5942 12173 -5908
rect 12451 -5942 12745 -5908
rect 13023 -5942 13317 -5908
rect 13595 -5942 13889 -5908
rect 14167 -5942 14461 -5908
rect 14739 -5942 15033 -5908
rect 15260 -5878 16602 -5776
rect 16776 -5878 17510 -5762
rect 17700 -5864 18728 -5762
rect 18808 -5790 18862 -5712
rect 18964 -5706 20532 -5672
rect 20732 -5486 21246 -5352
rect 20732 -5776 21214 -5486
rect 22086 -5288 25134 -5218
rect 22086 -5298 23356 -5288
rect 23356 -5298 23662 -5288
rect 23662 -5298 25134 -5288
rect 21445 -5368 21579 -5334
rect 21703 -5368 21837 -5334
rect 21366 -5494 21400 -5418
rect 21624 -5494 21658 -5418
rect 21882 -5494 21916 -5418
rect 21445 -5578 21579 -5544
rect 21703 -5578 21837 -5544
rect 21366 -5704 21400 -5628
rect 21624 -5704 21658 -5628
rect 21882 -5704 21916 -5628
rect 21445 -5788 21579 -5754
rect 21703 -5788 21837 -5754
rect 17700 -5878 20504 -5864
rect 15260 -5888 16176 -5878
rect 16176 -5888 16602 -5878
rect 16776 -5888 17510 -5878
rect 17700 -5886 18118 -5878
rect 18118 -5886 20504 -5878
rect 8878 -6378 10522 -6000
rect 10522 -6378 10556 -6000
rect 10556 -6001 11242 -6000
rect 10556 -6377 10636 -6001
rect 10636 -6377 10670 -6001
rect 10670 -6377 11094 -6001
rect 11094 -6377 11128 -6001
rect 11128 -6377 11208 -6001
rect 11208 -6377 11242 -6001
rect 10556 -6378 11242 -6377
rect 8878 -6528 10492 -6378
rect 11602 -6001 11878 -6000
rect 11602 -6377 11666 -6001
rect 11666 -6377 11700 -6001
rect 11700 -6377 11780 -6001
rect 11780 -6377 11814 -6001
rect 11814 -6377 11878 -6001
rect 11602 -6378 11878 -6377
rect 12176 -6001 12452 -6000
rect 12176 -6377 12238 -6001
rect 12238 -6377 12272 -6001
rect 12272 -6377 12352 -6001
rect 12352 -6377 12386 -6001
rect 12386 -6377 12452 -6001
rect 12176 -6378 12452 -6377
rect 12924 -6001 13252 -5982
rect 12924 -6377 12958 -6001
rect 12958 -6377 13252 -6001
rect 12924 -6392 13252 -6377
rect 13316 -6001 13592 -6000
rect 13316 -6377 13382 -6001
rect 13382 -6377 13416 -6001
rect 13416 -6377 13496 -6001
rect 13496 -6377 13530 -6001
rect 13530 -6377 13592 -6001
rect 13316 -6378 13592 -6377
rect 13886 -6001 14162 -6000
rect 13886 -6377 13954 -6001
rect 13954 -6377 13988 -6001
rect 13988 -6377 14068 -6001
rect 14068 -6377 14102 -6001
rect 14102 -6377 14162 -6001
rect 13886 -6378 14162 -6377
rect 15260 -6000 15938 -5888
rect 14526 -6001 15212 -6000
rect 14526 -6377 14560 -6001
rect 14560 -6377 14640 -6001
rect 14640 -6377 14674 -6001
rect 14674 -6377 15098 -6001
rect 15098 -6377 15132 -6001
rect 15132 -6377 15212 -6001
rect 14526 -6378 15212 -6377
rect 15212 -6378 15246 -6000
rect 15246 -6378 15938 -6000
rect 10735 -6470 11029 -6436
rect 11307 -6470 11601 -6436
rect 11879 -6470 12173 -6436
rect 12451 -6470 12745 -6436
rect 13023 -6470 13317 -6436
rect 13595 -6470 13889 -6436
rect 14167 -6470 14461 -6436
rect 14739 -6470 15033 -6436
rect 8878 -6906 10522 -6528
rect 10522 -6906 10556 -6528
rect 10556 -6529 11242 -6528
rect 10556 -6905 10636 -6529
rect 10636 -6905 10670 -6529
rect 10670 -6905 11094 -6529
rect 11094 -6905 11128 -6529
rect 11128 -6905 11208 -6529
rect 11208 -6905 11242 -6529
rect 10556 -6906 11242 -6905
rect 8878 -7114 10492 -6906
rect 11602 -6529 11878 -6528
rect 11602 -6905 11666 -6529
rect 11666 -6905 11700 -6529
rect 11700 -6905 11780 -6529
rect 11780 -6905 11814 -6529
rect 11814 -6905 11878 -6529
rect 11602 -6906 11878 -6905
rect 12238 -6529 12388 -6528
rect 12174 -6905 12238 -6530
rect 12238 -6905 12272 -6529
rect 12272 -6905 12352 -6529
rect 12352 -6905 12386 -6529
rect 12386 -6530 12388 -6529
rect 12386 -6905 12450 -6530
rect 12174 -6908 12450 -6905
rect 12742 -6529 13018 -6528
rect 12742 -6905 12810 -6529
rect 12810 -6905 12844 -6529
rect 12844 -6905 12924 -6529
rect 12924 -6905 12958 -6529
rect 12958 -6905 13018 -6529
rect 12742 -6906 13018 -6905
rect 13316 -6529 13592 -6528
rect 13316 -6905 13382 -6529
rect 13382 -6905 13416 -6529
rect 13416 -6905 13496 -6529
rect 13496 -6905 13530 -6529
rect 13530 -6905 13592 -6529
rect 13316 -6906 13592 -6905
rect 13888 -6529 14164 -6528
rect 13888 -6905 13954 -6529
rect 13954 -6905 13988 -6529
rect 13988 -6905 14068 -6529
rect 14068 -6905 14102 -6529
rect 14102 -6905 14164 -6529
rect 13888 -6906 14164 -6905
rect 15260 -6528 15938 -6378
rect 14526 -6529 15212 -6528
rect 14526 -6905 14560 -6529
rect 14560 -6905 14640 -6529
rect 14640 -6905 14674 -6529
rect 14674 -6905 15098 -6529
rect 15098 -6905 15132 -6529
rect 15132 -6905 15212 -6529
rect 14526 -6906 15212 -6905
rect 15212 -6906 15246 -6528
rect 15246 -6906 15938 -6528
rect 10735 -6998 11029 -6964
rect 11307 -6998 11601 -6964
rect 11879 -6998 12173 -6964
rect 12451 -6998 12745 -6964
rect 13023 -6998 13317 -6964
rect 13595 -6998 13889 -6964
rect 14167 -6998 14461 -6964
rect 14739 -6998 15033 -6964
rect 15260 -7114 15938 -6906
rect 16162 -6016 16608 -5960
rect 16770 -6016 17066 -5956
rect 16162 -6050 16276 -6016
rect 16276 -6050 16608 -6016
rect 16770 -6050 17066 -6016
rect 17228 -6016 17524 -5956
rect 17686 -6016 18132 -5960
rect 17228 -6050 17524 -6016
rect 17686 -6050 18018 -6016
rect 18018 -6050 18132 -6016
rect 16224 -6109 16758 -6108
rect 16224 -6885 16248 -6109
rect 16248 -6885 16672 -6109
rect 16672 -6885 16706 -6109
rect 16706 -6885 16758 -6109
rect 16224 -6886 16758 -6885
rect 17014 -6109 17280 -6106
rect 17014 -6885 17130 -6109
rect 17130 -6885 17164 -6109
rect 17164 -6885 17280 -6109
rect 17014 -6890 17280 -6885
rect 17532 -6109 18066 -6108
rect 17532 -6885 17588 -6109
rect 17588 -6885 17622 -6109
rect 17622 -6885 18046 -6109
rect 18046 -6885 18066 -6109
rect 17532 -6886 18066 -6885
rect 16162 -6978 16276 -6944
rect 16276 -6978 16644 -6944
rect 16644 -6978 16734 -6944
rect 16734 -6978 17078 -6944
rect 16162 -7034 17078 -6978
rect 17216 -6978 17560 -6944
rect 17560 -6978 17650 -6944
rect 17650 -6978 18018 -6944
rect 18018 -6978 18132 -6944
rect 17216 -7034 18132 -6978
rect 18330 -6354 20504 -5886
rect 18330 -6460 18834 -6354
rect 18330 -6734 18768 -6460
rect 18768 -6734 18802 -6460
rect 18802 -6734 18834 -6460
rect 18944 -6500 20512 -6466
rect 18882 -6635 18916 -6559
rect 20540 -6635 20574 -6559
rect 18330 -6844 18834 -6734
rect 18944 -6728 20512 -6694
rect 20736 -6580 21184 -5870
rect 22086 -5384 23274 -5298
rect 22086 -5406 23260 -5384
rect 23260 -5406 23274 -5384
rect 22086 -5758 22816 -5406
rect 23446 -5436 23572 -5402
rect 23362 -5632 23396 -5464
rect 23622 -5632 23656 -5464
rect 23446 -5694 23572 -5660
rect 22086 -5852 22638 -5758
rect 23778 -5834 25134 -5298
rect 22398 -6224 22620 -5948
rect 20736 -6844 21202 -6580
rect 21445 -6364 21579 -6330
rect 21703 -6364 21837 -6330
rect 21366 -6499 21400 -6423
rect 21624 -6499 21658 -6423
rect 21882 -6499 21916 -6423
rect 21445 -6592 21579 -6558
rect 21703 -6592 21837 -6558
rect 21366 -6727 21400 -6651
rect 21624 -6727 21658 -6651
rect 21882 -6727 21916 -6651
rect 21445 -6820 21579 -6786
rect 21703 -6820 21837 -6786
rect 18330 -6930 21202 -6844
rect 22118 -6694 22620 -6224
rect 24312 -6246 25178 -5946
rect 22118 -6802 22930 -6694
rect 23143 -6438 23919 -6404
rect 23050 -6634 23084 -6466
rect 23978 -6634 24012 -6466
rect 23143 -6696 23919 -6662
rect 24114 -6802 25178 -6246
rect 22118 -6810 23044 -6802
rect 23044 -6810 24018 -6802
rect 24018 -6810 25180 -6802
rect 22118 -6930 25180 -6810
rect 18330 -7114 25180 -6930
rect 8878 -7116 16176 -7114
rect 16176 -7116 18118 -7114
rect 18118 -7116 25180 -7114
rect 8878 -7248 25180 -7116
rect 8878 -7250 21202 -7248
rect 8878 -7320 10008 -7250
rect 8878 -7354 9710 -7320
rect 9710 -7354 9984 -7320
rect 9984 -7354 10008 -7320
rect 8878 -7366 10008 -7354
rect 8940 -7682 9046 -7608
rect 8940 -9410 9034 -7682
rect 9034 -9410 9046 -7682
rect 9220 -7734 9296 -7700
rect 9136 -9330 9170 -7762
rect 9208 -9240 9304 -7774
rect 9346 -9330 9380 -7762
rect 8940 -9442 9046 -9410
rect 9220 -9392 9296 -9358
rect 9809 -7468 9885 -7434
rect 9716 -9064 9750 -7496
rect 9788 -9050 9904 -7570
rect 9944 -9064 9978 -7496
rect 9809 -9126 9885 -9092
rect 10162 -9408 10362 -9088
rect 9466 -9410 9482 -9408
rect 9482 -9410 10362 -9408
rect 9466 -9442 10362 -9410
rect 8940 -9472 10362 -9442
rect 8940 -9506 9130 -9472
rect 9130 -9506 9386 -9472
rect 9386 -9506 10362 -9472
rect 8940 -9960 10362 -9506
rect 10638 -7492 11035 -7454
rect 24237 -7492 24634 -7454
rect 10638 -7658 11035 -7620
rect 24237 -7658 24634 -7620
rect 10638 -7824 11035 -7786
rect 24237 -7824 24634 -7786
rect 10638 -7990 11035 -7952
rect 24237 -7990 24634 -7952
rect 10638 -8156 11035 -8118
rect 24237 -8156 24634 -8118
rect 10638 -8322 11035 -8284
rect 24237 -8322 24634 -8284
rect 10638 -8488 11035 -8450
rect 24237 -8488 24634 -8450
rect 10638 -8654 11035 -8616
rect 24237 -8654 24634 -8616
rect 10638 -8820 11035 -8782
rect 24237 -8820 24634 -8782
rect 10638 -8986 11035 -8948
rect 24237 -8986 24634 -8948
rect 10638 -9152 11035 -9114
rect 24237 -9152 24634 -9114
rect 10638 -9318 11035 -9280
rect 24237 -9318 24634 -9280
rect 10638 -9484 11035 -9446
rect 24237 -9484 24634 -9446
rect 10638 -9650 11035 -9612
rect 24237 -9650 24634 -9612
rect 10638 -9816 11035 -9778
rect 24237 -9816 24634 -9778
rect 24788 -9960 25116 -7404
rect 8940 -9962 10586 -9960
rect 10586 -9962 24686 -9960
rect 24686 -9962 25116 -9960
rect 8940 -10142 25116 -9962
rect 1996 -12792 7070 -11824
rect 7814 -12034 21870 -11798
rect 7342 -12212 7510 -12178
rect 7280 -12438 7314 -12262
rect 7538 -12438 7572 -12262
rect 7342 -12522 7510 -12488
rect 13436 -12194 21870 -12034
rect 8284 -12272 9852 -12238
rect 9942 -12272 11510 -12238
rect 11600 -12272 13168 -12238
rect 8222 -12382 8256 -12322
rect 8348 -12382 9840 -12322
rect 9880 -12382 9914 -12322
rect 11538 -12382 11572 -12322
rect 13196 -12382 13230 -12322
rect 8284 -12466 9852 -12432
rect 9942 -12466 11510 -12432
rect 11600 -12466 13168 -12432
rect 13436 -12566 20150 -12510
rect 20656 -12566 21870 -12194
rect 22152 -11672 25426 -11668
rect 22152 -12538 25428 -11672
rect 13436 -12600 19884 -12566
rect 19884 -12600 20150 -12566
rect 20656 -12600 21822 -12566
rect 21822 -12600 21870 -12566
rect 13436 -12662 20150 -12600
rect 20656 -12646 21870 -12600
rect 13436 -12680 19788 -12662
rect 7778 -12792 19788 -12680
rect 19788 -12752 19822 -12662
rect 19822 -12700 20150 -12662
rect 19822 -12734 20010 -12700
rect 20010 -12734 20150 -12700
rect 19822 -12752 20150 -12734
rect 1996 -12826 3100 -12792
rect 3100 -12826 7070 -12792
rect 7778 -12826 19000 -12792
rect 19000 -12826 19788 -12792
rect 1996 -12862 7070 -12826
rect 1996 -13538 2982 -12862
rect 7778 -12888 19788 -12826
rect 7778 -12898 19062 -12888
rect 19062 -12898 19096 -12888
rect 3152 -12976 3549 -12938
rect 18551 -12976 18948 -12938
rect 3152 -13142 3549 -13104
rect 18551 -13142 18948 -13104
rect 19070 -13098 19096 -12898
rect 19096 -13098 19788 -12888
rect 19788 -13098 19808 -12752
rect 3152 -13308 3549 -13270
rect 18551 -13308 18948 -13270
rect 3152 -13474 3549 -13436
rect 18551 -13474 18948 -13436
rect 1996 -13586 19328 -13538
rect 1996 -13620 3100 -13586
rect 3100 -13620 19000 -13586
rect 19000 -13620 19328 -13586
rect 1996 -13730 19328 -13620
rect 1996 -13764 2098 -13730
rect 2098 -13764 19328 -13730
rect 1996 -13814 19328 -13764
rect 2150 -13914 2547 -13876
rect 18949 -13914 19346 -13876
rect 2150 -14080 2547 -14042
rect 18949 -14080 19346 -14042
rect 2150 -14246 2547 -14208
rect 18949 -14246 19346 -14208
rect 2150 -14412 2547 -14374
rect 18949 -14412 19346 -14374
rect 2150 -14578 2547 -14540
rect 18949 -14578 19346 -14540
rect 2150 -14744 2547 -14706
rect 18949 -14744 19346 -14706
rect 2150 -14910 2547 -14872
rect 18949 -14910 19346 -14872
rect 2150 -15076 2547 -15038
rect 18949 -15076 19346 -15038
rect 2150 -15242 2547 -15204
rect 18949 -15242 19346 -15204
rect 2150 -15408 2547 -15370
rect 18949 -15408 19346 -15370
rect 2150 -15574 2547 -15536
rect 18949 -15574 19346 -15536
rect 2150 -15740 2547 -15702
rect 18949 -15740 19346 -15702
rect 2150 -15906 2547 -15868
rect 18949 -15906 19346 -15868
rect 2150 -16072 2547 -16034
rect 18949 -16072 19346 -16034
rect 2150 -16238 2547 -16200
rect 18949 -16238 19346 -16200
rect 2150 -16404 2547 -16366
rect 18949 -16404 19346 -16366
rect 2150 -16570 2547 -16532
rect 18949 -16570 19346 -16532
rect 2150 -16736 2547 -16698
rect 18949 -16736 19346 -16698
rect 2150 -16902 2547 -16864
rect 18949 -16902 19346 -16864
rect 2150 -17068 2547 -17030
rect 18949 -17068 19346 -17030
rect 2150 -17234 2547 -17196
rect 18949 -17234 19346 -17196
rect 2150 -17400 2547 -17362
rect 18949 -17400 19346 -17362
rect 2150 -17566 2547 -17528
rect 18949 -17566 19346 -17528
rect 2150 -17732 2547 -17694
rect 18949 -17732 19346 -17694
rect 2150 -17898 2547 -17860
rect 18949 -17898 19346 -17860
rect 2150 -18064 2547 -18026
rect 18949 -18064 19346 -18026
rect 19926 -13093 19960 -12799
rect 20836 -13093 20870 -12799
rect 21746 -13093 21780 -12799
rect 20008 -13278 20788 -13244
rect 20008 -13312 20010 -13278
rect 20010 -13312 20786 -13278
rect 20786 -13312 20788 -13278
rect 20918 -13278 21698 -13242
rect 20008 -13352 20788 -13312
rect 19926 -13671 19960 -13377
rect 20918 -13312 20920 -13278
rect 20920 -13312 21696 -13278
rect 21696 -13312 21698 -13278
rect 20918 -13350 21698 -13312
rect 19998 -13600 20798 -13452
rect 20836 -13671 20870 -13377
rect 20908 -13600 21708 -13452
rect 20010 -13736 20786 -13702
rect 20010 -13770 20786 -13736
rect 21746 -13671 21780 -13377
rect 20920 -13736 21696 -13700
rect 20010 -13856 20786 -13770
rect 20920 -13770 21696 -13736
rect 20920 -13800 21696 -13770
rect 20010 -13870 20786 -13856
rect 20204 -13890 20622 -13870
rect 19926 -14249 19960 -13955
rect 20204 -14314 20622 -13890
rect 20836 -14249 20870 -13955
rect 20920 -13890 21696 -13856
rect 20920 -13952 21696 -13890
rect 21828 -13874 21884 -13758
rect 21884 -13874 21918 -13758
rect 21918 -13874 21944 -13758
rect 20916 -14308 21698 -14052
rect 21746 -14249 21780 -13955
rect 20204 -14336 20622 -14314
rect 20010 -14348 20786 -14336
rect 20010 -14434 20786 -14348
rect 20010 -14468 20786 -14434
rect 20920 -14434 21696 -14404
rect 20010 -14500 20786 -14468
rect 19926 -14827 19960 -14533
rect 20920 -14468 21696 -14434
rect 20920 -14504 21696 -14468
rect 19998 -14750 20798 -14602
rect 20836 -14827 20870 -14533
rect 20908 -14748 21708 -14600
rect 20008 -14892 20788 -14854
rect 20008 -14926 20010 -14892
rect 20010 -14926 20786 -14892
rect 20786 -14926 20788 -14892
rect 21746 -14827 21780 -14533
rect 20920 -14892 21700 -14854
rect 20008 -14962 20788 -14926
rect 20920 -14926 21696 -14892
rect 21696 -14926 21700 -14892
rect 20920 -14962 21700 -14926
rect 19926 -15405 19960 -15111
rect 20836 -15405 20870 -15111
rect 21746 -15405 21780 -15111
rect 19534 -15604 21862 -15548
rect 19534 -15638 19884 -15604
rect 19884 -15638 21822 -15604
rect 21822 -15638 21862 -15604
rect 19534 -15878 21862 -15638
rect 19534 -16020 20220 -15878
rect 19534 -17992 20222 -16020
rect 19534 -18128 20220 -17992
rect 20474 -16044 21252 -16008
rect 20474 -16078 20476 -16044
rect 20476 -16078 21252 -16044
rect 20392 -16174 20426 -16106
rect 20474 -16202 21252 -16078
rect 21302 -16174 21336 -16106
rect 20474 -16236 20476 -16202
rect 20476 -16236 21252 -16202
rect 20392 -16332 20426 -16264
rect 20474 -16268 21252 -16236
rect 20476 -16360 21252 -16332
rect 21302 -16332 21336 -16264
rect 20476 -16394 21252 -16360
rect 20392 -16490 20426 -16422
rect 20476 -16424 21252 -16394
rect 20476 -16518 21252 -16490
rect 21302 -16490 21336 -16422
rect 20476 -16552 21252 -16518
rect 20392 -16648 20426 -16580
rect 20476 -16582 21252 -16552
rect 20476 -16676 21252 -16648
rect 21302 -16648 21336 -16580
rect 20476 -16710 21252 -16676
rect 20392 -16806 20426 -16738
rect 20476 -16740 21252 -16710
rect 20476 -16834 21252 -16806
rect 21302 -16806 21336 -16738
rect 20476 -16868 21252 -16834
rect 20392 -16964 20426 -16896
rect 20476 -16898 21252 -16868
rect 20476 -16992 21252 -16964
rect 21302 -16964 21336 -16896
rect 20476 -17026 21252 -16992
rect 20392 -17122 20426 -17054
rect 20476 -17056 21252 -17026
rect 20476 -17150 21252 -17122
rect 21302 -17122 21336 -17054
rect 20476 -17184 21252 -17150
rect 20392 -17280 20426 -17212
rect 20476 -17214 21252 -17184
rect 20476 -17308 21252 -17280
rect 21302 -17280 21336 -17212
rect 20476 -17342 21252 -17308
rect 20392 -17438 20426 -17370
rect 20476 -17372 21252 -17342
rect 20476 -17466 21252 -17438
rect 21302 -17438 21336 -17370
rect 20476 -17500 21252 -17466
rect 20392 -17596 20426 -17528
rect 20476 -17530 21252 -17500
rect 20476 -17624 21252 -17596
rect 21302 -17596 21336 -17528
rect 20476 -17658 21252 -17624
rect 20392 -17754 20426 -17686
rect 20476 -17688 21252 -17658
rect 20472 -17782 21252 -17756
rect 21302 -17754 21336 -17686
rect 20472 -17816 20476 -17782
rect 20476 -17816 21252 -17782
rect 20392 -17912 20426 -17844
rect 20472 -17940 21252 -17816
rect 21302 -17912 21336 -17844
rect 20472 -17974 20476 -17940
rect 20476 -17974 21252 -17940
rect 20472 -17996 21252 -17974
rect 20474 -18010 21252 -17996
rect 21532 -16254 21862 -15878
rect 22520 -13101 22554 -12807
rect 22520 -13679 22554 -13385
rect 22608 -13138 23388 -13092
rect 22608 -13166 23390 -13138
rect 23448 -13101 23482 -12807
rect 22608 -13200 22613 -13166
rect 22613 -13200 23389 -13166
rect 23389 -13200 23390 -13166
rect 22608 -13286 23390 -13200
rect 22608 -13320 22613 -13286
rect 22613 -13320 23389 -13286
rect 23389 -13320 23390 -13286
rect 22608 -13344 23390 -13320
rect 22608 -13392 23388 -13344
rect 22520 -14257 22554 -13963
rect 22610 -13744 23390 -13668
rect 23448 -13679 23482 -13385
rect 23538 -13166 24318 -13090
rect 24376 -13101 24410 -12807
rect 23538 -13200 23541 -13166
rect 23541 -13200 24317 -13166
rect 24317 -13200 24318 -13166
rect 23538 -13286 24318 -13200
rect 23538 -13320 23541 -13286
rect 23541 -13320 24317 -13286
rect 24317 -13320 24318 -13286
rect 23538 -13390 24318 -13320
rect 22610 -13778 22613 -13744
rect 22613 -13778 23389 -13744
rect 23389 -13778 23390 -13744
rect 22610 -13864 23390 -13778
rect 22610 -13898 22613 -13864
rect 22613 -13898 23389 -13864
rect 23389 -13898 23390 -13864
rect 22610 -13968 23390 -13898
rect 22520 -14835 22554 -14541
rect 22608 -14298 23388 -14242
rect 22608 -14322 23390 -14298
rect 23448 -14257 23482 -13963
rect 23536 -13716 24316 -13666
rect 24376 -13679 24410 -13385
rect 23536 -13744 24318 -13716
rect 23536 -13778 23541 -13744
rect 23541 -13778 24317 -13744
rect 24317 -13778 24318 -13744
rect 23536 -13864 24318 -13778
rect 23536 -13898 23541 -13864
rect 23541 -13898 24317 -13864
rect 24317 -13898 24318 -13864
rect 23536 -13922 24318 -13898
rect 23536 -13966 24316 -13922
rect 22608 -14356 22613 -14322
rect 22613 -14356 23389 -14322
rect 23389 -14356 23390 -14322
rect 22608 -14442 23390 -14356
rect 22608 -14476 22613 -14442
rect 22613 -14476 23389 -14442
rect 23389 -14476 23390 -14442
rect 22608 -14504 23390 -14476
rect 22608 -14542 23388 -14504
rect 22610 -14900 23390 -14814
rect 23448 -14835 23482 -14541
rect 23538 -14322 24318 -14238
rect 24376 -14257 24410 -13963
rect 23538 -14356 23541 -14322
rect 23541 -14356 24317 -14322
rect 24317 -14356 24318 -14322
rect 23538 -14442 24318 -14356
rect 23538 -14476 23541 -14442
rect 23541 -14476 24317 -14442
rect 24317 -14476 24318 -14442
rect 23538 -14538 24318 -14476
rect 22610 -14934 22613 -14900
rect 22613 -14934 23389 -14900
rect 23389 -14934 23390 -14900
rect 22610 -14976 23390 -14934
rect 22520 -15413 22554 -15119
rect 24376 -14835 24410 -14541
rect 23448 -15413 23482 -15119
rect 22612 -15632 22613 -15598
rect 22613 -15632 23389 -15598
rect 23389 -15632 23390 -15598
rect 22612 -15642 23390 -15632
rect 23570 -14934 24284 -14908
rect 23570 -15020 24284 -14934
rect 23570 -15054 24284 -15020
rect 23570 -15478 24284 -15054
rect 24376 -15413 24410 -15119
rect 23570 -15512 24284 -15478
rect 23570 -15598 24284 -15512
rect 23570 -15622 24284 -15598
rect 22520 -15991 22554 -15697
rect 22610 -15914 23392 -15642
rect 22520 -16569 22554 -16275
rect 22610 -16056 23390 -15988
rect 23448 -15991 23482 -15697
rect 22610 -16090 22613 -16056
rect 22613 -16090 23389 -16056
rect 23389 -16090 23390 -16056
rect 22610 -16176 23390 -16090
rect 22610 -16210 22613 -16176
rect 22613 -16210 23389 -16176
rect 23389 -16210 23390 -16176
rect 22610 -16288 23390 -16210
rect 22520 -17147 22554 -16853
rect 22610 -16634 23390 -16552
rect 23448 -16569 23482 -16275
rect 23538 -16056 24318 -15988
rect 24376 -15991 24410 -15697
rect 23538 -16090 23541 -16056
rect 23541 -16090 24317 -16056
rect 24317 -16090 24318 -16056
rect 23538 -16176 24318 -16090
rect 23538 -16210 23541 -16176
rect 23541 -16210 24317 -16176
rect 24317 -16210 24318 -16176
rect 23538 -16288 24318 -16210
rect 22610 -16668 22613 -16634
rect 22613 -16668 23389 -16634
rect 23389 -16668 23390 -16634
rect 22610 -16754 23390 -16668
rect 22610 -16788 22613 -16754
rect 22613 -16788 23389 -16754
rect 23389 -16788 23390 -16754
rect 22610 -16852 23390 -16788
rect 22520 -17725 22554 -17431
rect 22610 -17212 23390 -17138
rect 23448 -17147 23482 -16853
rect 23536 -16606 24316 -16552
rect 23536 -16634 24318 -16606
rect 24376 -16569 24410 -16275
rect 23536 -16668 23541 -16634
rect 23541 -16668 24317 -16634
rect 24317 -16668 24318 -16634
rect 23536 -16754 24318 -16668
rect 23536 -16788 23541 -16754
rect 23541 -16788 24317 -16754
rect 24317 -16788 24318 -16754
rect 23536 -16812 24318 -16788
rect 23536 -16852 24316 -16812
rect 22610 -17246 22613 -17212
rect 22613 -17246 23389 -17212
rect 23389 -17246 23390 -17212
rect 22610 -17332 23390 -17246
rect 22610 -17366 22613 -17332
rect 22613 -17366 23389 -17332
rect 23389 -17366 23390 -17332
rect 22610 -17438 23390 -17366
rect 23448 -17725 23482 -17431
rect 23538 -17212 24318 -17136
rect 24376 -17147 24410 -16853
rect 23538 -17246 23541 -17212
rect 23541 -17246 24317 -17212
rect 24317 -17246 24318 -17212
rect 23538 -17332 24318 -17246
rect 23538 -17366 23541 -17332
rect 23541 -17366 24317 -17332
rect 24317 -17366 24318 -17332
rect 23538 -17436 24318 -17366
rect 24376 -17725 24410 -17431
rect 24616 -17924 25428 -12538
rect 1996 -18176 18346 -18128
rect 18856 -18176 20220 -18128
rect 1996 -18210 2098 -18176
rect 2098 -18210 18346 -18176
rect 18856 -18210 19398 -18176
rect 19398 -18210 20220 -18176
rect 1996 -18320 18346 -18210
rect 18856 -18320 20220 -18210
rect 1996 -18354 2096 -18320
rect 2096 -18354 18346 -18320
rect 18856 -18354 20220 -18320
rect 1996 -18408 18346 -18354
rect 18856 -18408 20220 -18354
rect 19534 -18466 20220 -18408
rect 2148 -18504 2545 -18466
rect 24547 -18504 24944 -18466
rect 2148 -18670 2545 -18632
rect 24547 -18670 24944 -18632
rect 2148 -18836 2545 -18798
rect 24547 -18836 24944 -18798
rect 2148 -19002 2545 -18964
rect 24547 -19002 24944 -18964
rect 2148 -19168 2545 -19130
rect 24547 -19168 24944 -19130
rect 2148 -19334 2545 -19296
rect 24547 -19334 24944 -19296
rect 2148 -19500 2545 -19462
rect 24547 -19500 24944 -19462
rect 2148 -19666 2545 -19628
rect 24547 -19666 24944 -19628
rect 2148 -19832 2545 -19794
rect 24547 -19832 24944 -19794
rect 2148 -19998 2545 -19960
rect 24547 -19998 24944 -19960
rect 2148 -20164 2545 -20126
rect 24547 -20164 24944 -20126
rect 2148 -20330 2545 -20292
rect 24547 -20330 24944 -20292
rect 2148 -20496 2545 -20458
rect 24547 -20496 24944 -20458
rect 2148 -20662 2545 -20624
rect 24547 -20662 24944 -20624
rect 2148 -20828 2545 -20790
rect 24547 -20828 24944 -20790
rect 2148 -20994 2545 -20956
rect 24547 -20994 24944 -20956
rect 2148 -21160 2545 -21122
rect 24547 -21160 24944 -21122
rect 2148 -21326 2545 -21288
rect 24547 -21326 24944 -21288
rect 2148 -21492 2545 -21454
rect 24547 -21492 24944 -21454
rect 2148 -21658 2545 -21620
rect 24547 -21658 24944 -21620
rect 2148 -21824 2545 -21786
rect 24547 -21824 24944 -21786
rect 2148 -21990 2545 -21952
rect 24547 -21990 24944 -21952
rect 2148 -22156 2545 -22118
rect 24547 -22156 24944 -22118
rect 2148 -22322 2545 -22284
rect 24547 -22322 24944 -22284
rect 2148 -22488 2545 -22450
rect 24547 -22488 24944 -22450
rect 1890 -23440 20268 -22710
rect 20472 -23018 20538 -22952
rect 21482 -22924 21544 -22828
rect 21328 -23008 21394 -22942
rect 21482 -23026 21508 -22924
rect 21508 -23026 21544 -22924
rect 21482 -23096 21544 -23026
rect 21226 -23122 21310 -23096
rect 21310 -23122 21412 -23096
rect 21412 -23122 21544 -23096
rect 21226 -23158 21544 -23122
rect 21764 -23598 22366 -23090
rect 22604 -22926 22666 -22830
rect 22604 -23028 22640 -22926
rect 22640 -23028 22666 -22926
rect 22754 -23010 22820 -22944
rect 22604 -23098 22666 -23028
rect 22604 -23124 22736 -23098
rect 22736 -23124 22838 -23098
rect 22838 -23124 22922 -23098
rect 22604 -23160 22922 -23124
rect 23580 -23020 23646 -22954
rect 24070 -23568 25410 -22730
<< metal1 >>
rect 1626 -826 2026 -812
rect 1626 -1200 1638 -826
rect 2012 -1200 2026 -826
rect 1626 -1212 2026 -1200
rect 2178 -826 2578 -812
rect 2178 -1200 2190 -826
rect 2564 -1200 2578 -826
rect 3592 -826 3992 -812
rect 2178 -1212 2578 -1200
rect 2676 -864 2820 -850
rect 2676 -1182 2748 -864
rect 2806 -1110 2820 -864
rect 3592 -946 3606 -826
rect 2882 -956 3606 -946
rect 2882 -964 3156 -956
rect 2882 -1030 2900 -964
rect 2966 -1030 3156 -964
rect 2882 -1046 3156 -1030
rect 2806 -1128 3046 -1110
rect 3018 -1182 3046 -1128
rect 2676 -1236 3046 -1182
rect 3146 -1180 3156 -1046
rect 3236 -1046 3606 -956
rect 3236 -1180 3246 -1046
rect 3146 -1194 3246 -1180
rect 3592 -1200 3606 -1046
rect 3980 -1200 3992 -826
rect 3592 -1212 3992 -1200
rect 4338 -824 4738 -812
rect 4338 -1198 4350 -824
rect 4724 -948 4738 -824
rect 8076 -822 8476 -812
rect 5516 -852 6032 -850
rect 5516 -884 6112 -852
rect 4724 -958 5454 -948
rect 4724 -1048 5096 -958
rect 4724 -1198 4738 -1048
rect 5086 -1180 5096 -1048
rect 5176 -964 5454 -958
rect 5176 -1030 5370 -964
rect 5436 -1030 5454 -964
rect 5176 -1048 5454 -1030
rect 5176 -1180 5186 -1048
rect 5516 -1110 5530 -884
rect 5086 -1192 5186 -1180
rect 5290 -1126 5530 -1110
rect 5290 -1180 5316 -1126
rect 5586 -1180 6112 -884
rect 4338 -1212 4738 -1198
rect 2676 -1261 2998 -1236
rect 2676 -1295 2933 -1261
rect 2967 -1295 2998 -1261
rect 2676 -1353 2998 -1295
rect 2676 -1354 2933 -1353
rect 2084 -1387 2933 -1354
rect 2967 -1387 2998 -1353
rect 2084 -1445 2998 -1387
rect 2084 -1479 2933 -1445
rect 2967 -1479 2998 -1445
rect 2084 -1537 2998 -1479
rect 2084 -1571 2933 -1537
rect 2967 -1571 2998 -1537
rect 2084 -1600 2998 -1571
rect 3446 -1261 3542 -1232
rect 3446 -1295 3477 -1261
rect 3511 -1286 3542 -1261
rect 4788 -1261 4884 -1232
rect 5290 -1236 6112 -1180
rect 8076 -1200 8088 -822
rect 8464 -1200 8476 -822
rect 8076 -1212 8476 -1200
rect 9976 -818 10376 -812
rect 9976 -1206 9982 -818
rect 10370 -1206 10376 -818
rect 9976 -1212 10376 -1206
rect 11192 -822 11592 -812
rect 11192 -1204 11200 -822
rect 11580 -1204 11592 -822
rect 23912 -820 24312 -812
rect 22388 -842 23808 -840
rect 14212 -846 23808 -842
rect 11192 -1212 11592 -1204
rect 12558 -960 23808 -846
rect 4788 -1286 4819 -1261
rect 3511 -1295 4819 -1286
rect 4853 -1295 4884 -1261
rect 3446 -1353 4884 -1295
rect 3446 -1387 3477 -1353
rect 3511 -1387 4819 -1353
rect 4853 -1387 4884 -1353
rect 3446 -1445 4884 -1387
rect 3446 -1479 3477 -1445
rect 3511 -1479 4819 -1445
rect 4853 -1479 4884 -1445
rect 3446 -1537 4884 -1479
rect 3446 -1571 3477 -1537
rect 3511 -1571 4819 -1537
rect 4853 -1571 4884 -1537
rect 3446 -1600 4884 -1571
rect 5332 -1261 6112 -1236
rect 5332 -1295 5363 -1261
rect 5397 -1295 6112 -1261
rect 5332 -1353 6112 -1295
rect 7372 -1344 7472 -1338
rect 5332 -1387 5363 -1353
rect 5397 -1387 6112 -1353
rect 5332 -1445 6112 -1387
rect 7234 -1444 7372 -1344
rect 7472 -1444 12358 -1344
rect 12458 -1444 12464 -1344
rect 5332 -1479 5363 -1445
rect 5397 -1479 6112 -1445
rect 5332 -1537 6112 -1479
rect 5332 -1571 5363 -1537
rect 5397 -1571 6112 -1537
rect 5332 -1600 6112 -1571
rect 2084 -1856 2756 -1600
rect 3038 -1690 3426 -1680
rect 3038 -1772 3046 -1690
rect 3414 -1772 3426 -1690
rect 3038 -1780 3426 -1772
rect 3038 -1842 3278 -1780
rect 2084 -1948 2754 -1856
rect 2084 -2496 2652 -1948
rect 2748 -1982 2754 -1948
rect 2686 -1994 2754 -1982
rect 2686 -2148 2698 -1994
rect 2894 -2010 3278 -1842
rect 3518 -1864 4838 -1600
rect 4904 -1682 5292 -1672
rect 4904 -1764 4912 -1682
rect 5280 -1764 5292 -1682
rect 4904 -1772 5292 -1764
rect 3670 -1866 4838 -1864
rect 5058 -1842 5292 -1772
rect 3670 -1940 4666 -1866
rect 3670 -1974 3676 -1940
rect 3670 -1986 3738 -1974
rect 2862 -2036 3562 -2010
rect 2862 -2042 3608 -2036
rect 2862 -2044 3428 -2042
rect 2816 -2050 3428 -2044
rect 2816 -2084 2828 -2050
rect 2996 -2076 3428 -2050
rect 3596 -2076 3608 -2042
rect 2996 -2082 3608 -2076
rect 2996 -2084 3562 -2082
rect 2816 -2090 3562 -2084
rect 2758 -2134 2806 -2122
rect 2758 -2148 2766 -2134
rect 2686 -2294 2766 -2148
rect 2686 -2450 2698 -2294
rect 2758 -2310 2766 -2294
rect 2800 -2310 2806 -2134
rect 2758 -2322 2806 -2310
rect 2862 -2354 2962 -2090
rect 3018 -2134 3064 -2122
rect 3018 -2310 3024 -2134
rect 3058 -2172 3064 -2134
rect 3360 -2135 3406 -2123
rect 3360 -2172 3366 -2135
rect 3058 -2272 3366 -2172
rect 3058 -2310 3064 -2272
rect 3018 -2322 3064 -2310
rect 3162 -2350 3262 -2272
rect 3360 -2311 3366 -2272
rect 3400 -2311 3406 -2135
rect 3360 -2323 3406 -2311
rect 2816 -2360 3008 -2354
rect 2816 -2394 2828 -2360
rect 2996 -2394 3008 -2360
rect 2816 -2400 3008 -2394
rect 2686 -2462 2754 -2450
rect 2748 -2476 2754 -2462
rect 2748 -2496 3056 -2476
rect 2084 -2854 3056 -2496
rect 3162 -2656 3168 -2350
rect 3256 -2656 3262 -2350
rect 3462 -2364 3562 -2090
rect 3624 -2123 3664 -2122
rect 3618 -2135 3664 -2123
rect 3618 -2311 3624 -2135
rect 3658 -2150 3664 -2135
rect 3724 -2150 3738 -1986
rect 3658 -2296 3738 -2150
rect 3658 -2311 3664 -2296
rect 3618 -2323 3664 -2311
rect 3624 -2324 3664 -2323
rect 3416 -2370 3608 -2364
rect 3416 -2404 3428 -2370
rect 3596 -2404 3608 -2370
rect 3416 -2410 3468 -2404
rect 3162 -2662 3262 -2656
rect 3462 -2654 3468 -2410
rect 3556 -2410 3608 -2404
rect 3556 -2654 3562 -2410
rect 3724 -2460 3738 -2296
rect 3670 -2472 3738 -2460
rect 3772 -2044 4564 -1940
rect 4660 -1974 4666 -1940
rect 3670 -2488 3676 -2472
rect 3462 -2662 3562 -2654
rect 3632 -2506 3676 -2488
rect 3772 -2506 3788 -2044
rect 3632 -2726 3788 -2506
rect 4544 -2506 4564 -2044
rect 4598 -1986 4666 -1974
rect 4598 -2150 4612 -1986
rect 5058 -2010 5442 -1842
rect 5578 -1846 6112 -1600
rect 5582 -1948 6112 -1846
rect 5582 -1982 5588 -1948
rect 5582 -1994 5650 -1982
rect 4774 -2036 5474 -2010
rect 4728 -2042 5474 -2036
rect 4728 -2076 4740 -2042
rect 4908 -2044 5474 -2042
rect 4908 -2050 5520 -2044
rect 4908 -2076 5340 -2050
rect 4728 -2082 5340 -2076
rect 4774 -2084 5340 -2082
rect 5508 -2084 5520 -2050
rect 4774 -2090 5520 -2084
rect 4672 -2123 4712 -2122
rect 4672 -2135 4718 -2123
rect 4672 -2150 4678 -2135
rect 4598 -2296 4678 -2150
rect 4598 -2460 4612 -2296
rect 4672 -2311 4678 -2296
rect 4712 -2311 4718 -2135
rect 4672 -2323 4718 -2311
rect 4672 -2324 4712 -2323
rect 4774 -2364 4874 -2090
rect 4930 -2135 4976 -2123
rect 4930 -2311 4936 -2135
rect 4970 -2172 4976 -2135
rect 5272 -2134 5318 -2122
rect 5272 -2172 5278 -2134
rect 4970 -2272 5278 -2172
rect 4970 -2311 4976 -2272
rect 4930 -2323 4976 -2311
rect 5074 -2350 5174 -2272
rect 5272 -2310 5278 -2272
rect 5312 -2310 5318 -2134
rect 5272 -2322 5318 -2310
rect 4728 -2370 4920 -2364
rect 4728 -2404 4740 -2370
rect 4908 -2404 4920 -2370
rect 4728 -2410 4780 -2404
rect 4598 -2472 4666 -2460
rect 4660 -2488 4666 -2472
rect 4660 -2506 4692 -2488
rect 4544 -2726 4692 -2506
rect 4774 -2654 4780 -2410
rect 4868 -2410 4920 -2404
rect 4868 -2654 4874 -2410
rect 4774 -2662 4874 -2654
rect 5074 -2656 5080 -2350
rect 5168 -2656 5174 -2350
rect 5374 -2354 5474 -2090
rect 5530 -2134 5578 -2122
rect 5530 -2310 5536 -2134
rect 5570 -2148 5578 -2134
rect 5638 -2148 5650 -1994
rect 5570 -2294 5650 -2148
rect 5570 -2310 5578 -2294
rect 5530 -2322 5578 -2310
rect 5328 -2360 5520 -2354
rect 5328 -2394 5340 -2360
rect 5508 -2394 5520 -2360
rect 5328 -2400 5520 -2394
rect 5638 -2450 5650 -2294
rect 5582 -2462 5650 -2450
rect 5582 -2482 5588 -2462
rect 5074 -2662 5174 -2656
rect 5276 -2496 5588 -2482
rect 5684 -2496 6112 -1948
rect 7235 -2028 7334 -1444
rect 7372 -1450 7472 -1444
rect 12558 -1490 12730 -960
rect 13494 -1280 23808 -960
rect 23912 -1200 23924 -820
rect 24302 -1200 24312 -820
rect 23912 -1212 24312 -1200
rect 13494 -1484 14010 -1280
rect 14434 -1282 23808 -1280
rect 13494 -1490 13562 -1484
rect 7378 -1500 7478 -1494
rect 7478 -1600 12184 -1500
rect 12284 -1600 12290 -1500
rect 12558 -1582 13562 -1490
rect 7378 -1606 7478 -1600
rect 7378 -1684 7478 -1678
rect 7478 -1784 12006 -1684
rect 12106 -1784 12112 -1684
rect 12424 -1740 13562 -1582
rect 7378 -1790 7478 -1784
rect 7234 -2082 9044 -2028
rect 7234 -2128 7514 -2082
rect 9032 -2128 9044 -2082
rect 7234 -2136 9044 -2128
rect 9222 -2048 9322 -1784
rect 9222 -2092 10966 -2048
rect 3632 -2770 4692 -2726
rect 5276 -2854 6112 -2496
rect 7235 -2612 7334 -2136
rect 9222 -2140 9438 -2092
rect 10952 -2140 10966 -2092
rect 11484 -2088 11576 -2082
rect 11484 -2122 11496 -2088
rect 11564 -2122 11576 -2088
rect 11484 -2128 11576 -2122
rect 9222 -2148 10966 -2140
rect 7432 -2194 7552 -2188
rect 7235 -2685 7336 -2612
rect 2084 -2870 6112 -2854
rect 2084 -3308 3880 -2870
rect 4452 -3308 6112 -2870
rect 7236 -3038 7336 -2685
rect 7432 -2982 7434 -2194
rect 7550 -2982 7552 -2194
rect 7432 -2988 7552 -2982
rect 7592 -2194 7712 -2188
rect 7592 -2982 7594 -2194
rect 7710 -2982 7712 -2194
rect 7592 -2988 7712 -2982
rect 7750 -2194 7870 -2188
rect 7750 -2982 7752 -2194
rect 7868 -2982 7870 -2194
rect 7750 -2988 7870 -2982
rect 7908 -2194 8028 -2188
rect 7908 -2982 7910 -2194
rect 8026 -2982 8028 -2194
rect 7908 -2988 8028 -2982
rect 8066 -2194 8186 -2188
rect 8066 -2982 8068 -2194
rect 8184 -2982 8186 -2194
rect 8066 -2988 8186 -2982
rect 8222 -2192 8342 -2186
rect 8222 -2980 8224 -2192
rect 8340 -2980 8342 -2192
rect 8222 -2986 8342 -2980
rect 8380 -2194 8500 -2188
rect 8380 -2982 8382 -2194
rect 8498 -2982 8500 -2194
rect 8380 -2988 8500 -2982
rect 8540 -2192 8660 -2186
rect 8540 -2980 8542 -2192
rect 8658 -2980 8660 -2192
rect 8540 -2986 8660 -2980
rect 8696 -2194 8816 -2188
rect 8696 -2982 8698 -2194
rect 8814 -2982 8816 -2194
rect 8696 -2988 8816 -2982
rect 8854 -2194 8974 -2188
rect 8854 -2982 8856 -2194
rect 8972 -2982 8974 -2194
rect 8854 -2988 8974 -2982
rect 9012 -2194 9132 -2188
rect 9012 -2982 9014 -2194
rect 9130 -2982 9132 -2194
rect 9012 -2988 9132 -2982
rect 9222 -3036 9322 -2148
rect 11300 -2176 11474 -2164
rect 9358 -2198 9478 -2192
rect 9358 -2986 9360 -2198
rect 9476 -2986 9478 -2198
rect 9358 -2992 9478 -2986
rect 9516 -2198 9636 -2192
rect 9516 -2986 9518 -2198
rect 9634 -2986 9636 -2198
rect 9516 -2992 9636 -2986
rect 9676 -2198 9796 -2192
rect 9676 -2986 9678 -2198
rect 9794 -2986 9796 -2198
rect 9676 -2992 9796 -2986
rect 9834 -2198 9954 -2192
rect 9834 -2986 9836 -2198
rect 9952 -2986 9954 -2198
rect 9834 -2992 9954 -2986
rect 9990 -2198 10110 -2192
rect 9990 -2986 9992 -2198
rect 10108 -2986 10110 -2198
rect 9990 -2992 10110 -2986
rect 10150 -2198 10270 -2192
rect 10150 -2986 10152 -2198
rect 10268 -2986 10270 -2198
rect 10150 -2992 10270 -2986
rect 10306 -2198 10426 -2192
rect 10306 -2986 10308 -2198
rect 10424 -2986 10426 -2198
rect 10306 -2992 10426 -2986
rect 10464 -2198 10584 -2192
rect 10464 -2986 10466 -2198
rect 10582 -2986 10584 -2198
rect 10464 -2992 10584 -2986
rect 10624 -2198 10744 -2192
rect 10624 -2986 10626 -2198
rect 10742 -2986 10744 -2198
rect 10624 -2992 10744 -2986
rect 10780 -2198 10900 -2192
rect 10780 -2986 10782 -2198
rect 10898 -2986 10900 -2198
rect 10780 -2992 10900 -2986
rect 10938 -2198 11058 -2192
rect 10938 -2986 10940 -2198
rect 11056 -2986 11058 -2198
rect 11300 -2964 11310 -2176
rect 11462 -2180 11474 -2176
rect 11468 -2958 11474 -2180
rect 11462 -2964 11474 -2958
rect 11300 -2974 11474 -2964
rect 10938 -2992 11058 -2986
rect 11504 -3010 11550 -2128
rect 12262 -2154 13562 -1740
rect 13662 -1576 13862 -1566
rect 13662 -1756 13672 -1576
rect 13852 -1756 13862 -1576
rect 13914 -1658 14010 -1484
rect 14070 -1362 14782 -1350
rect 14070 -1538 14082 -1362
rect 14770 -1538 14782 -1362
rect 14070 -1542 14782 -1538
rect 13914 -1687 14036 -1658
rect 13914 -1721 13971 -1687
rect 14005 -1721 14036 -1687
rect 13914 -1749 14036 -1721
rect 13662 -1766 13862 -1756
rect 12262 -2156 13048 -2154
rect 11592 -2182 11980 -2170
rect 11592 -2956 11606 -2182
rect 11666 -2956 11980 -2182
rect 11592 -2968 11980 -2956
rect 11772 -2980 11980 -2968
rect 11484 -3012 11576 -3010
rect 11480 -3016 11580 -3012
rect 7236 -3046 9046 -3038
rect 7236 -3092 7512 -3046
rect 9034 -3092 9046 -3046
rect 7236 -3138 9046 -3092
rect 9222 -3044 10966 -3036
rect 9222 -3092 9436 -3044
rect 10952 -3092 10966 -3044
rect 9222 -3136 10966 -3092
rect 11480 -3050 11496 -3016
rect 11564 -3050 11580 -3016
rect 11480 -3198 11580 -3050
rect 11772 -3164 11780 -2980
rect 11972 -3164 11980 -2980
rect 12262 -2224 12634 -2156
rect 12770 -2206 12878 -2156
rect 12770 -2224 12786 -2206
rect 12262 -3148 12616 -2224
rect 12774 -2240 12786 -2224
rect 12862 -2224 12878 -2206
rect 13014 -2224 13048 -2156
rect 12862 -2240 12874 -2224
rect 12774 -2246 12874 -2240
rect 12696 -2268 12742 -2256
rect 12696 -3036 12702 -2268
rect 12736 -2300 12742 -2268
rect 12906 -2268 12952 -2256
rect 12906 -2300 12912 -2268
rect 12736 -2400 12912 -2300
rect 12736 -3036 12742 -2400
rect 12696 -3048 12742 -3036
rect 12906 -3036 12912 -2400
rect 12946 -2300 12952 -2268
rect 13700 -2300 13800 -1766
rect 12946 -2400 13800 -2300
rect 13940 -1779 14036 -1749
rect 13940 -1813 13971 -1779
rect 14005 -1813 14036 -1779
rect 13940 -1871 14036 -1813
rect 14484 -1687 14580 -1542
rect 14484 -1721 14515 -1687
rect 14549 -1721 14580 -1687
rect 14484 -1779 14580 -1721
rect 14866 -1733 23808 -1282
rect 14866 -1750 14897 -1733
rect 14484 -1813 14515 -1779
rect 14549 -1813 14580 -1779
rect 14868 -1767 14897 -1750
rect 14931 -1767 14989 -1733
rect 15023 -1767 15081 -1733
rect 15115 -1767 15173 -1733
rect 15207 -1767 15265 -1733
rect 15299 -1767 15357 -1733
rect 15391 -1767 15449 -1733
rect 15483 -1767 15541 -1733
rect 15575 -1767 15633 -1733
rect 15667 -1767 15725 -1733
rect 15759 -1767 15817 -1733
rect 15851 -1767 15909 -1733
rect 15943 -1767 16001 -1733
rect 16035 -1767 16093 -1733
rect 16127 -1767 16185 -1733
rect 16219 -1767 16277 -1733
rect 16311 -1767 16369 -1733
rect 16403 -1767 16461 -1733
rect 16495 -1767 16553 -1733
rect 16587 -1767 16645 -1733
rect 16679 -1767 16737 -1733
rect 16771 -1767 16829 -1733
rect 16863 -1767 16921 -1733
rect 16955 -1767 17013 -1733
rect 17047 -1767 17105 -1733
rect 17139 -1767 17197 -1733
rect 17231 -1767 17289 -1733
rect 17323 -1767 17381 -1733
rect 17415 -1767 17473 -1733
rect 17507 -1767 17565 -1733
rect 17599 -1767 17657 -1733
rect 17691 -1767 17749 -1733
rect 17783 -1767 17841 -1733
rect 17875 -1767 17933 -1733
rect 17967 -1767 18025 -1733
rect 18059 -1767 18117 -1733
rect 18151 -1767 18209 -1733
rect 18243 -1767 18301 -1733
rect 18335 -1767 18393 -1733
rect 18427 -1767 18485 -1733
rect 18519 -1767 18577 -1733
rect 18611 -1767 18669 -1733
rect 18703 -1767 18761 -1733
rect 18795 -1767 18853 -1733
rect 18887 -1767 18945 -1733
rect 18979 -1767 19037 -1733
rect 19071 -1767 19129 -1733
rect 19163 -1767 19221 -1733
rect 19255 -1767 19313 -1733
rect 19347 -1767 19405 -1733
rect 19439 -1767 19497 -1733
rect 19531 -1767 19589 -1733
rect 19623 -1767 19681 -1733
rect 19715 -1767 19773 -1733
rect 19807 -1767 19865 -1733
rect 19899 -1767 19957 -1733
rect 19991 -1767 20049 -1733
rect 20083 -1767 20141 -1733
rect 20175 -1767 20233 -1733
rect 20267 -1767 20325 -1733
rect 20359 -1767 20417 -1733
rect 20451 -1767 20509 -1733
rect 20543 -1767 20601 -1733
rect 20635 -1767 20693 -1733
rect 20727 -1767 20785 -1733
rect 20819 -1767 20877 -1733
rect 20911 -1767 20969 -1733
rect 21003 -1767 21061 -1733
rect 21095 -1767 21153 -1733
rect 21187 -1767 21245 -1733
rect 21279 -1767 21337 -1733
rect 21371 -1767 21429 -1733
rect 21463 -1767 21521 -1733
rect 21555 -1767 21613 -1733
rect 21647 -1767 21705 -1733
rect 21739 -1767 21797 -1733
rect 21831 -1767 21889 -1733
rect 21923 -1767 21981 -1733
rect 22015 -1767 22073 -1733
rect 22107 -1767 23808 -1733
rect 14868 -1798 23808 -1767
rect 13940 -1905 13971 -1871
rect 14005 -1905 14036 -1871
rect 13940 -1963 14036 -1905
rect 13940 -1997 13971 -1963
rect 14005 -1997 14036 -1963
rect 14188 -1872 14436 -1858
rect 14188 -1964 14202 -1872
rect 14422 -1964 14436 -1872
rect 14188 -1978 14436 -1964
rect 14484 -1871 14580 -1813
rect 14484 -1905 14515 -1871
rect 14549 -1905 14580 -1871
rect 14484 -1963 14580 -1905
rect 14726 -1848 14826 -1836
rect 14726 -1924 14738 -1848
rect 14814 -1860 14826 -1848
rect 14814 -1897 21452 -1860
rect 14814 -1903 21455 -1897
rect 14814 -1910 16273 -1903
rect 14814 -1924 14826 -1910
rect 14726 -1936 14826 -1924
rect 16261 -1937 16273 -1910
rect 16307 -1937 16345 -1903
rect 16379 -1934 16993 -1903
rect 16379 -1937 16391 -1934
rect 16261 -1943 16391 -1937
rect 16896 -1937 16993 -1934
rect 17027 -1910 18481 -1903
rect 17027 -1937 17039 -1910
rect 16896 -1943 17039 -1937
rect 18469 -1937 18481 -1910
rect 18515 -1937 18553 -1903
rect 18587 -1934 19201 -1903
rect 18587 -1937 18599 -1934
rect 18469 -1943 18599 -1937
rect 19104 -1937 19201 -1934
rect 19235 -1910 20689 -1903
rect 19235 -1937 19247 -1910
rect 19104 -1943 19247 -1937
rect 20677 -1937 20689 -1910
rect 20723 -1937 20761 -1903
rect 20795 -1934 21409 -1903
rect 20795 -1937 20807 -1934
rect 20677 -1943 20807 -1937
rect 21312 -1937 21409 -1934
rect 21443 -1937 21455 -1903
rect 21312 -1943 21455 -1937
rect 13940 -2055 14036 -1997
rect 14484 -1997 14515 -1963
rect 14549 -1997 14580 -1963
rect 15622 -1971 15680 -1965
rect 13940 -2089 13971 -2055
rect 14005 -2089 14036 -2055
rect 14124 -2024 14244 -2018
rect 14124 -2076 14132 -2024
rect 14238 -2076 14244 -2024
rect 14124 -2082 14244 -2076
rect 14484 -2055 14580 -1997
rect 14968 -1988 15052 -1976
rect 13940 -2147 14036 -2089
rect 14484 -2089 14515 -2055
rect 14549 -2089 14580 -2055
rect 13940 -2181 13971 -2147
rect 14005 -2181 14036 -2147
rect 13940 -2239 14036 -2181
rect 14124 -2150 14244 -2144
rect 14124 -2202 14132 -2150
rect 14238 -2202 14244 -2150
rect 14124 -2208 14244 -2202
rect 14484 -2147 14580 -2089
rect 14726 -2022 14826 -2012
rect 14968 -2022 14980 -1988
rect 14726 -2026 14980 -2022
rect 14726 -2098 14740 -2026
rect 14812 -2098 14980 -2026
rect 14726 -2102 14980 -2098
rect 14726 -2112 14826 -2102
rect 14484 -2181 14515 -2147
rect 14549 -2181 14580 -2147
rect 14968 -2140 14980 -2102
rect 15040 -2140 15052 -1988
rect 15148 -1982 15232 -1976
rect 15148 -2090 15154 -1982
rect 15226 -2090 15232 -1982
rect 15622 -2005 15634 -1971
rect 15668 -1974 15680 -1971
rect 15989 -1971 16047 -1965
rect 15989 -1974 16001 -1971
rect 15668 -2002 16001 -1974
rect 15668 -2005 15680 -2002
rect 15622 -2011 15680 -2005
rect 15989 -2005 16001 -2002
rect 16035 -1974 16047 -1971
rect 16705 -1971 16763 -1965
rect 16705 -1974 16717 -1971
rect 16035 -2002 16717 -1974
rect 16035 -2005 16047 -2002
rect 15989 -2011 16047 -2005
rect 16705 -2005 16717 -2002
rect 16751 -2005 16763 -1971
rect 16896 -1966 17036 -1943
rect 16896 -2000 16933 -1966
rect 16967 -2000 17036 -1966
rect 16896 -2004 17036 -2000
rect 17830 -1971 17888 -1965
rect 16705 -2011 16763 -2005
rect 16921 -2006 16979 -2004
rect 17830 -2005 17842 -1971
rect 17876 -1974 17888 -1971
rect 18197 -1971 18255 -1965
rect 18197 -1974 18209 -1971
rect 17876 -2002 18209 -1974
rect 17876 -2005 17888 -2002
rect 17830 -2011 17888 -2005
rect 18197 -2005 18209 -2002
rect 18243 -1974 18255 -1971
rect 18913 -1971 18971 -1965
rect 18913 -1974 18925 -1971
rect 18243 -2002 18925 -1974
rect 18243 -2005 18255 -2002
rect 18197 -2011 18255 -2005
rect 18913 -2005 18925 -2002
rect 18959 -2005 18971 -1971
rect 19104 -1966 19244 -1943
rect 19104 -2000 19141 -1966
rect 19175 -2000 19244 -1966
rect 19104 -2004 19244 -2000
rect 20038 -1971 20096 -1965
rect 18913 -2011 18971 -2005
rect 19129 -2006 19187 -2004
rect 20038 -2005 20050 -1971
rect 20084 -1974 20096 -1971
rect 20405 -1971 20463 -1965
rect 20405 -1974 20417 -1971
rect 20084 -2002 20417 -1974
rect 20084 -2005 20096 -2002
rect 20038 -2011 20096 -2005
rect 20405 -2005 20417 -2002
rect 20451 -1974 20463 -1971
rect 21121 -1971 21179 -1965
rect 21121 -1974 21133 -1971
rect 20451 -2002 21133 -1974
rect 20451 -2005 20463 -2002
rect 20405 -2011 20463 -2005
rect 21121 -2005 21133 -2002
rect 21167 -2005 21179 -1971
rect 21312 -1966 21452 -1943
rect 21312 -2000 21349 -1966
rect 21383 -2000 21452 -1966
rect 21312 -2004 21452 -2000
rect 21954 -1952 22034 -1942
rect 21121 -2011 21179 -2005
rect 21337 -2006 21395 -2004
rect 15796 -2036 15886 -2030
rect 15796 -2076 15814 -2036
rect 15854 -2040 15886 -2036
rect 18004 -2036 18094 -2030
rect 15854 -2050 17608 -2040
rect 15854 -2072 17556 -2050
rect 15854 -2076 15886 -2072
rect 15796 -2082 15886 -2076
rect 15148 -2096 15232 -2090
rect 17548 -2088 17556 -2072
rect 17594 -2088 17608 -2050
rect 18004 -2076 18022 -2036
rect 18062 -2040 18094 -2036
rect 20212 -2036 20302 -2030
rect 18062 -2050 19816 -2040
rect 18062 -2072 19766 -2050
rect 18062 -2076 18094 -2072
rect 18004 -2082 18094 -2076
rect 17548 -2100 17608 -2088
rect 19756 -2088 19766 -2072
rect 19804 -2088 19816 -2050
rect 20212 -2076 20230 -2036
rect 20270 -2040 20302 -2036
rect 21954 -2040 21962 -1952
rect 20270 -2072 21962 -2040
rect 20270 -2076 20302 -2072
rect 20212 -2082 20302 -2076
rect 19756 -2100 19816 -2088
rect 14968 -2152 15052 -2140
rect 15703 -2107 15761 -2101
rect 15703 -2141 15715 -2107
rect 15749 -2110 15761 -2107
rect 16081 -2107 16139 -2101
rect 16081 -2110 16093 -2107
rect 15749 -2138 16093 -2110
rect 15749 -2141 15761 -2138
rect 15703 -2147 15761 -2141
rect 16081 -2141 16093 -2138
rect 16127 -2110 16139 -2107
rect 16705 -2107 16763 -2101
rect 16705 -2110 16717 -2107
rect 16127 -2138 16717 -2110
rect 16127 -2141 16139 -2138
rect 16081 -2147 16139 -2141
rect 16705 -2141 16717 -2138
rect 16751 -2141 16763 -2107
rect 16705 -2147 16763 -2141
rect 17911 -2107 17969 -2101
rect 17911 -2141 17923 -2107
rect 17957 -2110 17969 -2107
rect 18289 -2107 18347 -2101
rect 18289 -2110 18301 -2107
rect 17957 -2138 18301 -2110
rect 17957 -2141 17969 -2138
rect 17911 -2147 17969 -2141
rect 18289 -2141 18301 -2138
rect 18335 -2110 18347 -2107
rect 18913 -2107 18971 -2101
rect 18913 -2110 18925 -2107
rect 18335 -2138 18925 -2110
rect 18335 -2141 18347 -2138
rect 18289 -2147 18347 -2141
rect 18913 -2141 18925 -2138
rect 18959 -2141 18971 -2107
rect 18913 -2147 18971 -2141
rect 20119 -2107 20177 -2101
rect 20119 -2141 20131 -2107
rect 20165 -2110 20177 -2107
rect 20497 -2107 20555 -2101
rect 20497 -2110 20509 -2107
rect 20165 -2138 20509 -2110
rect 20165 -2141 20177 -2138
rect 20119 -2147 20177 -2141
rect 20497 -2141 20509 -2138
rect 20543 -2110 20555 -2107
rect 21121 -2107 21179 -2101
rect 21121 -2110 21133 -2107
rect 20543 -2138 21133 -2110
rect 20543 -2141 20555 -2138
rect 20497 -2147 20555 -2141
rect 21121 -2141 21133 -2138
rect 21167 -2141 21179 -2107
rect 21121 -2147 21179 -2141
rect 13940 -2273 13971 -2239
rect 14005 -2273 14036 -2239
rect 14484 -2239 14580 -2181
rect 21954 -2174 21962 -2072
rect 22026 -2174 22034 -1952
rect 21954 -2182 22034 -2174
rect 13940 -2331 14036 -2273
rect 13940 -2365 13971 -2331
rect 14005 -2365 14036 -2331
rect 14186 -2250 14434 -2244
rect 14186 -2258 14204 -2250
rect 14242 -2258 14434 -2250
rect 14186 -2350 14200 -2258
rect 14420 -2350 14434 -2258
rect 14186 -2364 14434 -2350
rect 14484 -2273 14515 -2239
rect 14549 -2246 14580 -2239
rect 22136 -2246 22146 -1854
rect 14549 -2273 22146 -2246
rect 14484 -2277 22146 -2273
rect 14484 -2311 14897 -2277
rect 14931 -2311 14989 -2277
rect 15023 -2311 15081 -2277
rect 15115 -2311 15173 -2277
rect 15207 -2311 15265 -2277
rect 15299 -2311 15357 -2277
rect 15391 -2311 15449 -2277
rect 15483 -2311 15541 -2277
rect 15575 -2311 15633 -2277
rect 15667 -2311 15725 -2277
rect 15759 -2311 15817 -2277
rect 15851 -2311 15909 -2277
rect 15943 -2311 16001 -2277
rect 16035 -2311 16093 -2277
rect 16127 -2311 16185 -2277
rect 16219 -2311 16277 -2277
rect 16311 -2311 16369 -2277
rect 16403 -2311 16461 -2277
rect 16495 -2311 16553 -2277
rect 16587 -2311 16645 -2277
rect 16679 -2311 16737 -2277
rect 16771 -2311 16829 -2277
rect 16863 -2311 16921 -2277
rect 16955 -2311 17013 -2277
rect 17047 -2311 17105 -2277
rect 17139 -2311 17197 -2277
rect 17231 -2311 17289 -2277
rect 17323 -2311 17381 -2277
rect 17415 -2311 17473 -2277
rect 17507 -2311 17565 -2277
rect 17599 -2311 17657 -2277
rect 17691 -2311 17749 -2277
rect 17783 -2311 17841 -2277
rect 17875 -2311 17933 -2277
rect 17967 -2311 18025 -2277
rect 18059 -2311 18117 -2277
rect 18151 -2311 18209 -2277
rect 18243 -2311 18301 -2277
rect 18335 -2311 18393 -2277
rect 18427 -2311 18485 -2277
rect 18519 -2311 18577 -2277
rect 18611 -2311 18669 -2277
rect 18703 -2311 18761 -2277
rect 18795 -2311 18853 -2277
rect 18887 -2311 18945 -2277
rect 18979 -2311 19037 -2277
rect 19071 -2311 19129 -2277
rect 19163 -2311 19221 -2277
rect 19255 -2311 19313 -2277
rect 19347 -2311 19405 -2277
rect 19439 -2311 19497 -2277
rect 19531 -2311 19589 -2277
rect 19623 -2311 19681 -2277
rect 19715 -2311 19773 -2277
rect 19807 -2311 19865 -2277
rect 19899 -2311 19957 -2277
rect 19991 -2311 20049 -2277
rect 20083 -2311 20141 -2277
rect 20175 -2311 20233 -2277
rect 20267 -2311 20325 -2277
rect 20359 -2311 20417 -2277
rect 20451 -2311 20509 -2277
rect 20543 -2311 20601 -2277
rect 20635 -2311 20693 -2277
rect 20727 -2311 20785 -2277
rect 20819 -2311 20877 -2277
rect 20911 -2311 20969 -2277
rect 21003 -2311 21061 -2277
rect 21095 -2311 21153 -2277
rect 21187 -2311 21245 -2277
rect 21279 -2311 21337 -2277
rect 21371 -2311 21429 -2277
rect 21463 -2311 21521 -2277
rect 21555 -2311 21613 -2277
rect 21647 -2311 21705 -2277
rect 21739 -2311 21797 -2277
rect 21831 -2311 21889 -2277
rect 21923 -2311 21981 -2277
rect 22015 -2311 22073 -2277
rect 22107 -2311 22146 -2277
rect 14484 -2331 22146 -2311
rect 12946 -3036 12952 -2400
rect 13940 -2423 14036 -2365
rect 13940 -2446 13971 -2423
rect 12906 -3048 12952 -3036
rect 13028 -2457 13971 -2446
rect 14005 -2457 14036 -2423
rect 14484 -2365 14515 -2331
rect 14549 -2342 22146 -2331
rect 14549 -2365 14580 -2342
rect 14484 -2423 14580 -2365
rect 13028 -2468 14036 -2457
rect 13028 -3026 13052 -2468
rect 13648 -2515 14036 -2468
rect 13648 -2549 13971 -2515
rect 14005 -2549 14036 -2515
rect 13648 -2607 14036 -2549
rect 13648 -2641 13971 -2607
rect 14005 -2641 14036 -2607
rect 13648 -2699 14036 -2641
rect 13648 -2733 13971 -2699
rect 14005 -2733 14036 -2699
rect 13648 -2791 14036 -2733
rect 13648 -2825 13971 -2791
rect 14005 -2825 14036 -2791
rect 14186 -2472 14332 -2450
rect 14186 -2572 14208 -2472
rect 14308 -2572 14332 -2472
rect 14186 -2616 14332 -2572
rect 14484 -2457 14515 -2423
rect 14549 -2457 14580 -2423
rect 21954 -2414 22034 -2406
rect 14484 -2515 14580 -2457
rect 14968 -2448 15052 -2436
rect 14484 -2549 14515 -2515
rect 14549 -2549 14580 -2515
rect 14484 -2607 14580 -2549
rect 14726 -2486 14826 -2476
rect 14968 -2486 14980 -2448
rect 14726 -2490 14980 -2486
rect 14726 -2562 14740 -2490
rect 14812 -2562 14980 -2490
rect 14726 -2566 14980 -2562
rect 14726 -2576 14826 -2566
rect 14186 -2748 14266 -2616
rect 14186 -2816 14192 -2748
rect 14260 -2816 14266 -2748
rect 14186 -2822 14266 -2816
rect 14484 -2641 14515 -2607
rect 14549 -2641 14580 -2607
rect 14968 -2600 14980 -2566
rect 15040 -2600 15052 -2448
rect 15703 -2447 15761 -2441
rect 15703 -2481 15715 -2447
rect 15749 -2450 15761 -2447
rect 16081 -2447 16139 -2441
rect 16081 -2450 16093 -2447
rect 15749 -2478 16093 -2450
rect 15749 -2481 15761 -2478
rect 15703 -2487 15761 -2481
rect 16081 -2481 16093 -2478
rect 16127 -2450 16139 -2447
rect 16705 -2447 16763 -2441
rect 16705 -2450 16717 -2447
rect 16127 -2478 16717 -2450
rect 16127 -2481 16139 -2478
rect 16081 -2487 16139 -2481
rect 16705 -2481 16717 -2478
rect 16751 -2481 16763 -2447
rect 16705 -2487 16763 -2481
rect 17911 -2447 17969 -2441
rect 17911 -2481 17923 -2447
rect 17957 -2450 17969 -2447
rect 18289 -2447 18347 -2441
rect 18289 -2450 18301 -2447
rect 17957 -2478 18301 -2450
rect 17957 -2481 17969 -2478
rect 17911 -2487 17969 -2481
rect 18289 -2481 18301 -2478
rect 18335 -2450 18347 -2447
rect 18913 -2447 18971 -2441
rect 18913 -2450 18925 -2447
rect 18335 -2478 18925 -2450
rect 18335 -2481 18347 -2478
rect 18289 -2487 18347 -2481
rect 18913 -2481 18925 -2478
rect 18959 -2481 18971 -2447
rect 18913 -2487 18971 -2481
rect 20119 -2447 20177 -2441
rect 20119 -2481 20131 -2447
rect 20165 -2450 20177 -2447
rect 20497 -2447 20555 -2441
rect 20497 -2450 20509 -2447
rect 20165 -2478 20509 -2450
rect 20165 -2481 20177 -2478
rect 20119 -2487 20177 -2481
rect 20497 -2481 20509 -2478
rect 20543 -2450 20555 -2447
rect 21121 -2447 21179 -2441
rect 21121 -2450 21133 -2447
rect 20543 -2478 21133 -2450
rect 20543 -2481 20555 -2478
rect 20497 -2487 20555 -2481
rect 21121 -2481 21133 -2478
rect 21167 -2481 21179 -2447
rect 21121 -2487 21179 -2481
rect 14968 -2612 15052 -2600
rect 15148 -2498 15232 -2492
rect 15148 -2606 15154 -2498
rect 15226 -2606 15232 -2498
rect 17548 -2500 17608 -2488
rect 15796 -2512 15886 -2506
rect 15796 -2552 15814 -2512
rect 15854 -2516 15886 -2512
rect 17548 -2516 17556 -2500
rect 15854 -2538 17556 -2516
rect 17594 -2538 17608 -2500
rect 19756 -2500 19816 -2488
rect 15854 -2548 17608 -2538
rect 18004 -2512 18094 -2506
rect 15854 -2552 15886 -2548
rect 15796 -2558 15886 -2552
rect 18004 -2552 18022 -2512
rect 18062 -2516 18094 -2512
rect 19756 -2516 19766 -2500
rect 18062 -2538 19766 -2516
rect 19804 -2538 19816 -2500
rect 18062 -2548 19816 -2538
rect 20212 -2512 20302 -2506
rect 18062 -2552 18094 -2548
rect 18004 -2558 18094 -2552
rect 20212 -2552 20230 -2512
rect 20270 -2516 20302 -2512
rect 21954 -2516 21962 -2414
rect 20270 -2548 21962 -2516
rect 20270 -2552 20302 -2548
rect 20212 -2558 20302 -2552
rect 15148 -2612 15232 -2606
rect 15622 -2583 15680 -2577
rect 15622 -2617 15634 -2583
rect 15668 -2586 15680 -2583
rect 15989 -2583 16047 -2577
rect 15989 -2586 16001 -2583
rect 15668 -2614 16001 -2586
rect 15668 -2617 15680 -2614
rect 15622 -2623 15680 -2617
rect 15989 -2617 16001 -2614
rect 16035 -2586 16047 -2583
rect 16705 -2583 16763 -2577
rect 16705 -2586 16717 -2583
rect 16035 -2614 16717 -2586
rect 16035 -2617 16047 -2614
rect 15989 -2623 16047 -2617
rect 16705 -2617 16717 -2614
rect 16751 -2617 16763 -2583
rect 16921 -2584 16979 -2582
rect 17830 -2583 17888 -2577
rect 16705 -2623 16763 -2617
rect 16896 -2588 17036 -2584
rect 16896 -2622 16933 -2588
rect 16967 -2622 17036 -2588
rect 14484 -2699 14580 -2641
rect 16896 -2645 17036 -2622
rect 17830 -2617 17842 -2583
rect 17876 -2586 17888 -2583
rect 18197 -2583 18255 -2577
rect 18197 -2586 18209 -2583
rect 17876 -2614 18209 -2586
rect 17876 -2617 17888 -2614
rect 17830 -2623 17888 -2617
rect 18197 -2617 18209 -2614
rect 18243 -2586 18255 -2583
rect 18913 -2583 18971 -2577
rect 18913 -2586 18925 -2583
rect 18243 -2614 18925 -2586
rect 18243 -2617 18255 -2614
rect 18197 -2623 18255 -2617
rect 18913 -2617 18925 -2614
rect 18959 -2617 18971 -2583
rect 19129 -2584 19187 -2582
rect 20038 -2583 20096 -2577
rect 18913 -2623 18971 -2617
rect 19104 -2588 19244 -2584
rect 19104 -2622 19141 -2588
rect 19175 -2622 19244 -2588
rect 19104 -2645 19244 -2622
rect 20038 -2617 20050 -2583
rect 20084 -2586 20096 -2583
rect 20405 -2583 20463 -2577
rect 20405 -2586 20417 -2583
rect 20084 -2614 20417 -2586
rect 20084 -2617 20096 -2614
rect 20038 -2623 20096 -2617
rect 20405 -2617 20417 -2614
rect 20451 -2586 20463 -2583
rect 21121 -2583 21179 -2577
rect 21121 -2586 21133 -2583
rect 20451 -2614 21133 -2586
rect 20451 -2617 20463 -2614
rect 20405 -2623 20463 -2617
rect 21121 -2617 21133 -2614
rect 21167 -2617 21179 -2583
rect 21337 -2584 21395 -2582
rect 21121 -2623 21179 -2617
rect 21312 -2588 21452 -2584
rect 21312 -2622 21349 -2588
rect 21383 -2622 21452 -2588
rect 21312 -2645 21452 -2622
rect 21954 -2636 21962 -2548
rect 22026 -2636 22034 -2414
rect 16261 -2651 16391 -2645
rect 14484 -2733 14515 -2699
rect 14549 -2733 14580 -2699
rect 14484 -2791 14580 -2733
rect 14726 -2664 14826 -2652
rect 14726 -2740 14738 -2664
rect 14814 -2678 14826 -2664
rect 16261 -2678 16273 -2651
rect 14814 -2685 16273 -2678
rect 16307 -2685 16345 -2651
rect 16379 -2654 16391 -2651
rect 16896 -2651 17039 -2645
rect 16896 -2654 16993 -2651
rect 16379 -2685 16993 -2654
rect 17027 -2678 17039 -2651
rect 18469 -2651 18599 -2645
rect 18469 -2678 18481 -2651
rect 17027 -2685 18481 -2678
rect 18515 -2685 18553 -2651
rect 18587 -2654 18599 -2651
rect 19104 -2651 19247 -2645
rect 19104 -2654 19201 -2651
rect 18587 -2685 19201 -2654
rect 19235 -2678 19247 -2651
rect 20677 -2651 20807 -2645
rect 20677 -2678 20689 -2651
rect 19235 -2685 20689 -2678
rect 20723 -2685 20761 -2651
rect 20795 -2654 20807 -2651
rect 21312 -2651 21455 -2645
rect 21954 -2646 22034 -2636
rect 21312 -2654 21409 -2651
rect 20795 -2685 21409 -2654
rect 21443 -2685 21455 -2651
rect 14814 -2691 21455 -2685
rect 14814 -2728 21452 -2691
rect 14814 -2740 14826 -2728
rect 22136 -2734 22146 -2342
rect 22288 -2734 22300 -1854
rect 14726 -2752 14826 -2740
rect 22362 -2790 23808 -1798
rect 13648 -2854 14036 -2825
rect 14484 -2825 14515 -2791
rect 14549 -2825 14580 -2791
rect 14484 -2854 14580 -2825
rect 14868 -2821 23808 -2790
rect 13648 -3026 13960 -2854
rect 14868 -2855 14897 -2821
rect 14931 -2855 14989 -2821
rect 15023 -2855 15081 -2821
rect 15115 -2855 15173 -2821
rect 15207 -2855 15265 -2821
rect 15299 -2855 15357 -2821
rect 15391 -2855 15449 -2821
rect 15483 -2855 15541 -2821
rect 15575 -2855 15633 -2821
rect 15667 -2855 15725 -2821
rect 15759 -2855 15817 -2821
rect 15851 -2855 15909 -2821
rect 15943 -2855 16001 -2821
rect 16035 -2855 16093 -2821
rect 16127 -2855 16185 -2821
rect 16219 -2855 16277 -2821
rect 16311 -2855 16369 -2821
rect 16403 -2855 16461 -2821
rect 16495 -2855 16553 -2821
rect 16587 -2855 16645 -2821
rect 16679 -2855 16737 -2821
rect 16771 -2855 16829 -2821
rect 16863 -2855 16921 -2821
rect 16955 -2855 17013 -2821
rect 17047 -2855 17105 -2821
rect 17139 -2855 17197 -2821
rect 17231 -2855 17289 -2821
rect 17323 -2855 17381 -2821
rect 17415 -2855 17473 -2821
rect 17507 -2855 17565 -2821
rect 17599 -2855 17657 -2821
rect 17691 -2855 17749 -2821
rect 17783 -2855 17841 -2821
rect 17875 -2855 17933 -2821
rect 17967 -2855 18025 -2821
rect 18059 -2855 18117 -2821
rect 18151 -2855 18209 -2821
rect 18243 -2855 18301 -2821
rect 18335 -2855 18393 -2821
rect 18427 -2855 18485 -2821
rect 18519 -2855 18577 -2821
rect 18611 -2855 18669 -2821
rect 18703 -2855 18761 -2821
rect 18795 -2855 18853 -2821
rect 18887 -2855 18945 -2821
rect 18979 -2855 19037 -2821
rect 19071 -2855 19129 -2821
rect 19163 -2855 19221 -2821
rect 19255 -2855 19313 -2821
rect 19347 -2855 19405 -2821
rect 19439 -2855 19497 -2821
rect 19531 -2855 19589 -2821
rect 19623 -2855 19681 -2821
rect 19715 -2855 19773 -2821
rect 19807 -2855 19865 -2821
rect 19899 -2855 19957 -2821
rect 19991 -2855 20049 -2821
rect 20083 -2855 20141 -2821
rect 20175 -2855 20233 -2821
rect 20267 -2855 20325 -2821
rect 20359 -2855 20417 -2821
rect 20451 -2855 20509 -2821
rect 20543 -2855 20601 -2821
rect 20635 -2855 20693 -2821
rect 20727 -2855 20785 -2821
rect 20819 -2855 20877 -2821
rect 20911 -2855 20969 -2821
rect 21003 -2855 21061 -2821
rect 21095 -2855 21153 -2821
rect 21187 -2855 21245 -2821
rect 21279 -2855 21337 -2821
rect 21371 -2855 21429 -2821
rect 21463 -2855 21521 -2821
rect 21555 -2855 21613 -2821
rect 21647 -2855 21705 -2821
rect 21739 -2855 21797 -2821
rect 21831 -2855 21889 -2821
rect 21923 -2855 21981 -2821
rect 22015 -2855 22073 -2821
rect 22107 -2855 23808 -2821
rect 14868 -2886 23808 -2855
rect 14022 -2902 14532 -2886
rect 14022 -2982 14040 -2902
rect 14140 -2982 14414 -2902
rect 14514 -2982 14532 -2902
rect 14022 -2998 14532 -2982
rect 13028 -3044 13960 -3026
rect 12774 -3062 12874 -3058
rect 11772 -3172 11980 -3164
rect 2084 -3330 6112 -3308
rect 11416 -3208 11616 -3198
rect 11416 -3386 11426 -3208
rect 11604 -3386 11616 -3208
rect 11416 -3398 11616 -3386
rect 12260 -3216 12616 -3148
rect 2300 -3594 6034 -3578
rect 1626 -3600 6034 -3594
rect 1626 -5026 1636 -3600
rect 1920 -3770 6034 -3600
rect 12260 -3630 12462 -3216
rect 12588 -3390 12616 -3216
rect 12772 -3064 12874 -3062
rect 12772 -3098 12786 -3064
rect 12862 -3098 12874 -3064
rect 12772 -3176 12874 -3098
rect 13936 -3124 14136 -3116
rect 13936 -3176 13942 -3124
rect 12772 -3294 13942 -3176
rect 12588 -3416 13840 -3390
rect 13646 -3630 13840 -3416
rect 13936 -3470 13942 -3294
rect 14128 -3470 14136 -3124
rect 13936 -3476 14136 -3470
rect 14332 -3152 14532 -2998
rect 16052 -3004 23808 -2886
rect 15160 -3048 15950 -3036
rect 15160 -3128 15172 -3048
rect 15938 -3088 15950 -3048
rect 15938 -3094 15952 -3088
rect 15940 -3128 15952 -3094
rect 15160 -3134 15952 -3128
rect 14332 -3464 14344 -3152
rect 14520 -3166 14532 -3152
rect 16052 -3166 16120 -3004
rect 16212 -3136 23808 -3004
rect 14520 -3178 15150 -3166
rect 14520 -3254 15110 -3178
rect 15144 -3254 15150 -3178
rect 14520 -3266 15150 -3254
rect 15962 -3178 16120 -3166
rect 15962 -3254 15968 -3178
rect 16002 -3254 16120 -3178
rect 15962 -3266 16120 -3254
rect 14520 -3464 14532 -3266
rect 15160 -3304 15952 -3298
rect 15160 -3338 15172 -3304
rect 15940 -3338 15952 -3304
rect 15160 -3344 15952 -3338
rect 16104 -3422 16120 -3266
rect 14332 -3476 14532 -3464
rect 15008 -3442 16120 -3422
rect 15008 -3516 15034 -3442
rect 17524 -3514 23808 -3136
rect 16212 -3516 23808 -3514
rect 15008 -3534 23808 -3516
rect 1920 -3916 6036 -3770
rect 1920 -3918 3162 -3916
rect 1920 -4936 2456 -3918
rect 2552 -3962 3162 -3918
rect 2552 -4326 2592 -3962
rect 2662 -4034 2728 -4028
rect 2662 -4088 2668 -4034
rect 2722 -4036 2728 -4034
rect 2722 -4054 2982 -4036
rect 2722 -4088 2744 -4054
rect 2812 -4088 2902 -4054
rect 2970 -4088 2982 -4054
rect 2662 -4094 2982 -4088
rect 2672 -4138 2724 -4126
rect 2672 -4326 2682 -4138
rect 2552 -4526 2682 -4326
rect 2552 -4890 2592 -4526
rect 2672 -4714 2682 -4526
rect 2716 -4714 2724 -4138
rect 2672 -4726 2724 -4714
rect 2756 -4134 2958 -4126
rect 2756 -4716 2766 -4134
rect 2950 -4716 2958 -4134
rect 2756 -4724 2958 -4716
rect 2992 -4138 3038 -4126
rect 2992 -4714 2998 -4138
rect 3032 -4326 3038 -4138
rect 3118 -4326 3162 -3962
rect 3032 -4526 3162 -4326
rect 3032 -4714 3038 -4526
rect 2834 -4726 2880 -4724
rect 2992 -4726 3038 -4714
rect 2662 -4764 2982 -4758
rect 2662 -4818 2668 -4764
rect 2722 -4798 2744 -4764
rect 2812 -4798 2902 -4764
rect 2970 -4798 2982 -4764
rect 2722 -4816 2982 -4798
rect 2722 -4818 2728 -4816
rect 2662 -4824 2728 -4818
rect 3118 -4890 3162 -4526
rect 2552 -4934 3162 -4890
rect 3258 -3962 3870 -3916
rect 3258 -4326 3302 -3962
rect 3692 -4034 3758 -4028
rect 3692 -4036 3698 -4034
rect 3438 -4054 3698 -4036
rect 3438 -4088 3450 -4054
rect 3518 -4088 3608 -4054
rect 3676 -4088 3698 -4054
rect 3752 -4088 3758 -4034
rect 3438 -4094 3758 -4088
rect 3382 -4138 3428 -4126
rect 3382 -4326 3388 -4138
rect 3258 -4526 3388 -4326
rect 3258 -4890 3302 -4526
rect 3382 -4714 3388 -4526
rect 3422 -4714 3428 -4138
rect 3382 -4726 3428 -4714
rect 3462 -4134 3664 -4126
rect 3462 -4716 3472 -4134
rect 3656 -4716 3664 -4134
rect 3462 -4724 3664 -4716
rect 3698 -4138 3748 -4126
rect 3698 -4714 3704 -4138
rect 3738 -4326 3748 -4138
rect 3828 -4326 3870 -3962
rect 3738 -4526 3870 -4326
rect 3738 -4714 3748 -4526
rect 3540 -4726 3586 -4724
rect 3698 -4726 3748 -4714
rect 3438 -4764 3758 -4758
rect 3438 -4798 3450 -4764
rect 3518 -4798 3608 -4764
rect 3676 -4798 3698 -4764
rect 3438 -4816 3698 -4798
rect 3692 -4818 3698 -4816
rect 3752 -4818 3758 -4764
rect 3692 -4824 3758 -4818
rect 3828 -4890 3870 -4526
rect 3258 -4934 3870 -4890
rect 3966 -4934 4370 -3916
rect 4466 -3962 5078 -3916
rect 4466 -4326 4508 -3962
rect 4578 -4034 4644 -4028
rect 4578 -4088 4584 -4034
rect 4638 -4036 4644 -4034
rect 4638 -4054 4898 -4036
rect 4638 -4088 4660 -4054
rect 4728 -4088 4818 -4054
rect 4886 -4088 4898 -4054
rect 4578 -4094 4898 -4088
rect 4588 -4138 4638 -4126
rect 4588 -4326 4598 -4138
rect 4466 -4526 4598 -4326
rect 4466 -4890 4508 -4526
rect 4588 -4714 4598 -4526
rect 4632 -4714 4638 -4138
rect 4588 -4726 4638 -4714
rect 4672 -4134 4874 -4126
rect 4672 -4716 4680 -4134
rect 4864 -4716 4874 -4134
rect 4672 -4724 4874 -4716
rect 4908 -4138 4954 -4126
rect 4908 -4714 4914 -4138
rect 4948 -4326 4954 -4138
rect 5034 -4326 5078 -3962
rect 4948 -4526 5078 -4326
rect 4948 -4714 4954 -4526
rect 4750 -4726 4796 -4724
rect 4908 -4726 4954 -4714
rect 4578 -4764 4898 -4758
rect 4578 -4818 4584 -4764
rect 4638 -4798 4660 -4764
rect 4728 -4798 4818 -4764
rect 4886 -4798 4898 -4764
rect 4638 -4816 4898 -4798
rect 4638 -4818 4644 -4816
rect 4578 -4824 4644 -4818
rect 5034 -4890 5078 -4526
rect 4466 -4934 5078 -4890
rect 5174 -3918 6036 -3916
rect 5174 -3962 5784 -3918
rect 5174 -4326 5218 -3962
rect 5608 -4034 5674 -4028
rect 5608 -4036 5614 -4034
rect 5354 -4054 5614 -4036
rect 5354 -4088 5366 -4054
rect 5434 -4088 5524 -4054
rect 5592 -4088 5614 -4054
rect 5668 -4088 5674 -4034
rect 5354 -4094 5674 -4088
rect 5298 -4138 5344 -4126
rect 5298 -4326 5304 -4138
rect 5174 -4526 5304 -4326
rect 5174 -4890 5218 -4526
rect 5298 -4714 5304 -4526
rect 5338 -4714 5344 -4138
rect 5298 -4726 5344 -4714
rect 5378 -4134 5580 -4126
rect 5378 -4716 5386 -4134
rect 5570 -4716 5580 -4134
rect 5378 -4724 5580 -4716
rect 5612 -4138 5664 -4126
rect 5612 -4714 5620 -4138
rect 5654 -4326 5664 -4138
rect 5744 -4326 5784 -3962
rect 5654 -4526 5784 -4326
rect 5654 -4714 5664 -4526
rect 5456 -4726 5502 -4724
rect 5612 -4726 5664 -4714
rect 5354 -4764 5674 -4758
rect 5354 -4798 5366 -4764
rect 5434 -4798 5524 -4764
rect 5592 -4798 5614 -4764
rect 5354 -4816 5614 -4798
rect 5608 -4818 5614 -4816
rect 5668 -4818 5674 -4764
rect 5608 -4824 5674 -4818
rect 5744 -4890 5784 -4526
rect 5174 -4934 5784 -4890
rect 2552 -4936 5784 -4934
rect 5880 -4936 6036 -3918
rect 9140 -4152 9146 -4052
rect 9246 -4152 11462 -4052
rect 11562 -4152 11568 -4052
rect 12260 -4066 13840 -3630
rect 1920 -5026 6036 -4936
rect 1626 -5036 6036 -5026
rect 2300 -5042 6036 -5036
rect 8880 -4310 25158 -4298
rect 8880 -4316 12112 -4310
rect 15250 -4316 25158 -4310
rect 4108 -5044 4226 -5042
rect 1936 -5104 6036 -5102
rect 1936 -5116 6416 -5104
rect 1936 -5122 3952 -5116
rect 1936 -5154 2048 -5122
rect 2454 -5154 3952 -5122
rect 1936 -6772 1990 -5154
rect 2476 -5174 3952 -5154
rect 2476 -5848 2586 -5174
rect 2706 -5276 3952 -5174
rect 2706 -5428 2730 -5276
rect 2964 -5342 3464 -5338
rect 2814 -5348 3606 -5342
rect 2814 -5382 2826 -5348
rect 3594 -5382 3606 -5348
rect 2814 -5388 3606 -5382
rect 2706 -5441 2804 -5428
rect 2706 -5617 2764 -5441
rect 2798 -5617 2804 -5441
rect 2706 -5630 2804 -5617
rect 2964 -5438 3464 -5388
rect 2964 -5618 3020 -5438
rect 3400 -5618 3464 -5438
rect 2706 -5778 2730 -5630
rect 2964 -5670 3464 -5618
rect 3612 -5430 3812 -5420
rect 3612 -5630 3622 -5430
rect 3802 -5630 3812 -5430
rect 3612 -5640 3812 -5630
rect 2814 -5676 3606 -5670
rect 2814 -5710 2826 -5676
rect 3594 -5710 3606 -5676
rect 2814 -5716 3606 -5710
rect 2964 -5718 3464 -5716
rect 3872 -5778 3952 -5276
rect 2706 -5812 3952 -5778
rect 2706 -5848 3714 -5812
rect 2476 -5886 3714 -5848
rect 2476 -6386 2550 -5886
rect 2814 -5952 3606 -5946
rect 2814 -5986 2826 -5952
rect 3594 -5986 3606 -5952
rect 2814 -5992 3606 -5986
rect 2610 -6032 2810 -6022
rect 2610 -6232 2620 -6032
rect 2800 -6232 2810 -6032
rect 2610 -6242 2810 -6232
rect 2962 -6042 3462 -5992
rect 3690 -6032 3714 -5886
rect 2962 -6222 3022 -6042
rect 3402 -6222 3462 -6042
rect 2962 -6274 3462 -6222
rect 3616 -6045 3714 -6032
rect 3616 -6221 3622 -6045
rect 3656 -6221 3714 -6045
rect 3616 -6234 3714 -6221
rect 2814 -6280 3606 -6274
rect 2814 -6314 2826 -6280
rect 3594 -6314 3606 -6280
rect 2814 -6320 3606 -6314
rect 2962 -6326 3462 -6320
rect 3690 -6386 3714 -6234
rect 2476 -6486 3714 -6386
rect 3834 -6486 3952 -5812
rect 2476 -6772 3952 -6486
rect 1936 -6798 2048 -6772
rect 2454 -6798 3952 -6772
rect 1936 -6808 3952 -6798
rect 4374 -5156 6416 -5116
rect 4374 -5174 5838 -5156
rect 4374 -5276 5630 -5174
rect 4374 -5778 4464 -5276
rect 4872 -5342 5372 -5338
rect 4730 -5348 5522 -5342
rect 4730 -5382 4742 -5348
rect 5510 -5382 5522 -5348
rect 4730 -5388 5522 -5382
rect 4524 -5430 4724 -5420
rect 4524 -5630 4534 -5430
rect 4714 -5630 4724 -5430
rect 4524 -5640 4724 -5630
rect 4872 -5438 5372 -5388
rect 5606 -5428 5630 -5276
rect 4872 -5618 4936 -5438
rect 5316 -5618 5372 -5438
rect 4872 -5670 5372 -5618
rect 5532 -5441 5630 -5428
rect 5532 -5617 5538 -5441
rect 5572 -5617 5630 -5441
rect 5532 -5630 5630 -5617
rect 4730 -5676 5522 -5670
rect 4730 -5710 4742 -5676
rect 5510 -5710 5522 -5676
rect 4730 -5716 5522 -5710
rect 4872 -5718 5372 -5716
rect 5606 -5778 5630 -5630
rect 4374 -5812 5630 -5778
rect 4374 -6486 4502 -5812
rect 4622 -5848 5630 -5812
rect 5750 -5848 5838 -5174
rect 4622 -5886 5838 -5848
rect 4622 -6032 4646 -5886
rect 4730 -5952 5522 -5946
rect 4730 -5986 4742 -5952
rect 5510 -5986 5522 -5952
rect 4730 -5992 5522 -5986
rect 4622 -6045 4720 -6032
rect 4622 -6221 4680 -6045
rect 4714 -6221 4720 -6045
rect 4622 -6234 4720 -6221
rect 4874 -6042 5374 -5992
rect 4874 -6222 4934 -6042
rect 5314 -6222 5374 -6042
rect 4622 -6386 4646 -6234
rect 4874 -6274 5374 -6222
rect 5526 -6032 5726 -6022
rect 5526 -6232 5536 -6032
rect 5716 -6232 5726 -6032
rect 5526 -6242 5726 -6232
rect 4730 -6280 5522 -6274
rect 4730 -6314 4742 -6280
rect 5510 -6314 5522 -6280
rect 4730 -6320 5522 -6314
rect 4874 -6326 5374 -6320
rect 5786 -6386 5838 -5886
rect 4622 -6486 5838 -6386
rect 4374 -6774 5838 -6486
rect 6324 -6774 6416 -5156
rect 8880 -5476 8900 -4316
rect 11694 -4574 12058 -4548
rect 11694 -4734 11724 -4574
rect 10476 -4768 11724 -4734
rect 11772 -4626 11980 -4616
rect 10476 -4958 10494 -4768
rect 11772 -4810 11780 -4626
rect 11972 -4810 11980 -4626
rect 12034 -4750 12058 -4574
rect 16094 -4556 16958 -4548
rect 17330 -4556 18192 -4548
rect 16094 -4574 18192 -4556
rect 12034 -4760 12112 -4750
rect 15250 -4760 15282 -4750
rect 12034 -4768 15282 -4760
rect 11772 -4816 11980 -4810
rect 10662 -4886 15100 -4816
rect 10662 -4920 10674 -4886
rect 11042 -4896 11252 -4886
rect 11042 -4920 11054 -4896
rect 10662 -4926 11054 -4920
rect 11240 -4920 11252 -4896
rect 11620 -4920 11830 -4886
rect 12198 -4896 12408 -4886
rect 12198 -4920 12210 -4896
rect 11240 -4926 12210 -4920
rect 12396 -4920 12408 -4896
rect 12776 -4896 12986 -4886
rect 12776 -4920 12844 -4896
rect 12396 -4926 12844 -4920
rect 12974 -4920 12986 -4896
rect 13354 -4896 13564 -4886
rect 13354 -4920 13366 -4896
rect 12974 -4926 13366 -4920
rect 13552 -4920 13564 -4896
rect 13932 -4920 14142 -4886
rect 14510 -4896 14720 -4886
rect 14510 -4920 14522 -4896
rect 13552 -4926 14522 -4920
rect 14708 -4920 14720 -4896
rect 15088 -4920 15100 -4886
rect 14708 -4926 15100 -4920
rect 11436 -4958 12014 -4926
rect 12592 -4958 12844 -4926
rect 13748 -4958 14326 -4926
rect 15264 -4958 15282 -4768
rect 10476 -4970 11230 -4958
rect 11224 -5346 11230 -4970
rect 10462 -5358 11230 -5346
rect 11436 -5354 11452 -4958
rect 11992 -5354 12014 -4958
rect 10462 -5476 10494 -5358
rect 11436 -5390 12014 -5354
rect 12104 -4970 12504 -4958
rect 12104 -5346 12122 -4970
rect 12488 -5346 12504 -4970
rect 12104 -5358 12504 -5346
rect 12592 -5358 12604 -4958
rect 12826 -5358 12844 -4958
rect 12918 -4970 13178 -4958
rect 12918 -5346 12924 -4970
rect 13168 -5346 13178 -4970
rect 12918 -5358 13178 -5346
rect 13260 -4970 13660 -4958
rect 13260 -5346 13276 -4970
rect 13642 -5346 13660 -4970
rect 13260 -5358 13660 -5346
rect 13748 -5354 13768 -4958
rect 14308 -5354 14326 -4958
rect 12592 -5390 12844 -5358
rect 13748 -5390 14326 -5354
rect 14532 -4970 15282 -4958
rect 14532 -5346 14538 -4970
rect 14532 -5358 15282 -5346
rect 8880 -5494 10494 -5476
rect 10662 -5396 11054 -5390
rect 10662 -5430 10674 -5396
rect 11042 -5420 11054 -5396
rect 11240 -5396 12210 -5390
rect 11240 -5420 11252 -5396
rect 11042 -5430 11252 -5420
rect 11620 -5430 11830 -5396
rect 12198 -5420 12210 -5396
rect 12396 -5396 12844 -5390
rect 12396 -5420 12408 -5396
rect 12198 -5430 12408 -5420
rect 12776 -5420 12844 -5396
rect 12974 -5396 13366 -5390
rect 12974 -5420 12986 -5396
rect 12776 -5430 12986 -5420
rect 13354 -5420 13366 -5396
rect 13552 -5396 14522 -5390
rect 13552 -5420 13564 -5396
rect 13354 -5430 13564 -5420
rect 13932 -5430 14142 -5396
rect 14510 -5420 14522 -5396
rect 14708 -5396 15100 -5390
rect 14708 -5420 14720 -5396
rect 14510 -5430 14720 -5420
rect 15088 -5430 15100 -5396
rect 10662 -5500 15100 -5430
rect 15264 -5530 15282 -5358
rect 16094 -5530 16118 -4574
rect 16260 -4660 17076 -4640
rect 16260 -4666 17077 -4660
rect 16260 -4700 16313 -4666
rect 16607 -4700 16771 -4666
rect 17065 -4700 17077 -4666
rect 16301 -4706 16619 -4700
rect 16648 -4706 17077 -4700
rect 16648 -4744 16924 -4706
rect 17106 -4734 17186 -4574
rect 17218 -4660 18034 -4640
rect 17217 -4666 18034 -4660
rect 17217 -4700 17229 -4666
rect 17523 -4700 17687 -4666
rect 17981 -4700 18034 -4666
rect 17217 -4706 17535 -4700
rect 17675 -4706 17993 -4700
rect 16648 -4776 16666 -4744
rect 16210 -4794 16666 -4776
rect 16210 -5484 16228 -4794
rect 16210 -5502 16666 -5484
rect 15264 -5548 16118 -5530
rect 16648 -5530 16666 -5502
rect 16878 -5530 16924 -4744
rect 16648 -5570 16924 -5530
rect 17026 -4750 17266 -4734
rect 17026 -5526 17044 -4750
rect 17246 -5526 17266 -4750
rect 17026 -5542 17266 -5526
rect 17328 -5570 17424 -4706
rect 17498 -4742 18082 -4734
rect 17498 -5530 17508 -4742
rect 17702 -4750 18082 -4742
rect 18064 -5526 18082 -4750
rect 18002 -5530 18082 -5526
rect 17498 -5542 18082 -5530
rect 16301 -5576 16619 -5570
rect 4374 -6808 6416 -6774
rect 1936 -6822 6416 -6808
rect 3364 -7116 3370 -6962
rect 2496 -7126 3370 -7116
rect 2496 -7214 2510 -7126
rect 3230 -7214 3370 -7126
rect 2496 -7222 3370 -7214
rect 3478 -7222 3484 -6962
rect 3614 -7214 3620 -6954
rect 3728 -7110 3734 -6954
rect 3728 -7120 4600 -7110
rect 3728 -7208 3888 -7120
rect 4588 -7208 4600 -7120
rect 3728 -7214 4600 -7208
rect 2406 -8054 2412 -7254
rect 2520 -8054 2526 -7254
rect 2564 -8054 2570 -7254
rect 2678 -8054 2684 -7254
rect 2722 -8054 2728 -7254
rect 2836 -8054 2842 -7254
rect 2880 -8054 2886 -7254
rect 2994 -8054 3000 -7254
rect 3036 -8054 3042 -7254
rect 3150 -8054 3156 -7254
rect 3196 -8054 3202 -7254
rect 3310 -8054 3316 -7254
rect 3364 -8078 3370 -7906
rect 3478 -8078 3484 -7906
rect 3364 -8086 3484 -8078
rect 2496 -8092 3484 -8086
rect 2496 -8172 2512 -8092
rect 3212 -8172 3484 -8092
rect 2496 -8184 3484 -8172
rect 3614 -8078 3620 -7916
rect 3728 -8078 3734 -7916
rect 3782 -8054 3790 -7254
rect 3894 -8054 3902 -7254
rect 3940 -8054 3946 -7254
rect 4054 -8054 4060 -7254
rect 4098 -8054 4104 -7254
rect 4212 -8054 4218 -7254
rect 4256 -8054 4262 -7254
rect 4370 -8054 4376 -7254
rect 4414 -8054 4420 -7254
rect 4528 -8054 4534 -7254
rect 4572 -8054 4578 -7254
rect 4686 -8054 4692 -7254
rect 7588 -7438 7604 -5608
rect 8962 -5636 16060 -5608
rect 16301 -5610 16313 -5576
rect 16607 -5610 16619 -5576
rect 16301 -5616 16619 -5610
rect 16648 -5576 17077 -5570
rect 17217 -5576 17535 -5570
rect 16648 -5610 16771 -5576
rect 17065 -5610 17229 -5576
rect 17523 -5610 17535 -5576
rect 16648 -5616 17535 -5610
rect 8962 -5640 15260 -5636
rect 15938 -5752 16060 -5636
rect 16648 -5636 17534 -5616
rect 15938 -5758 16614 -5752
rect 10492 -5814 15260 -5776
rect 10492 -5988 10580 -5814
rect 10682 -5908 15086 -5888
rect 10682 -5942 10735 -5908
rect 11029 -5942 11307 -5908
rect 11601 -5942 11879 -5908
rect 12173 -5942 12451 -5908
rect 12745 -5942 13023 -5908
rect 13317 -5942 13595 -5908
rect 13889 -5942 14167 -5908
rect 14461 -5942 14739 -5908
rect 15033 -5942 15086 -5908
rect 10682 -5948 15086 -5942
rect 10492 -6000 11248 -5988
rect 11242 -6378 11248 -6000
rect 10492 -6388 11248 -6378
rect 10492 -6390 10680 -6388
rect 10492 -6516 10580 -6390
rect 10723 -6436 11041 -6430
rect 10723 -6470 10735 -6436
rect 11029 -6470 11041 -6436
rect 10723 -6476 11041 -6470
rect 10492 -6518 10680 -6516
rect 11088 -6518 11248 -6388
rect 11362 -6430 11542 -5948
rect 11588 -5990 11892 -5984
rect 11588 -6000 11666 -5990
rect 11814 -6000 11892 -5990
rect 11588 -6378 11602 -6000
rect 11878 -6378 11892 -6000
rect 11588 -6388 11666 -6378
rect 11814 -6388 11892 -6378
rect 11588 -6394 11892 -6388
rect 11295 -6436 11613 -6430
rect 11295 -6470 11307 -6436
rect 11601 -6470 11613 -6436
rect 11295 -6476 11613 -6470
rect 10492 -6528 11248 -6518
rect 11242 -6906 11248 -6528
rect 10492 -6918 11248 -6906
rect 10492 -7086 10580 -6918
rect 10723 -6964 11041 -6958
rect 10723 -6998 10735 -6964
rect 11029 -6998 11041 -6964
rect 10723 -7004 11041 -6998
rect 11088 -7056 11248 -6918
rect 11362 -6958 11542 -6476
rect 11660 -6512 11820 -6394
rect 11936 -6430 12116 -5948
rect 12912 -5982 13260 -5948
rect 12164 -5988 12468 -5984
rect 12164 -6000 12850 -5988
rect 12164 -6378 12176 -6000
rect 12452 -6378 12850 -6000
rect 12164 -6394 12850 -6378
rect 11867 -6436 12185 -6430
rect 11867 -6470 11879 -6436
rect 12173 -6470 12185 -6436
rect 11867 -6476 12185 -6470
rect 11586 -6518 11890 -6512
rect 11586 -6528 11666 -6518
rect 11814 -6528 11890 -6518
rect 11586 -6906 11602 -6528
rect 11878 -6906 11890 -6528
rect 11586 -6916 11666 -6906
rect 11814 -6916 11890 -6906
rect 11586 -6922 11890 -6916
rect 11936 -6958 12116 -6476
rect 12234 -6512 12394 -6394
rect 12912 -6430 12924 -5982
rect 13252 -6392 13260 -5982
rect 12439 -6436 12924 -6430
rect 13250 -6430 13260 -6392
rect 13300 -6000 13604 -5984
rect 13300 -6378 13316 -6000
rect 13592 -6378 13604 -6000
rect 13300 -6394 13604 -6378
rect 13250 -6436 13329 -6430
rect 12439 -6470 12451 -6436
rect 12745 -6468 12924 -6436
rect 12745 -6470 13023 -6468
rect 13317 -6470 13329 -6436
rect 12439 -6476 13329 -6470
rect 12160 -6528 12464 -6512
rect 12160 -6530 12238 -6528
rect 12388 -6530 12464 -6528
rect 12160 -6908 12174 -6530
rect 12450 -6908 12464 -6530
rect 12160 -6922 12464 -6908
rect 11294 -6964 12185 -6958
rect 11294 -6998 11307 -6964
rect 11601 -6998 11879 -6964
rect 12173 -6998 12185 -6964
rect 11294 -7004 12185 -6998
rect 11294 -7018 12184 -7004
rect 12234 -7056 12394 -6922
rect 12508 -6958 12688 -6476
rect 12730 -6518 13034 -6512
rect 12730 -6528 12810 -6518
rect 12958 -6528 13034 -6518
rect 12730 -6906 12742 -6528
rect 13018 -6906 13034 -6528
rect 12730 -6916 12810 -6906
rect 12958 -6916 13034 -6906
rect 12730 -6922 13034 -6916
rect 13080 -6958 13260 -6476
rect 13376 -6512 13536 -6394
rect 13650 -6430 13830 -5948
rect 13874 -5990 14178 -5984
rect 13874 -6000 13954 -5990
rect 14102 -6000 14178 -5990
rect 13874 -6378 13886 -6000
rect 14162 -6378 14178 -6000
rect 13874 -6388 13954 -6378
rect 14102 -6388 14178 -6378
rect 13874 -6394 14178 -6388
rect 13583 -6436 13901 -6430
rect 13583 -6470 13595 -6436
rect 13889 -6470 13901 -6436
rect 13583 -6476 13901 -6470
rect 13304 -6528 13608 -6512
rect 13304 -6906 13316 -6528
rect 13592 -6906 13608 -6528
rect 13304 -6922 13608 -6906
rect 12439 -6964 13330 -6958
rect 12439 -6998 12451 -6964
rect 12745 -6998 13023 -6964
rect 13317 -6998 13330 -6964
rect 12439 -7004 13330 -6998
rect 12440 -7018 13330 -7004
rect 13376 -7056 13536 -6922
rect 13650 -6958 13830 -6476
rect 13948 -6512 14108 -6394
rect 14222 -6430 14402 -5948
rect 15228 -5988 15260 -5814
rect 16602 -5888 16614 -5758
rect 14520 -6000 15260 -5988
rect 15938 -5894 16614 -5888
rect 14520 -6378 14526 -6000
rect 14520 -6388 15260 -6378
rect 14155 -6436 14473 -6430
rect 14155 -6470 14167 -6436
rect 14461 -6470 14473 -6436
rect 14155 -6476 14473 -6470
rect 13876 -6518 14180 -6512
rect 13876 -6528 13954 -6518
rect 14102 -6528 14180 -6518
rect 13876 -6906 13888 -6528
rect 14164 -6906 14180 -6528
rect 13876 -6916 13954 -6906
rect 14102 -6916 14180 -6906
rect 13876 -6922 14180 -6916
rect 14222 -6958 14402 -6476
rect 14520 -6518 14680 -6388
rect 14727 -6436 15045 -6430
rect 14727 -6470 14739 -6436
rect 15033 -6470 15045 -6436
rect 14727 -6476 15045 -6470
rect 15228 -6518 15260 -6388
rect 14520 -6528 15260 -6518
rect 14520 -6906 14526 -6528
rect 14520 -6918 15260 -6906
rect 13583 -6964 14474 -6958
rect 13583 -6998 13595 -6964
rect 13889 -6998 14167 -6964
rect 14461 -6998 14474 -6964
rect 13583 -7004 14474 -6998
rect 13584 -7018 14474 -7004
rect 14520 -7056 14680 -6918
rect 14727 -6964 15045 -6958
rect 14727 -6998 14739 -6964
rect 15033 -6998 15045 -6964
rect 14727 -7004 15045 -6998
rect 11088 -7086 14680 -7056
rect 15228 -7086 15260 -6918
rect 10492 -7114 15260 -7086
rect 15938 -7086 15964 -5894
rect 16036 -5960 16620 -5950
rect 16036 -6050 16162 -5960
rect 16608 -6050 16620 -5960
rect 16036 -6056 16620 -6050
rect 16036 -6554 16156 -6056
rect 16648 -6092 16728 -5636
rect 16762 -5762 17524 -5752
rect 16762 -5888 16776 -5762
rect 17510 -5888 17524 -5762
rect 16762 -5894 17524 -5888
rect 16758 -5956 17078 -5950
rect 16758 -6050 16770 -5956
rect 17066 -6050 17078 -5956
rect 16758 -6056 17078 -6050
rect 17216 -5956 17536 -5950
rect 17216 -6050 17228 -5956
rect 17524 -6050 17536 -5956
rect 17216 -6056 17536 -6050
rect 16036 -7036 16044 -6554
rect 16148 -6938 16156 -6554
rect 16208 -6108 16770 -6092
rect 16208 -6886 16224 -6108
rect 16758 -6886 16770 -6108
rect 16208 -6902 16770 -6886
rect 16830 -6938 16954 -6056
rect 16998 -6106 17298 -6092
rect 16998 -6890 17014 -6106
rect 17280 -6890 17298 -6106
rect 16998 -6902 17298 -6890
rect 17340 -6938 17464 -6056
rect 17564 -6092 17644 -5542
rect 17675 -5576 17993 -5570
rect 17675 -5610 17687 -5576
rect 17981 -5610 17993 -5576
rect 17675 -5616 17993 -5610
rect 18174 -5674 18192 -4574
rect 21246 -5244 22086 -5218
rect 21246 -5274 21272 -5244
rect 18848 -5382 20732 -5352
rect 18848 -5530 18878 -5382
rect 18952 -5462 20544 -5456
rect 18952 -5496 18964 -5462
rect 20532 -5496 20544 -5462
rect 18952 -5502 19090 -5496
rect 18848 -5534 18900 -5530
rect 18848 -5546 18942 -5534
rect 18848 -5548 18902 -5546
rect 18862 -5622 18902 -5548
rect 18936 -5622 18942 -5546
rect 18862 -5634 18942 -5622
rect 18174 -5694 18808 -5674
rect 17684 -5762 18742 -5752
rect 17684 -5886 17700 -5762
rect 18728 -5850 18742 -5762
rect 18788 -5790 18808 -5694
rect 18862 -5790 18900 -5634
rect 19036 -5666 19090 -5502
rect 18952 -5672 19090 -5666
rect 19230 -5502 20544 -5496
rect 19230 -5666 20470 -5502
rect 20574 -5534 20674 -5530
rect 20554 -5546 20674 -5534
rect 20554 -5622 20560 -5546
rect 20594 -5622 20674 -5546
rect 20554 -5634 20674 -5622
rect 19230 -5672 20544 -5666
rect 18952 -5706 18964 -5672
rect 20532 -5706 20544 -5672
rect 18952 -5712 20544 -5706
rect 18788 -5808 18900 -5790
rect 18728 -5864 20528 -5850
rect 17684 -5894 18330 -5886
rect 17674 -5960 18258 -5950
rect 17674 -6050 17686 -5960
rect 18132 -6050 18258 -5960
rect 17674 -6056 18258 -6050
rect 17520 -6100 18082 -6092
rect 17520 -6894 17528 -6100
rect 17782 -6108 18082 -6100
rect 18066 -6886 18082 -6108
rect 17782 -6894 18082 -6886
rect 17520 -6902 18082 -6894
rect 18138 -6554 18258 -6056
rect 18138 -6938 18146 -6554
rect 16148 -6944 17118 -6938
rect 16148 -7034 16162 -6944
rect 17078 -7034 17118 -6944
rect 16148 -7036 17118 -7034
rect 16036 -7044 17118 -7036
rect 16160 -7046 17118 -7044
rect 17176 -6944 18146 -6938
rect 17176 -7034 17216 -6944
rect 18132 -7034 18146 -6944
rect 17176 -7036 18146 -7034
rect 18250 -7036 18258 -6554
rect 17176 -7046 18258 -7036
rect 18304 -7086 18330 -5894
rect 20504 -6354 20528 -5864
rect 18834 -6382 20528 -6354
rect 20574 -6016 20674 -5634
rect 20714 -5776 20732 -5382
rect 21246 -5402 21270 -5274
rect 21433 -5334 21591 -5328
rect 21433 -5368 21445 -5334
rect 21579 -5368 21591 -5334
rect 21433 -5374 21468 -5368
rect 21246 -5406 21400 -5402
rect 21246 -5418 21406 -5406
rect 21246 -5486 21366 -5418
rect 21214 -5494 21366 -5486
rect 21400 -5494 21406 -5418
rect 21214 -5506 21406 -5494
rect 21214 -5508 21400 -5506
rect 21214 -5776 21232 -5508
rect 21462 -5538 21468 -5374
rect 21433 -5544 21468 -5538
rect 21556 -5374 21591 -5368
rect 21556 -5538 21562 -5374
rect 21620 -5406 21662 -5244
rect 21691 -5334 21849 -5328
rect 21691 -5368 21703 -5334
rect 21837 -5368 21849 -5334
rect 21691 -5374 21849 -5368
rect 21618 -5418 21664 -5406
rect 21618 -5494 21624 -5418
rect 21658 -5494 21664 -5418
rect 21618 -5506 21664 -5494
rect 21556 -5544 21591 -5538
rect 21433 -5578 21445 -5544
rect 21579 -5578 21591 -5544
rect 21433 -5584 21468 -5578
rect 20714 -5790 21232 -5776
rect 21290 -5616 21390 -5610
rect 21290 -5628 21406 -5616
rect 21290 -5704 21366 -5628
rect 21400 -5704 21406 -5628
rect 21290 -5716 21406 -5704
rect 20574 -6104 20580 -6016
rect 20668 -6104 20674 -6016
rect 18834 -6547 18898 -6382
rect 18932 -6466 20524 -6460
rect 18932 -6500 18944 -6466
rect 20512 -6500 20524 -6466
rect 18932 -6506 19092 -6500
rect 18834 -6559 18922 -6547
rect 18834 -6635 18882 -6559
rect 18916 -6635 18922 -6559
rect 18834 -6647 18922 -6635
rect 18834 -6816 18898 -6647
rect 19036 -6688 19092 -6506
rect 18932 -6694 19092 -6688
rect 19232 -6506 20524 -6500
rect 19232 -6688 20460 -6506
rect 20574 -6547 20674 -6104
rect 20534 -6559 20674 -6547
rect 20534 -6635 20540 -6559
rect 20574 -6635 20674 -6559
rect 20534 -6647 20674 -6635
rect 20574 -6654 20674 -6647
rect 20712 -5870 21212 -5850
rect 19232 -6694 20524 -6688
rect 18932 -6728 18944 -6694
rect 20512 -6728 20524 -6694
rect 18932 -6734 20524 -6728
rect 20712 -6816 20736 -5870
rect 21184 -6560 21212 -5870
rect 21290 -6010 21390 -5716
rect 21462 -5748 21468 -5584
rect 21433 -5754 21468 -5748
rect 21556 -5584 21591 -5578
rect 21556 -5748 21562 -5584
rect 21620 -5616 21662 -5506
rect 21718 -5538 21818 -5374
rect 21876 -5418 22000 -5406
rect 21876 -5494 21882 -5418
rect 21916 -5494 22000 -5418
rect 21876 -5506 22000 -5494
rect 21691 -5544 21849 -5538
rect 21691 -5578 21703 -5544
rect 21837 -5578 21849 -5544
rect 21691 -5584 21849 -5578
rect 21618 -5628 21664 -5616
rect 21618 -5704 21624 -5628
rect 21658 -5704 21664 -5628
rect 21618 -5716 21664 -5704
rect 21718 -5748 21818 -5584
rect 21900 -5616 22000 -5506
rect 21876 -5628 22000 -5616
rect 21876 -5704 21882 -5628
rect 21916 -5704 22000 -5628
rect 21876 -5716 22000 -5704
rect 21556 -5754 21591 -5748
rect 21433 -5788 21445 -5754
rect 21579 -5788 21591 -5754
rect 21433 -5794 21591 -5788
rect 21691 -5754 21849 -5748
rect 21691 -5788 21703 -5754
rect 21837 -5788 21849 -5754
rect 21691 -5794 21849 -5788
rect 21718 -6010 21818 -5794
rect 21290 -6110 21818 -6010
rect 21290 -6411 21390 -6110
rect 21718 -6324 21818 -6110
rect 21900 -5990 22000 -5716
rect 22066 -5852 22086 -5244
rect 23274 -5322 23778 -5298
rect 23274 -5406 23294 -5322
rect 23376 -5402 23642 -5322
rect 23376 -5404 23446 -5402
rect 22816 -5422 23294 -5406
rect 22816 -5758 22836 -5422
rect 23434 -5436 23446 -5404
rect 23572 -5404 23642 -5402
rect 23724 -5404 23778 -5322
rect 23572 -5436 23584 -5404
rect 23434 -5442 23584 -5436
rect 23356 -5464 23402 -5452
rect 23356 -5494 23362 -5464
rect 22638 -5776 22836 -5758
rect 22914 -5594 23362 -5494
rect 22638 -5852 22654 -5776
rect 22914 -5842 23014 -5594
rect 23356 -5632 23362 -5594
rect 23396 -5494 23402 -5464
rect 23616 -5464 23662 -5452
rect 23616 -5494 23622 -5464
rect 23396 -5594 23622 -5494
rect 23396 -5632 23402 -5594
rect 23356 -5644 23402 -5632
rect 23616 -5632 23622 -5594
rect 23656 -5494 23662 -5464
rect 23656 -5594 23666 -5494
rect 23656 -5632 23662 -5594
rect 23616 -5644 23662 -5632
rect 22066 -5872 22654 -5852
rect 22714 -5852 23014 -5842
rect 22374 -5948 22652 -5924
rect 21900 -5996 22308 -5990
rect 21900 -6124 22006 -5996
rect 22302 -6124 22308 -5996
rect 21900 -6130 22308 -6124
rect 21433 -6330 21591 -6324
rect 21433 -6364 21445 -6330
rect 21579 -6364 21591 -6330
rect 21433 -6370 21470 -6364
rect 21290 -6423 21406 -6411
rect 21290 -6499 21366 -6423
rect 21400 -6499 21406 -6423
rect 21290 -6511 21406 -6499
rect 21290 -6516 21390 -6511
rect 21464 -6552 21470 -6370
rect 21433 -6558 21470 -6552
rect 21560 -6370 21591 -6364
rect 21691 -6330 21849 -6324
rect 21691 -6364 21703 -6330
rect 21837 -6364 21849 -6330
rect 21691 -6370 21849 -6364
rect 21560 -6552 21564 -6370
rect 21618 -6423 21664 -6411
rect 21618 -6499 21624 -6423
rect 21658 -6499 21664 -6423
rect 21618 -6511 21664 -6499
rect 21560 -6558 21591 -6552
rect 21184 -6580 21272 -6560
rect 18834 -6844 20736 -6816
rect 21202 -6636 21272 -6580
rect 21433 -6592 21445 -6558
rect 21579 -6592 21591 -6558
rect 21433 -6598 21470 -6592
rect 21202 -6639 21400 -6636
rect 21202 -6651 21406 -6639
rect 21202 -6727 21366 -6651
rect 21400 -6727 21406 -6651
rect 21202 -6739 21406 -6727
rect 21202 -6742 21400 -6739
rect 21202 -6878 21272 -6742
rect 21464 -6780 21470 -6598
rect 21433 -6786 21470 -6780
rect 21560 -6598 21591 -6592
rect 21560 -6780 21564 -6598
rect 21620 -6639 21662 -6511
rect 21718 -6552 21818 -6370
rect 21900 -6411 22000 -6130
rect 22374 -6188 22398 -5948
rect 21876 -6423 22000 -6411
rect 21876 -6499 21882 -6423
rect 21916 -6499 22000 -6423
rect 21876 -6511 22000 -6499
rect 21691 -6558 21849 -6552
rect 21691 -6592 21703 -6558
rect 21837 -6592 21849 -6558
rect 21691 -6598 21849 -6592
rect 21618 -6651 21664 -6639
rect 21618 -6727 21624 -6651
rect 21658 -6727 21664 -6651
rect 21618 -6739 21664 -6727
rect 21560 -6786 21591 -6780
rect 21433 -6820 21445 -6786
rect 21579 -6820 21591 -6786
rect 21433 -6826 21591 -6820
rect 21202 -6902 21274 -6878
rect 21620 -6902 21662 -6739
rect 21718 -6780 21818 -6598
rect 21900 -6639 22000 -6511
rect 21876 -6651 22000 -6639
rect 21876 -6727 21882 -6651
rect 21916 -6727 22000 -6651
rect 21876 -6738 22000 -6727
rect 22070 -6224 22398 -6188
rect 21876 -6739 21922 -6738
rect 21691 -6786 21849 -6780
rect 21691 -6820 21703 -6786
rect 21837 -6820 21849 -6786
rect 21691 -6826 21849 -6820
rect 21718 -6828 21818 -6826
rect 22070 -6902 22118 -6224
rect 22620 -6674 22652 -5948
rect 22714 -6132 22726 -5852
rect 23002 -6132 23014 -5852
rect 22714 -6142 23014 -6132
rect 23434 -5660 23584 -5654
rect 23434 -5694 23446 -5660
rect 23572 -5694 23584 -5660
rect 23434 -5930 23584 -5694
rect 23756 -5834 23778 -5404
rect 25134 -5834 25158 -4316
rect 23756 -5858 25158 -5834
rect 24010 -5930 24210 -5924
rect 23434 -6130 24010 -5930
rect 22714 -6496 22814 -6142
rect 23434 -6398 23584 -6130
rect 24010 -6136 24210 -6130
rect 24286 -5946 25202 -5924
rect 24286 -6220 24312 -5946
rect 24082 -6246 24312 -6220
rect 23131 -6404 23931 -6398
rect 23131 -6438 23143 -6404
rect 23919 -6438 23931 -6404
rect 23131 -6444 23931 -6438
rect 23044 -6466 23090 -6454
rect 23044 -6496 23050 -6466
rect 22714 -6596 23050 -6496
rect 23044 -6634 23050 -6596
rect 23084 -6496 23090 -6466
rect 23972 -6466 24018 -6454
rect 23972 -6496 23978 -6466
rect 23084 -6596 23978 -6496
rect 23084 -6634 23090 -6596
rect 23044 -6646 23090 -6634
rect 23972 -6634 23978 -6596
rect 24012 -6634 24018 -6466
rect 23972 -6646 24018 -6634
rect 23131 -6662 23931 -6656
rect 22620 -6694 22982 -6674
rect 22930 -6776 22982 -6694
rect 23131 -6696 23143 -6662
rect 23919 -6696 23931 -6662
rect 24082 -6674 24114 -6246
rect 23131 -6702 23931 -6696
rect 23332 -6774 23730 -6702
rect 24080 -6774 24114 -6674
rect 23332 -6776 24114 -6774
rect 22930 -6802 24114 -6776
rect 25178 -6674 25202 -5946
rect 25178 -6802 25204 -6674
rect 21202 -6930 22118 -6902
rect 15938 -7114 18330 -7086
rect 25180 -7248 25204 -6802
rect 21202 -7250 25204 -7248
rect 10008 -7290 25204 -7250
rect 10008 -7366 10100 -7290
rect 8962 -7410 10100 -7366
rect 8962 -7438 9648 -7410
rect 7588 -7454 9648 -7438
rect 9792 -7434 9902 -7410
rect 9792 -7468 9809 -7434
rect 9885 -7468 9902 -7434
rect 10046 -7454 10100 -7410
rect 24218 -7402 24654 -7390
rect 10618 -7454 11048 -7438
rect 9792 -7474 9902 -7468
rect 9710 -7496 9756 -7484
rect 8920 -7608 9068 -7586
rect 3614 -8096 3734 -8078
rect 3614 -8102 4608 -8096
rect 3614 -8188 3888 -8102
rect 4594 -8188 4608 -8102
rect 3614 -8196 4608 -8188
rect 8920 -10142 8940 -7608
rect 9046 -9422 9068 -7608
rect 9148 -7700 9364 -7684
rect 9148 -7734 9220 -7700
rect 9296 -7734 9364 -7700
rect 9148 -7750 9364 -7734
rect 9130 -7762 9386 -7750
rect 9130 -9330 9136 -7762
rect 9170 -7774 9346 -7762
rect 9170 -9240 9208 -7774
rect 9304 -9240 9346 -7774
rect 9170 -9268 9346 -9240
rect 9170 -9330 9176 -9268
rect 9130 -9342 9176 -9330
rect 9340 -9330 9346 -9268
rect 9380 -8908 9386 -7762
rect 9710 -8908 9716 -7496
rect 9380 -9002 9716 -8908
rect 9380 -9330 9386 -9002
rect 9710 -9064 9716 -9002
rect 9750 -7548 9756 -7496
rect 9938 -7496 9984 -7484
rect 9938 -7548 9944 -7496
rect 9750 -7570 9944 -7548
rect 9750 -9050 9788 -7570
rect 9904 -9050 9944 -7570
rect 9750 -9064 9944 -9050
rect 9978 -8908 9984 -7496
rect 10618 -7492 10638 -7454
rect 11035 -7492 11048 -7454
rect 10618 -7620 11048 -7492
rect 24218 -7540 24230 -7402
rect 24644 -7540 24654 -7402
rect 24218 -7550 24654 -7540
rect 24760 -7404 25152 -7368
rect 10618 -7658 10638 -7620
rect 11035 -7658 11048 -7620
rect 10618 -7674 11048 -7658
rect 24220 -7620 24650 -7604
rect 24220 -7658 24237 -7620
rect 24634 -7658 24650 -7620
rect 10620 -7786 11050 -7770
rect 10620 -7824 10638 -7786
rect 11035 -7824 11050 -7786
rect 10620 -7952 11050 -7824
rect 24220 -7786 24650 -7658
rect 24220 -7824 24237 -7786
rect 24634 -7824 24650 -7786
rect 24220 -7840 24650 -7824
rect 10620 -7990 10638 -7952
rect 11035 -7990 11050 -7952
rect 10620 -8006 11050 -7990
rect 24220 -7952 24650 -7936
rect 24220 -7990 24237 -7952
rect 24634 -7990 24650 -7952
rect 10620 -8118 11050 -8102
rect 10620 -8156 10638 -8118
rect 11035 -8156 11050 -8118
rect 10620 -8284 11050 -8156
rect 24220 -8118 24650 -7990
rect 24220 -8156 24237 -8118
rect 24634 -8156 24650 -8118
rect 24220 -8172 24650 -8156
rect 10620 -8322 10638 -8284
rect 11035 -8322 11050 -8284
rect 10620 -8338 11050 -8322
rect 24220 -8284 24650 -8266
rect 24220 -8322 24237 -8284
rect 24634 -8322 24650 -8284
rect 10620 -8450 11050 -8434
rect 10620 -8488 10638 -8450
rect 11035 -8488 11050 -8450
rect 10620 -8616 11050 -8488
rect 24220 -8450 24650 -8322
rect 24220 -8488 24237 -8450
rect 24634 -8488 24650 -8450
rect 24220 -8502 24650 -8488
rect 10620 -8654 10638 -8616
rect 11035 -8654 11050 -8616
rect 10620 -8670 11050 -8654
rect 24220 -8616 24650 -8598
rect 24220 -8654 24237 -8616
rect 24634 -8654 24650 -8616
rect 10620 -8782 11050 -8766
rect 10620 -8820 10638 -8782
rect 11035 -8820 11050 -8782
rect 9978 -9002 10547 -8908
rect 10620 -8948 11050 -8820
rect 24220 -8782 24650 -8654
rect 24220 -8820 24237 -8782
rect 24634 -8820 24650 -8782
rect 24220 -8834 24650 -8820
rect 10620 -8986 10638 -8948
rect 11035 -8986 11050 -8948
rect 10620 -9002 11050 -8986
rect 24220 -8948 24650 -8930
rect 24220 -8986 24237 -8948
rect 24634 -8986 24650 -8948
rect 9978 -9064 9984 -9002
rect 9710 -9076 9984 -9064
rect 9736 -9092 9952 -9076
rect 9736 -9126 9809 -9092
rect 9885 -9126 9952 -9092
rect 9736 -9132 9952 -9126
rect 10146 -9088 10384 -9066
rect 9340 -9342 9386 -9330
rect 9208 -9358 9308 -9352
rect 9208 -9392 9220 -9358
rect 9296 -9392 9308 -9358
rect 10146 -9386 10162 -9088
rect 9208 -9422 9308 -9392
rect 9448 -9406 10162 -9386
rect 9448 -9408 9636 -9406
rect 10048 -9408 10162 -9406
rect 9448 -9422 9466 -9408
rect 9046 -9442 9466 -9422
rect 10362 -9940 10384 -9088
rect 10453 -9751 10547 -9002
rect 10620 -9114 11050 -9098
rect 10620 -9152 10638 -9114
rect 11035 -9152 11050 -9114
rect 10620 -9280 11050 -9152
rect 24220 -9114 24650 -8986
rect 24220 -9152 24237 -9114
rect 24634 -9152 24650 -9114
rect 24220 -9166 24650 -9152
rect 10620 -9318 10638 -9280
rect 11035 -9318 11050 -9280
rect 10620 -9334 11050 -9318
rect 24220 -9280 24650 -9264
rect 24220 -9318 24237 -9280
rect 24634 -9318 24650 -9280
rect 10620 -9446 11050 -9428
rect 10620 -9484 10638 -9446
rect 11035 -9484 11050 -9446
rect 10620 -9612 11050 -9484
rect 24220 -9446 24650 -9318
rect 24220 -9484 24237 -9446
rect 24634 -9484 24650 -9446
rect 24220 -9500 24650 -9484
rect 10620 -9650 10638 -9612
rect 11035 -9650 11050 -9612
rect 10620 -9664 11050 -9650
rect 24220 -9612 24650 -9596
rect 24220 -9650 24237 -9612
rect 24634 -9650 24650 -9612
rect 10453 -9778 11069 -9751
rect 10453 -9816 10638 -9778
rect 11035 -9816 11069 -9778
rect 10453 -9845 11069 -9816
rect 24220 -9778 24650 -9650
rect 24220 -9816 24237 -9778
rect 24634 -9816 24650 -9778
rect 24220 -9832 24650 -9816
rect 24760 -9940 24788 -7404
rect 10362 -9960 24788 -9940
rect 25116 -10142 25152 -7404
rect 8920 -10144 24792 -10142
rect 25112 -10144 25152 -10142
rect 8920 -10176 25152 -10144
rect 15968 -10464 25450 -10450
rect 15968 -11130 15988 -10464
rect 16648 -10898 17142 -10464
rect 18052 -10898 25450 -10464
rect 16648 -11130 25450 -10898
rect 15968 -11150 25450 -11130
rect 1844 -11310 21916 -11292
rect 1844 -11314 17714 -11310
rect 1844 -11824 2030 -11314
rect 3298 -11484 17714 -11314
rect 3298 -11798 15036 -11484
rect 15812 -11798 17714 -11484
rect 18284 -11798 21916 -11310
rect 3298 -11824 7814 -11798
rect 1844 -13814 1996 -11824
rect 7070 -12022 7814 -11824
rect 7070 -12862 7118 -12022
rect 7752 -12034 7814 -12022
rect 7752 -12082 13436 -12034
rect 7330 -12178 7522 -12172
rect 7330 -12212 7342 -12178
rect 7510 -12212 7522 -12178
rect 7330 -12218 7522 -12212
rect 13404 -12194 13436 -12082
rect 7274 -12262 7320 -12250
rect 7274 -12438 7280 -12262
rect 7314 -12438 7320 -12262
rect 7274 -12450 7320 -12438
rect 7370 -12482 7478 -12218
rect 13404 -12226 20656 -12194
rect 8272 -12238 9864 -12232
rect 7532 -12260 7578 -12250
rect 7532 -12262 7714 -12260
rect 7532 -12438 7538 -12262
rect 7572 -12270 7714 -12262
rect 7704 -12430 7714 -12270
rect 8272 -12272 8284 -12238
rect 9852 -12264 9864 -12238
rect 9930 -12238 11522 -12232
rect 9852 -12272 9886 -12264
rect 8272 -12278 9886 -12272
rect 9930 -12272 9942 -12238
rect 11510 -12272 11522 -12238
rect 9930 -12278 9998 -12272
rect 8336 -12310 9886 -12278
rect 8216 -12322 8262 -12310
rect 8216 -12382 8222 -12322
rect 8256 -12382 8262 -12322
rect 8216 -12394 8262 -12382
rect 8336 -12322 9920 -12310
rect 8336 -12382 8348 -12322
rect 9840 -12382 9880 -12322
rect 9914 -12382 9920 -12322
rect 8336 -12394 9920 -12382
rect 8336 -12426 9886 -12394
rect 9978 -12426 9998 -12278
rect 7572 -12438 7714 -12430
rect 7532 -12440 7714 -12438
rect 8272 -12432 9886 -12426
rect 7532 -12450 7578 -12440
rect 8272 -12466 8284 -12432
rect 9852 -12442 9886 -12432
rect 9930 -12432 9998 -12426
rect 11440 -12278 11522 -12272
rect 11588 -12238 13180 -12232
rect 11588 -12272 11600 -12238
rect 13168 -12272 13180 -12238
rect 11588 -12278 11662 -12272
rect 11440 -12426 11464 -12278
rect 11532 -12322 11578 -12310
rect 11532 -12382 11538 -12322
rect 11572 -12382 11578 -12322
rect 11532 -12394 11578 -12382
rect 11640 -12426 11662 -12278
rect 11440 -12432 11522 -12426
rect 9852 -12466 9864 -12442
rect 8272 -12472 9864 -12466
rect 9930 -12466 9942 -12432
rect 11510 -12466 11522 -12432
rect 9930 -12472 11522 -12466
rect 11588 -12432 11662 -12426
rect 13104 -12278 13180 -12272
rect 13104 -12426 13126 -12278
rect 20278 -12298 20478 -12284
rect 20278 -12302 20292 -12298
rect 13236 -12306 20292 -12302
rect 13190 -12322 20292 -12306
rect 13190 -12382 13196 -12322
rect 13230 -12382 20292 -12322
rect 13190 -12398 20292 -12382
rect 13236 -12402 20292 -12398
rect 13104 -12432 13180 -12426
rect 11588 -12466 11600 -12432
rect 13168 -12466 13180 -12432
rect 11588 -12472 13180 -12466
rect 20278 -12468 20292 -12402
rect 20464 -12468 20478 -12298
rect 7330 -12488 7522 -12482
rect 7330 -12522 7342 -12488
rect 7510 -12522 7522 -12488
rect 7330 -12528 7522 -12522
rect 13404 -12510 20194 -12474
rect 20278 -12484 20478 -12468
rect 2982 -12938 7118 -12862
rect 7339 -12620 7514 -12528
rect 13404 -12618 13436 -12510
rect 7339 -12910 7346 -12620
rect 7506 -12910 7514 -12620
rect 7339 -12916 7514 -12910
rect 7744 -12680 13436 -12618
rect 20150 -12618 20194 -12510
rect 20610 -12618 20656 -12226
rect 20150 -12646 20656 -12618
rect 21870 -12646 21916 -11798
rect 22120 -11596 25450 -11150
rect 22120 -11668 25512 -11596
rect 22120 -12538 22152 -11668
rect 25426 -11672 25512 -11668
rect 22120 -12574 24616 -12538
rect 7744 -12898 7778 -12680
rect 20150 -12752 21916 -12646
rect 19808 -12799 21916 -12752
rect 2982 -12958 3152 -12938
rect 2982 -13448 3002 -12958
rect 3140 -12976 3152 -12958
rect 3549 -12958 7118 -12938
rect 7744 -12938 19070 -12898
rect 7744 -12954 18551 -12938
rect 3549 -12976 3561 -12958
rect 3140 -12982 3561 -12976
rect 3134 -13104 3566 -13098
rect 3134 -13142 3152 -13104
rect 3549 -13142 3566 -13104
rect 3134 -13270 3566 -13142
rect 3134 -13308 3152 -13270
rect 3549 -13308 3566 -13270
rect 3134 -13314 3566 -13308
rect 3140 -13436 3561 -13430
rect 3140 -13448 3152 -13436
rect 2982 -13474 3152 -13448
rect 3549 -13448 3561 -13436
rect 4022 -13448 4422 -12958
rect 6016 -13448 6416 -12958
rect 8000 -13448 8400 -12954
rect 10006 -13448 10406 -12954
rect 12016 -13448 12416 -12954
rect 14008 -13448 14408 -12954
rect 16002 -13448 16402 -12954
rect 18008 -12976 18551 -12954
rect 18948 -12976 19070 -12938
rect 18008 -13098 19070 -12976
rect 19808 -13093 19926 -12799
rect 19960 -13093 20836 -12799
rect 20870 -13093 21746 -12799
rect 21780 -13093 21916 -12799
rect 19808 -13098 21916 -13093
rect 18008 -13104 21916 -13098
rect 18008 -13112 18551 -13104
rect 18008 -13448 18408 -13112
rect 18539 -13142 18551 -13112
rect 18948 -13112 21916 -13104
rect 22452 -12795 22556 -12794
rect 23444 -12795 23486 -12794
rect 24374 -12795 24416 -12794
rect 22452 -12807 22560 -12795
rect 22452 -13101 22520 -12807
rect 22554 -12834 22560 -12807
rect 23442 -12807 23488 -12795
rect 23442 -12834 23448 -12807
rect 22554 -13028 23448 -12834
rect 22554 -13101 22560 -13028
rect 18948 -13142 18960 -13112
rect 18539 -13148 18960 -13142
rect 22452 -13113 22560 -13101
rect 22596 -13092 23404 -13078
rect 18532 -13242 21712 -13228
rect 18532 -13244 20918 -13242
rect 18532 -13270 20008 -13244
rect 18532 -13308 18551 -13270
rect 18948 -13308 20008 -13270
rect 18532 -13322 20008 -13308
rect 18532 -13350 19822 -13322
rect 19460 -13368 19822 -13350
rect 19994 -13352 20008 -13322
rect 20788 -13330 20918 -13244
rect 20788 -13352 20802 -13330
rect 18539 -13436 18960 -13430
rect 18539 -13448 18551 -13436
rect 3549 -13474 18551 -13448
rect 18948 -13448 18960 -13436
rect 18948 -13474 19350 -13448
rect 2982 -13538 19350 -13474
rect 19328 -13814 19350 -13538
rect 1844 -13870 19350 -13814
rect 1844 -13876 19358 -13870
rect 1844 -13892 2150 -13876
rect 1844 -18044 1970 -13892
rect 2138 -13914 2150 -13892
rect 2547 -13888 18949 -13876
rect 2547 -13892 4972 -13888
rect 5450 -13890 18949 -13888
rect 5450 -13892 8958 -13890
rect 9436 -13892 18949 -13890
rect 2547 -13914 2559 -13892
rect 2138 -13920 2559 -13914
rect 2138 -14038 2559 -14036
rect 2132 -14042 2564 -14038
rect 2132 -14080 2150 -14042
rect 2547 -14080 2564 -14042
rect 2132 -14208 2564 -14080
rect 2132 -14246 2150 -14208
rect 2547 -14246 2564 -14208
rect 2132 -14254 2564 -14246
rect 2134 -14374 2566 -14368
rect 2134 -14412 2150 -14374
rect 2547 -14412 2566 -14374
rect 2134 -14540 2566 -14412
rect 2134 -14578 2150 -14540
rect 2547 -14578 2566 -14540
rect 2134 -14584 2566 -14578
rect 2132 -14706 2564 -14700
rect 2132 -14744 2150 -14706
rect 2547 -14744 2564 -14706
rect 2132 -14872 2564 -14744
rect 2132 -14910 2150 -14872
rect 2547 -14910 2564 -14872
rect 2132 -14916 2564 -14910
rect 2132 -15038 2564 -15032
rect 2132 -15076 2150 -15038
rect 2547 -15076 2564 -15038
rect 2132 -15204 2564 -15076
rect 2132 -15242 2150 -15204
rect 2547 -15242 2564 -15204
rect 2132 -15248 2564 -15242
rect 2130 -15370 2562 -15362
rect 2130 -15408 2150 -15370
rect 2547 -15408 2562 -15370
rect 2130 -15536 2562 -15408
rect 2130 -15574 2150 -15536
rect 2547 -15574 2562 -15536
rect 2130 -15578 2562 -15574
rect 2138 -15580 2559 -15578
rect 2132 -15702 2564 -15696
rect 2132 -15740 2150 -15702
rect 2547 -15740 2564 -15702
rect 2132 -15868 2564 -15740
rect 2132 -15906 2150 -15868
rect 2547 -15906 2564 -15868
rect 2132 -15912 2564 -15906
rect 2132 -16034 2564 -16026
rect 2132 -16072 2150 -16034
rect 2547 -16072 2564 -16034
rect 2132 -16200 2564 -16072
rect 2132 -16238 2150 -16200
rect 2547 -16238 2564 -16200
rect 2132 -16242 2564 -16238
rect 2138 -16244 2559 -16242
rect 2132 -16366 2564 -16360
rect 2132 -16404 2150 -16366
rect 2547 -16404 2564 -16366
rect 2132 -16532 2564 -16404
rect 2132 -16570 2150 -16532
rect 2547 -16570 2564 -16532
rect 2132 -16576 2564 -16570
rect 2130 -16698 2562 -16692
rect 2130 -16736 2150 -16698
rect 2547 -16736 2562 -16698
rect 2130 -16864 2562 -16736
rect 2130 -16902 2150 -16864
rect 2547 -16902 2562 -16864
rect 2130 -16908 2562 -16902
rect 2130 -17030 2562 -17024
rect 2130 -17068 2150 -17030
rect 2547 -17068 2562 -17030
rect 2130 -17196 2562 -17068
rect 2130 -17234 2150 -17196
rect 2547 -17234 2562 -17196
rect 2130 -17240 2562 -17234
rect 2132 -17362 2564 -17354
rect 2132 -17400 2150 -17362
rect 2547 -17400 2564 -17362
rect 2132 -17528 2564 -17400
rect 2132 -17566 2150 -17528
rect 2547 -17566 2564 -17528
rect 2132 -17570 2564 -17566
rect 2138 -17572 2559 -17570
rect 2132 -17694 2564 -17688
rect 2132 -17732 2150 -17694
rect 2547 -17732 2564 -17694
rect 2132 -17860 2564 -17732
rect 2132 -17898 2150 -17860
rect 2547 -17898 2564 -17860
rect 2132 -17904 2564 -17898
rect 2138 -18026 2559 -18020
rect 2138 -18044 2150 -18026
rect 1844 -18064 2150 -18044
rect 2547 -18044 2559 -18026
rect 5008 -18044 5408 -18040
rect 7024 -18044 7424 -13892
rect 9006 -18044 9406 -18042
rect 11014 -18044 11414 -13892
rect 14994 -18044 15394 -13892
rect 18937 -13914 18949 -13892
rect 19346 -13914 19358 -13876
rect 18937 -13920 19358 -13914
rect 16042 -13978 16556 -13972
rect 16042 -13980 19366 -13978
rect 16042 -14472 16050 -13980
rect 16548 -13994 19366 -13980
rect 16548 -14456 18384 -13994
rect 19346 -14132 19366 -13994
rect 18848 -14146 19366 -14132
rect 18848 -14456 18870 -14146
rect 18932 -14208 19364 -14202
rect 18932 -14246 18949 -14208
rect 19346 -14246 19364 -14208
rect 18932 -14374 19364 -14246
rect 18932 -14412 18949 -14374
rect 19346 -14412 19364 -14374
rect 18932 -14418 19364 -14412
rect 16548 -14466 18870 -14456
rect 16548 -14472 16556 -14466
rect 16042 -14480 16556 -14472
rect 18932 -14540 19364 -14534
rect 18932 -14578 18949 -14540
rect 19346 -14578 19364 -14540
rect 18932 -14706 19364 -14578
rect 18932 -14744 18949 -14706
rect 19346 -14744 19364 -14706
rect 18932 -14750 19364 -14744
rect 19460 -14838 19640 -13368
rect 19920 -13377 19966 -13365
rect 19994 -13368 20802 -13352
rect 20904 -13350 20918 -13330
rect 21698 -13350 21712 -13242
rect 19920 -13426 19926 -13377
rect 19698 -13440 19926 -13426
rect 19698 -14762 19712 -13440
rect 19844 -13626 19926 -13440
rect 19844 -14576 19858 -13626
rect 19920 -13671 19926 -13626
rect 19960 -13426 19966 -13377
rect 20830 -13377 20876 -13365
rect 20904 -13368 21712 -13350
rect 20830 -13426 20836 -13377
rect 19960 -13452 20836 -13426
rect 19960 -13600 19998 -13452
rect 20798 -13600 20836 -13452
rect 19960 -13626 20836 -13600
rect 19960 -13671 19966 -13626
rect 19920 -13683 19966 -13671
rect 20830 -13671 20836 -13626
rect 20870 -13426 20876 -13377
rect 21740 -13377 21786 -13365
rect 21740 -13426 21746 -13377
rect 20870 -13452 21746 -13426
rect 20870 -13600 20908 -13452
rect 21708 -13600 21746 -13452
rect 20870 -13626 21746 -13600
rect 20870 -13671 20876 -13626
rect 19994 -13702 20802 -13680
rect 20830 -13683 20876 -13671
rect 21740 -13671 21746 -13626
rect 21780 -13671 21786 -13377
rect 19994 -13870 20010 -13702
rect 19994 -13896 20204 -13870
rect 19920 -13955 19966 -13943
rect 19920 -14249 19926 -13955
rect 19960 -14249 19966 -13955
rect 19920 -14261 19966 -14249
rect 20174 -14308 20204 -13896
rect 19994 -14336 20204 -14308
rect 19994 -14500 20010 -14336
rect 20786 -13718 20802 -13702
rect 20904 -13700 21712 -13680
rect 21740 -13683 21786 -13671
rect 22452 -13373 22554 -13113
rect 22452 -13385 22560 -13373
rect 22452 -13679 22520 -13385
rect 22554 -13450 22560 -13385
rect 22596 -13392 22608 -13092
rect 23388 -13138 23404 -13092
rect 23442 -13101 23448 -13028
rect 23482 -12836 23488 -12807
rect 24370 -12807 24416 -12795
rect 24370 -12836 24376 -12807
rect 23482 -13028 24376 -12836
rect 23482 -13101 23488 -13028
rect 23442 -13113 23488 -13101
rect 23524 -13090 24332 -13078
rect 23390 -13160 23404 -13138
rect 23524 -13160 23538 -13090
rect 23390 -13326 23538 -13160
rect 23390 -13344 23404 -13326
rect 23388 -13392 23404 -13344
rect 22596 -13402 23404 -13392
rect 23442 -13385 23488 -13373
rect 23442 -13450 23448 -13385
rect 22554 -13618 23448 -13450
rect 22554 -13679 22560 -13618
rect 20904 -13718 20920 -13700
rect 20786 -13800 20920 -13718
rect 21696 -13800 21712 -13700
rect 22452 -13691 22560 -13679
rect 22594 -13668 23402 -13656
rect 21816 -13758 21956 -13746
rect 20786 -13820 21712 -13800
rect 20786 -13870 20802 -13820
rect 21748 -13848 21828 -13758
rect 20622 -13896 20802 -13870
rect 20908 -13856 21828 -13848
rect 20622 -14308 20654 -13896
rect 20830 -13955 20876 -13943
rect 20830 -14249 20836 -13955
rect 20870 -14008 20876 -13955
rect 20908 -13952 20920 -13856
rect 21696 -13874 21828 -13856
rect 21944 -13874 21956 -13758
rect 21696 -13908 21956 -13874
rect 21696 -13952 21708 -13908
rect 20908 -13964 21708 -13952
rect 21740 -13955 21786 -13943
rect 21740 -14008 21746 -13955
rect 20870 -14030 21746 -14008
rect 20870 -14249 20882 -14030
rect 20830 -14261 20882 -14249
rect 20854 -14306 20882 -14261
rect 21736 -14249 21746 -14030
rect 21780 -14170 21786 -13955
rect 22452 -13951 22554 -13691
rect 22452 -13963 22560 -13951
rect 21780 -14249 22400 -14170
rect 21736 -14306 22400 -14249
rect 20854 -14308 20916 -14306
rect 21698 -14308 22400 -14306
rect 20622 -14336 20802 -14308
rect 20854 -14330 22400 -14308
rect 20786 -14384 20802 -14336
rect 20786 -14404 22156 -14384
rect 20786 -14486 20920 -14404
rect 20786 -14500 20802 -14486
rect 19920 -14533 19966 -14521
rect 19994 -14524 20802 -14500
rect 20904 -14504 20920 -14486
rect 21696 -14482 22156 -14404
rect 21696 -14504 21712 -14482
rect 19920 -14576 19926 -14533
rect 19844 -14762 19926 -14576
rect 19698 -14776 19926 -14762
rect 19920 -14827 19926 -14776
rect 19960 -14576 19966 -14533
rect 20830 -14533 20876 -14521
rect 20904 -14524 21712 -14504
rect 20830 -14576 20836 -14533
rect 19960 -14602 20836 -14576
rect 19960 -14750 19998 -14602
rect 20798 -14750 20836 -14602
rect 19960 -14776 20836 -14750
rect 19960 -14827 19966 -14776
rect 18932 -14872 19364 -14866
rect 18932 -14910 18949 -14872
rect 19346 -14910 19364 -14872
rect 18932 -15038 19364 -14910
rect 19460 -14884 19822 -14838
rect 19920 -14839 19966 -14827
rect 20830 -14827 20836 -14776
rect 20870 -14576 20876 -14533
rect 21740 -14533 21786 -14521
rect 21740 -14576 21746 -14533
rect 20870 -14600 21746 -14576
rect 20870 -14748 20908 -14600
rect 21708 -14748 21746 -14600
rect 20870 -14776 21746 -14748
rect 20870 -14827 20876 -14776
rect 19994 -14854 20802 -14838
rect 20830 -14839 20876 -14827
rect 21740 -14827 21746 -14776
rect 21780 -14827 21786 -14533
rect 19994 -14884 20008 -14854
rect 19460 -14962 20008 -14884
rect 20788 -14876 20802 -14854
rect 20904 -14854 21712 -14838
rect 21740 -14839 21786 -14827
rect 20904 -14876 20920 -14854
rect 20788 -14962 20920 -14876
rect 21700 -14962 21712 -14854
rect 19460 -14978 21712 -14962
rect 18932 -15076 18949 -15038
rect 19346 -15076 19364 -15038
rect 18932 -15082 19364 -15076
rect 19920 -15111 19966 -15099
rect 19920 -15122 19926 -15111
rect 18402 -15164 18802 -15148
rect 18402 -15530 18420 -15164
rect 18784 -15530 18802 -15164
rect 18932 -15204 19364 -15198
rect 18932 -15242 18949 -15204
rect 19346 -15242 19364 -15204
rect 18932 -15370 19364 -15242
rect 18932 -15408 18949 -15370
rect 19346 -15408 19364 -15370
rect 18932 -15414 19364 -15408
rect 19502 -15405 19926 -15122
rect 19960 -15122 19966 -15111
rect 20830 -15111 20876 -15099
rect 20830 -15122 20836 -15111
rect 19960 -15405 20836 -15122
rect 20870 -15122 20876 -15111
rect 21740 -15111 21786 -15099
rect 21740 -15122 21746 -15111
rect 20870 -15405 21746 -15122
rect 21780 -15122 21786 -15111
rect 21780 -15405 21878 -15122
rect 18402 -15548 18802 -15530
rect 18932 -15536 19364 -15530
rect 18426 -17798 18776 -15548
rect 18932 -15574 18949 -15536
rect 19346 -15574 19364 -15536
rect 18932 -15702 19364 -15574
rect 18932 -15740 18949 -15702
rect 19346 -15740 19364 -15702
rect 18932 -15746 19364 -15740
rect 19502 -15548 21878 -15405
rect 18932 -15868 19364 -15862
rect 18932 -15906 18949 -15868
rect 19346 -15906 19364 -15868
rect 18932 -16034 19364 -15906
rect 18932 -16072 18949 -16034
rect 19346 -16072 19364 -16034
rect 18932 -16078 19364 -16072
rect 18932 -16200 19364 -16194
rect 18932 -16238 18949 -16200
rect 19346 -16238 19364 -16200
rect 18932 -16366 19364 -16238
rect 18932 -16404 18949 -16366
rect 19346 -16404 19364 -16366
rect 18932 -16410 19364 -16404
rect 18932 -16532 19364 -16526
rect 18932 -16570 18949 -16532
rect 19346 -16570 19364 -16532
rect 18932 -16698 19364 -16570
rect 18932 -16736 18949 -16698
rect 19346 -16736 19364 -16698
rect 18932 -16742 19364 -16736
rect 18932 -16864 19364 -16858
rect 18932 -16902 18949 -16864
rect 19346 -16902 19364 -16864
rect 18932 -17030 19364 -16902
rect 18932 -17068 18949 -17030
rect 19346 -17068 19364 -17030
rect 18932 -17074 19364 -17068
rect 18932 -17196 19364 -17190
rect 18932 -17234 18949 -17196
rect 19346 -17234 19364 -17196
rect 18932 -17362 19364 -17234
rect 18932 -17400 18949 -17362
rect 19346 -17400 19364 -17362
rect 18932 -17406 19364 -17400
rect 18932 -17528 19364 -17522
rect 18932 -17566 18949 -17528
rect 19346 -17566 19364 -17528
rect 18932 -17694 19364 -17566
rect 18932 -17732 18949 -17694
rect 19346 -17732 19364 -17694
rect 18932 -17738 19364 -17732
rect 18426 -17860 19376 -17798
rect 18426 -17898 18949 -17860
rect 19346 -17898 19376 -17860
rect 18426 -17958 19376 -17898
rect 2547 -18064 18352 -18044
rect 1844 -18128 18352 -18064
rect 1844 -18408 1996 -18128
rect 18346 -18408 18352 -18128
rect 1844 -18466 18352 -18408
rect 1844 -18486 2148 -18466
rect 1844 -22670 1970 -18486
rect 2136 -18504 2148 -18486
rect 2545 -18484 18352 -18466
rect 2545 -18486 4962 -18484
rect 5456 -18486 18352 -18484
rect 2545 -18504 2557 -18486
rect 2136 -18510 2557 -18504
rect 2130 -18632 2564 -18616
rect 2130 -18670 2148 -18632
rect 2545 -18670 2564 -18632
rect 2130 -18798 2564 -18670
rect 2130 -18836 2148 -18798
rect 2545 -18836 2564 -18798
rect 2130 -18850 2564 -18836
rect 2130 -18964 2564 -18950
rect 2130 -19002 2148 -18964
rect 2545 -19002 2564 -18964
rect 2130 -19130 2564 -19002
rect 2130 -19168 2148 -19130
rect 2545 -19168 2564 -19130
rect 2130 -19184 2564 -19168
rect 2130 -19296 2564 -19280
rect 2130 -19334 2148 -19296
rect 2545 -19334 2564 -19296
rect 2130 -19462 2564 -19334
rect 2130 -19500 2148 -19462
rect 2545 -19500 2564 -19462
rect 2130 -19514 2564 -19500
rect 2130 -19628 2564 -19612
rect 2130 -19666 2148 -19628
rect 2545 -19666 2564 -19628
rect 2130 -19794 2564 -19666
rect 2130 -19832 2148 -19794
rect 2545 -19832 2564 -19794
rect 2130 -19846 2564 -19832
rect 2130 -19960 2564 -19946
rect 2130 -19998 2148 -19960
rect 2545 -19998 2564 -19960
rect 2130 -20126 2564 -19998
rect 2130 -20164 2148 -20126
rect 2545 -20164 2564 -20126
rect 2130 -20180 2564 -20164
rect 2130 -20292 2564 -20276
rect 2130 -20330 2148 -20292
rect 2545 -20330 2564 -20292
rect 2130 -20458 2564 -20330
rect 2130 -20496 2148 -20458
rect 2545 -20496 2564 -20458
rect 2130 -20510 2564 -20496
rect 2130 -20624 2564 -20608
rect 2130 -20662 2148 -20624
rect 2545 -20662 2564 -20624
rect 2130 -20790 2564 -20662
rect 2130 -20828 2148 -20790
rect 2545 -20828 2564 -20790
rect 2130 -20842 2564 -20828
rect 2128 -20956 2562 -20940
rect 2128 -20994 2148 -20956
rect 2545 -20994 2562 -20956
rect 2128 -21122 2562 -20994
rect 2128 -21160 2148 -21122
rect 2545 -21160 2562 -21122
rect 2128 -21174 2562 -21160
rect 2130 -21288 2564 -21272
rect 2130 -21326 2148 -21288
rect 2545 -21326 2564 -21288
rect 2130 -21454 2564 -21326
rect 2130 -21492 2148 -21454
rect 2545 -21492 2564 -21454
rect 2130 -21506 2564 -21492
rect 2130 -21620 2564 -21604
rect 2130 -21658 2148 -21620
rect 2545 -21658 2564 -21620
rect 2130 -21786 2564 -21658
rect 2130 -21824 2148 -21786
rect 2545 -21824 2564 -21786
rect 2130 -21838 2564 -21824
rect 2128 -21952 2562 -21936
rect 2128 -21990 2148 -21952
rect 2545 -21990 2562 -21952
rect 2128 -22118 2562 -21990
rect 2128 -22156 2148 -22118
rect 2545 -22156 2562 -22118
rect 2128 -22170 2562 -22156
rect 2136 -22232 2670 -22222
rect 2136 -22372 2148 -22232
rect 2654 -22372 2670 -22232
rect 2136 -22382 2670 -22372
rect 2136 -22450 2557 -22444
rect 2136 -22488 2148 -22450
rect 2545 -22488 2557 -22450
rect 2136 -22494 2557 -22488
rect 5008 -22670 5408 -22668
rect 9006 -22670 9406 -18486
rect 13040 -22670 13440 -18486
rect 16960 -22670 17360 -18486
rect 18426 -18578 18776 -17958
rect 18937 -18026 19358 -18020
rect 18937 -18044 18949 -18026
rect 18850 -18064 18949 -18044
rect 19346 -18044 19358 -18026
rect 19502 -18044 19534 -15548
rect 20220 -15918 21532 -15878
rect 20220 -15994 20252 -15918
rect 20220 -16020 20254 -15994
rect 20222 -17992 20254 -16020
rect 20464 -16008 21264 -15994
rect 19346 -18064 19534 -18044
rect 18850 -18128 19534 -18064
rect 20220 -18022 20254 -17992
rect 20332 -16106 20432 -16094
rect 20332 -16174 20392 -16106
rect 20426 -16174 20432 -16106
rect 20332 -16264 20432 -16174
rect 20332 -16332 20392 -16264
rect 20426 -16332 20432 -16264
rect 20464 -16268 20474 -16008
rect 21252 -16268 21264 -16008
rect 20464 -16284 21264 -16268
rect 21296 -16106 21396 -16094
rect 21296 -16174 21302 -16106
rect 21336 -16174 21396 -16106
rect 21296 -16264 21396 -16174
rect 20332 -16422 20432 -16332
rect 20332 -16490 20392 -16422
rect 20426 -16490 20432 -16422
rect 20464 -16324 21264 -16312
rect 20464 -16430 20474 -16324
rect 21252 -16430 21264 -16324
rect 20464 -16442 21264 -16430
rect 21296 -16332 21302 -16264
rect 21336 -16332 21396 -16264
rect 21520 -16254 21532 -15918
rect 21862 -16254 21878 -15548
rect 21956 -15590 22156 -14482
rect 22240 -14884 22400 -14330
rect 22452 -14257 22520 -13963
rect 22554 -14022 22560 -13963
rect 22594 -13968 22610 -13668
rect 23390 -13702 23402 -13668
rect 23442 -13679 23448 -13618
rect 23482 -13450 23488 -13385
rect 23524 -13390 23538 -13326
rect 24318 -13160 24332 -13090
rect 24370 -13101 24376 -13028
rect 24410 -13101 24416 -12807
rect 24370 -13113 24416 -13101
rect 24548 -13160 24616 -12574
rect 24318 -13326 24616 -13160
rect 24318 -13390 24332 -13326
rect 23524 -13402 24332 -13390
rect 24370 -13374 24416 -13373
rect 24370 -13385 24478 -13374
rect 24370 -13450 24376 -13385
rect 23482 -13618 24376 -13450
rect 23482 -13679 23488 -13618
rect 23442 -13691 23488 -13679
rect 23520 -13666 24328 -13656
rect 23390 -13738 23404 -13702
rect 23520 -13738 23536 -13666
rect 24316 -13702 24328 -13666
rect 24370 -13679 24376 -13618
rect 24410 -13679 24478 -13385
rect 24370 -13691 24478 -13679
rect 24316 -13714 24330 -13702
rect 23390 -13904 23536 -13738
rect 23390 -13942 23404 -13904
rect 23390 -13968 23402 -13942
rect 22594 -13980 23402 -13968
rect 23442 -13963 23488 -13951
rect 23442 -14022 23448 -13963
rect 22554 -14190 23448 -14022
rect 22554 -14257 22560 -14190
rect 22452 -14269 22560 -14257
rect 22596 -14242 23404 -14230
rect 22452 -14529 22554 -14269
rect 22452 -14541 22560 -14529
rect 22452 -14834 22520 -14541
rect 22514 -14835 22520 -14834
rect 22554 -14598 22560 -14541
rect 22596 -14542 22608 -14242
rect 23388 -14298 23404 -14242
rect 23442 -14257 23448 -14190
rect 23482 -14022 23488 -13963
rect 23520 -13966 23536 -13904
rect 24318 -13922 24330 -13714
rect 24316 -13942 24330 -13922
rect 24316 -13966 24328 -13942
rect 24376 -13951 24478 -13691
rect 23520 -13980 24328 -13966
rect 24370 -13963 24478 -13951
rect 24370 -14022 24376 -13963
rect 23482 -14190 24376 -14022
rect 23482 -14257 23488 -14190
rect 23442 -14269 23488 -14257
rect 23524 -14238 24332 -14230
rect 23390 -14316 23404 -14298
rect 23524 -14316 23538 -14238
rect 23390 -14482 23538 -14316
rect 23390 -14504 23404 -14482
rect 23388 -14542 23404 -14504
rect 22596 -14554 23404 -14542
rect 23442 -14541 23488 -14529
rect 23442 -14598 23448 -14541
rect 22554 -14766 23448 -14598
rect 22554 -14835 22560 -14766
rect 22514 -14847 22560 -14835
rect 22596 -14814 23404 -14802
rect 22596 -14884 22610 -14814
rect 22240 -14976 22610 -14884
rect 23390 -14976 23404 -14814
rect 23442 -14835 23448 -14766
rect 23482 -14598 23488 -14541
rect 23524 -14538 23538 -14482
rect 24318 -14316 24332 -14238
rect 24370 -14257 24376 -14190
rect 24410 -14257 24478 -13963
rect 24370 -14268 24478 -14257
rect 24370 -14269 24416 -14268
rect 24548 -14316 24616 -13326
rect 24318 -14482 24616 -14316
rect 24318 -14538 24332 -14482
rect 23524 -14554 24332 -14538
rect 24370 -14532 24416 -14529
rect 24370 -14541 24478 -14532
rect 24370 -14598 24376 -14541
rect 23482 -14766 24376 -14598
rect 23482 -14835 23488 -14766
rect 23442 -14847 23488 -14835
rect 24370 -14835 24376 -14766
rect 24410 -14835 24478 -14541
rect 24370 -14847 24478 -14835
rect 22240 -14982 23404 -14976
rect 23552 -14908 24300 -14894
rect 22452 -15107 22554 -15040
rect 22452 -15119 22560 -15107
rect 22452 -15413 22520 -15119
rect 22554 -15184 22560 -15119
rect 23442 -15119 23488 -15107
rect 23442 -15184 23448 -15119
rect 22554 -15352 23448 -15184
rect 22554 -15413 22560 -15352
rect 22452 -15425 22560 -15413
rect 23442 -15413 23448 -15352
rect 23482 -15413 23488 -15119
rect 23442 -15425 23488 -15413
rect 22452 -15560 22554 -15425
rect 22452 -15590 23486 -15560
rect 21956 -15598 23486 -15590
rect 21956 -15642 22612 -15598
rect 23390 -15642 23486 -15598
rect 23552 -15622 23570 -14908
rect 24284 -15622 24300 -14908
rect 24376 -15107 24478 -14847
rect 24370 -15119 24478 -15107
rect 24370 -15413 24376 -15119
rect 24410 -15413 24478 -15119
rect 24370 -15425 24478 -15413
rect 23552 -15638 24300 -15622
rect 21956 -15697 22610 -15642
rect 21956 -15750 22520 -15697
rect 21520 -16266 21878 -16254
rect 22452 -15991 22520 -15750
rect 22554 -15914 22610 -15697
rect 23392 -15685 23486 -15642
rect 24376 -15685 24478 -15425
rect 23392 -15697 23488 -15685
rect 23392 -15914 23448 -15697
rect 22554 -15946 23448 -15914
rect 22554 -15991 22560 -15946
rect 22452 -16003 22560 -15991
rect 22596 -15988 23404 -15978
rect 22452 -16263 22554 -16003
rect 21296 -16422 21396 -16332
rect 20332 -16580 20432 -16490
rect 20332 -16648 20392 -16580
rect 20426 -16648 20432 -16580
rect 20464 -16482 21264 -16470
rect 20464 -16588 20474 -16482
rect 21252 -16588 21264 -16482
rect 20464 -16600 21264 -16588
rect 21296 -16490 21302 -16422
rect 21336 -16490 21396 -16422
rect 21296 -16580 21396 -16490
rect 22452 -16275 22560 -16263
rect 22452 -16569 22520 -16275
rect 22554 -16332 22560 -16275
rect 22596 -16288 22610 -15988
rect 23390 -16050 23404 -15988
rect 23442 -15991 23448 -15946
rect 23482 -15752 23488 -15697
rect 24370 -15697 24478 -15685
rect 24370 -15752 24376 -15697
rect 23482 -15920 24376 -15752
rect 23482 -15991 23488 -15920
rect 23442 -16003 23488 -15991
rect 23522 -15988 24330 -15978
rect 23522 -16050 23538 -15988
rect 23390 -16216 23538 -16050
rect 23390 -16288 23404 -16216
rect 22596 -16302 23404 -16288
rect 23442 -16275 23488 -16263
rect 23442 -16332 23448 -16275
rect 22554 -16500 23448 -16332
rect 22554 -16569 22560 -16500
rect 20332 -16738 20432 -16648
rect 20332 -16806 20392 -16738
rect 20426 -16806 20432 -16738
rect 20464 -16640 21264 -16628
rect 20464 -16746 20474 -16640
rect 21252 -16746 21264 -16640
rect 20464 -16758 21264 -16746
rect 21296 -16648 21302 -16580
rect 21336 -16648 21396 -16580
rect 21296 -16738 21396 -16648
rect 20332 -16896 20432 -16806
rect 20332 -16964 20392 -16896
rect 20426 -16964 20432 -16896
rect 20464 -16798 21264 -16786
rect 20464 -16904 20474 -16798
rect 21252 -16904 21264 -16798
rect 20464 -16916 21264 -16904
rect 21296 -16806 21302 -16738
rect 21336 -16806 21396 -16738
rect 21296 -16896 21396 -16806
rect 20332 -17054 20432 -16964
rect 20332 -17122 20392 -17054
rect 20426 -17122 20432 -17054
rect 20464 -16956 21264 -16944
rect 20464 -17062 20474 -16956
rect 21252 -17062 21264 -16956
rect 20464 -17074 21264 -17062
rect 21296 -16964 21302 -16896
rect 21336 -16964 21396 -16896
rect 21296 -17054 21396 -16964
rect 20332 -17212 20432 -17122
rect 20332 -17280 20392 -17212
rect 20426 -17280 20432 -17212
rect 20464 -17114 21264 -17102
rect 20464 -17220 20476 -17114
rect 21254 -17220 21264 -17114
rect 20464 -17232 21264 -17220
rect 21296 -17122 21302 -17054
rect 21336 -17122 21396 -17054
rect 21704 -16590 22104 -16576
rect 21704 -17098 21718 -16590
rect 22090 -17098 22104 -16590
rect 21704 -17112 22104 -17098
rect 22452 -16581 22560 -16569
rect 22596 -16552 23404 -16540
rect 22452 -16841 22554 -16581
rect 22452 -16853 22560 -16841
rect 21296 -17212 21396 -17122
rect 20332 -17370 20432 -17280
rect 20332 -17438 20392 -17370
rect 20426 -17438 20432 -17370
rect 20464 -17272 21264 -17260
rect 20464 -17378 20474 -17272
rect 21252 -17378 21264 -17272
rect 20464 -17390 21264 -17378
rect 21296 -17280 21302 -17212
rect 21336 -17280 21396 -17212
rect 21296 -17370 21396 -17280
rect 20332 -17528 20432 -17438
rect 20332 -17596 20392 -17528
rect 20426 -17596 20432 -17528
rect 20464 -17430 21264 -17418
rect 20464 -17536 20474 -17430
rect 21252 -17536 21264 -17430
rect 20464 -17548 21264 -17536
rect 21296 -17438 21302 -17370
rect 21336 -17438 21396 -17370
rect 21296 -17528 21396 -17438
rect 20332 -17686 20432 -17596
rect 20332 -17754 20392 -17686
rect 20426 -17754 20432 -17686
rect 20464 -17588 21264 -17576
rect 20464 -17694 20474 -17588
rect 21252 -17694 21264 -17588
rect 20464 -17706 21264 -17694
rect 21296 -17596 21302 -17528
rect 21336 -17596 21396 -17528
rect 21296 -17686 21396 -17596
rect 20332 -17844 20432 -17754
rect 20332 -17912 20392 -17844
rect 20426 -17912 20432 -17844
rect 18850 -18408 18856 -18128
rect 18850 -18466 19534 -18408
rect 20220 -18466 20252 -18022
rect 20332 -18116 20432 -17912
rect 20464 -17750 21264 -17734
rect 20464 -17756 20476 -17750
rect 21250 -17756 21264 -17750
rect 20464 -17996 20472 -17756
rect 20464 -18010 20474 -17996
rect 21252 -18010 21264 -17756
rect 20464 -18022 21264 -18010
rect 21296 -17754 21302 -17686
rect 21336 -17754 21396 -17686
rect 21296 -17844 21396 -17754
rect 21296 -17912 21302 -17844
rect 21336 -17912 21396 -17844
rect 21296 -18116 21396 -17912
rect 20332 -18216 21396 -18116
rect 18850 -18486 20252 -18466
rect 17754 -18590 19608 -18578
rect 17754 -19030 17768 -18590
rect 19592 -19030 19608 -18590
rect 17754 -19040 19608 -19030
rect 19848 -22670 20248 -18486
rect 20776 -20592 20936 -18216
rect 21830 -18388 21990 -17112
rect 22452 -17147 22520 -16853
rect 22554 -16906 22560 -16853
rect 22596 -16852 22610 -16552
rect 23390 -16628 23404 -16552
rect 23442 -16569 23448 -16500
rect 23482 -16332 23488 -16275
rect 23522 -16288 23538 -16216
rect 24318 -16050 24330 -15988
rect 24370 -15991 24376 -15920
rect 24410 -15991 24478 -15697
rect 24370 -16000 24478 -15991
rect 24370 -16003 24416 -16000
rect 24548 -16050 24616 -14482
rect 24318 -16216 24616 -16050
rect 24318 -16288 24330 -16216
rect 23522 -16302 24330 -16288
rect 24370 -16264 24416 -16263
rect 24370 -16275 24478 -16264
rect 24370 -16332 24376 -16275
rect 23482 -16500 24376 -16332
rect 23482 -16569 23488 -16500
rect 23442 -16581 23488 -16569
rect 23524 -16552 24332 -16540
rect 23524 -16628 23536 -16552
rect 24316 -16604 24332 -16552
rect 24370 -16569 24376 -16500
rect 24410 -16569 24478 -16275
rect 24370 -16581 24478 -16569
rect 23390 -16794 23536 -16628
rect 23390 -16852 23404 -16794
rect 22596 -16864 23404 -16852
rect 23442 -16853 23488 -16841
rect 23442 -16906 23448 -16853
rect 22554 -17074 23448 -16906
rect 22554 -17147 22560 -17074
rect 22452 -17159 22560 -17147
rect 22596 -17138 23404 -17126
rect 22452 -17419 22554 -17159
rect 22452 -17431 22560 -17419
rect 22452 -17725 22520 -17431
rect 22554 -17502 22560 -17431
rect 22596 -17438 22610 -17138
rect 23390 -17206 23404 -17138
rect 23442 -17147 23448 -17074
rect 23482 -16906 23488 -16853
rect 23524 -16852 23536 -16794
rect 24318 -16812 24332 -16604
rect 24316 -16852 24332 -16812
rect 24376 -16841 24478 -16581
rect 23524 -16864 24332 -16852
rect 24370 -16853 24478 -16841
rect 24370 -16906 24376 -16853
rect 23482 -17074 24376 -16906
rect 23482 -17147 23488 -17074
rect 23442 -17159 23488 -17147
rect 23524 -17136 24332 -17126
rect 23524 -17206 23538 -17136
rect 23390 -17372 23538 -17206
rect 23390 -17438 23404 -17372
rect 22596 -17450 23404 -17438
rect 23442 -17431 23488 -17419
rect 23442 -17502 23448 -17431
rect 22554 -17696 23448 -17502
rect 22554 -17725 22560 -17696
rect 22452 -17736 22560 -17725
rect 22514 -17737 22560 -17736
rect 23442 -17725 23448 -17696
rect 23482 -17502 23488 -17431
rect 23524 -17436 23538 -17372
rect 24318 -17206 24332 -17136
rect 24370 -17147 24376 -17074
rect 24410 -17147 24478 -16853
rect 24370 -17158 24478 -17147
rect 24370 -17159 24416 -17158
rect 24548 -17206 24616 -16216
rect 24318 -17372 24616 -17206
rect 24318 -17436 24332 -17372
rect 23524 -17450 24332 -17436
rect 24370 -17431 24416 -17419
rect 24370 -17502 24376 -17431
rect 23482 -17694 24376 -17502
rect 23482 -17725 23488 -17694
rect 23442 -17737 23488 -17725
rect 24370 -17725 24376 -17694
rect 24410 -17725 24416 -17431
rect 24370 -17737 24416 -17725
rect 24548 -17820 24616 -17372
rect 22120 -17924 24616 -17820
rect 25428 -17924 25512 -11672
rect 22120 -17984 25512 -17924
rect 24548 -17986 25512 -17984
rect 21830 -18548 23334 -18388
rect 24535 -18466 24956 -18460
rect 24535 -18504 24547 -18466
rect 24944 -18504 24956 -18466
rect 24535 -18510 24956 -18504
rect 23174 -18572 23334 -18548
rect 23174 -18632 24982 -18572
rect 23174 -18670 24547 -18632
rect 24944 -18670 24982 -18632
rect 23174 -18732 24982 -18670
rect 23174 -19970 23334 -18732
rect 24530 -18798 24964 -18782
rect 24530 -18836 24547 -18798
rect 24944 -18836 24964 -18798
rect 24530 -18964 24964 -18836
rect 24530 -19002 24547 -18964
rect 24944 -19002 24964 -18964
rect 24530 -19016 24964 -19002
rect 24530 -19130 24964 -19114
rect 24530 -19168 24547 -19130
rect 24944 -19168 24964 -19130
rect 24530 -19296 24964 -19168
rect 24530 -19334 24547 -19296
rect 24944 -19334 24964 -19296
rect 24530 -19348 24964 -19334
rect 24530 -19462 24964 -19446
rect 24530 -19500 24547 -19462
rect 24944 -19500 24964 -19462
rect 24530 -19628 24964 -19500
rect 24530 -19666 24547 -19628
rect 24944 -19666 24964 -19628
rect 24530 -19680 24964 -19666
rect 24530 -19794 24964 -19778
rect 24530 -19832 24547 -19794
rect 24944 -19832 24964 -19794
rect 24530 -19960 24964 -19832
rect 23102 -19984 23402 -19970
rect 23102 -20260 23114 -19984
rect 23386 -20260 23402 -19984
rect 24530 -19998 24547 -19960
rect 24944 -19998 24964 -19960
rect 24530 -20012 24964 -19998
rect 23102 -20270 23402 -20260
rect 24530 -20126 24964 -20110
rect 24530 -20164 24547 -20126
rect 24944 -20164 24964 -20126
rect 20704 -20606 21004 -20592
rect 20704 -20882 20718 -20606
rect 20990 -20882 21004 -20606
rect 20704 -20892 21004 -20882
rect 20776 -22154 20936 -20892
rect 20706 -22168 21006 -22154
rect 20706 -22440 20720 -22168
rect 20992 -22440 21006 -22168
rect 20706 -22454 21006 -22440
rect 1844 -22710 20318 -22670
rect 1844 -23440 1890 -22710
rect 20268 -23440 20318 -22710
rect 20776 -22932 20936 -22454
rect 21474 -22828 22674 -22792
rect 20458 -22942 21408 -22932
rect 20458 -22952 21328 -22942
rect 20458 -23018 20472 -22952
rect 20538 -23008 21328 -22952
rect 21394 -23008 21408 -22942
rect 20538 -23018 21408 -23008
rect 20458 -23032 21408 -23018
rect 20776 -23304 20936 -23032
rect 21474 -23088 21482 -22828
rect 21214 -23096 21482 -23088
rect 21544 -22830 22674 -22828
rect 21544 -23090 22604 -22830
rect 21214 -23158 21226 -23096
rect 21544 -23158 21764 -23090
rect 21214 -23186 21764 -23158
rect 1844 -23486 20318 -23440
rect 20656 -23312 21056 -23304
rect 20656 -23696 20664 -23312
rect 21048 -23696 21056 -23312
rect 21288 -23598 21764 -23186
rect 22366 -23160 22604 -23090
rect 22666 -23090 22674 -22830
rect 23174 -22932 23334 -20270
rect 24530 -20292 24964 -20164
rect 24530 -20330 24547 -20292
rect 24944 -20330 24964 -20292
rect 24530 -20344 24964 -20330
rect 24530 -20458 24964 -20442
rect 24530 -20496 24547 -20458
rect 24944 -20496 24964 -20458
rect 24530 -20624 24964 -20496
rect 24530 -20662 24547 -20624
rect 24944 -20662 24964 -20624
rect 24530 -20676 24964 -20662
rect 24530 -20790 24964 -20774
rect 24530 -20828 24547 -20790
rect 24944 -20828 24964 -20790
rect 24530 -20956 24964 -20828
rect 24530 -20994 24547 -20956
rect 24944 -20994 24964 -20956
rect 24530 -21008 24964 -20994
rect 24528 -21122 24962 -21108
rect 24528 -21160 24547 -21122
rect 24944 -21160 24962 -21122
rect 24528 -21288 24962 -21160
rect 24528 -21326 24547 -21288
rect 24944 -21326 24962 -21288
rect 24528 -21342 24962 -21326
rect 24530 -21454 24964 -21438
rect 24530 -21492 24547 -21454
rect 24944 -21492 24964 -21454
rect 24530 -21620 24964 -21492
rect 24530 -21658 24547 -21620
rect 24944 -21658 24964 -21620
rect 24530 -21672 24964 -21658
rect 24528 -21786 24962 -21770
rect 24528 -21824 24547 -21786
rect 24944 -21824 24962 -21786
rect 24528 -21952 24962 -21824
rect 24528 -21990 24547 -21952
rect 24944 -21990 24962 -21952
rect 24528 -22004 24962 -21990
rect 24528 -22118 24962 -22104
rect 24528 -22156 24547 -22118
rect 24944 -22156 24962 -22118
rect 24528 -22284 24962 -22156
rect 24528 -22322 24547 -22284
rect 24944 -22322 24962 -22284
rect 24528 -22338 24962 -22322
rect 24535 -22450 24956 -22444
rect 24535 -22488 24547 -22450
rect 24944 -22488 24956 -22450
rect 24535 -22494 24956 -22488
rect 25198 -22706 25512 -17986
rect 24040 -22730 25512 -22706
rect 22740 -22944 23658 -22932
rect 22740 -23010 22754 -22944
rect 22820 -22954 23658 -22944
rect 22820 -23010 23580 -22954
rect 22740 -23020 23580 -23010
rect 23646 -23020 23658 -22954
rect 22740 -23032 23658 -23020
rect 22666 -23098 22934 -23090
rect 22922 -23160 22934 -23098
rect 22366 -23348 22934 -23160
rect 23174 -23304 23334 -23032
rect 24040 -23206 24070 -22730
rect 23054 -23316 23454 -23304
rect 22366 -23598 22968 -23348
rect 21288 -23646 22968 -23598
rect 20656 -23704 21056 -23696
rect 23054 -23690 23070 -23316
rect 23440 -23690 23454 -23316
rect 23544 -23568 24070 -23206
rect 25410 -23568 25512 -22730
rect 23544 -23646 25512 -23568
rect 23054 -23704 23454 -23690
<< via1 >>
rect 1638 -1200 2012 -826
rect 2190 -1200 2564 -826
rect 3606 -1200 3980 -826
rect 4350 -1198 4724 -824
rect 8088 -1200 8464 -822
rect 9982 -1206 10370 -818
rect 11200 -1204 11580 -822
rect 7372 -1444 7472 -1344
rect 12358 -1444 12458 -1344
rect 3046 -1694 3414 -1690
rect 3046 -1768 3050 -1694
rect 3050 -1768 3412 -1694
rect 3412 -1768 3414 -1694
rect 3046 -1772 3414 -1768
rect 4912 -1686 5280 -1682
rect 4912 -1760 4916 -1686
rect 4916 -1760 5278 -1686
rect 5278 -1760 5280 -1686
rect 4912 -1764 5280 -1760
rect 3168 -2656 3256 -2350
rect 3468 -2404 3556 -2370
rect 3468 -2654 3556 -2404
rect 3788 -2726 4544 -2044
rect 4780 -2404 4868 -2370
rect 4780 -2654 4868 -2404
rect 5080 -2656 5168 -2350
rect 12730 -1490 13494 -960
rect 23924 -1200 24302 -820
rect 7378 -1600 7478 -1500
rect 12184 -1600 12284 -1500
rect 7378 -1784 7478 -1684
rect 12006 -1784 12106 -1684
rect 3880 -3308 4452 -2870
rect 7434 -2198 7550 -2194
rect 7434 -2976 7444 -2198
rect 7444 -2976 7540 -2198
rect 7540 -2976 7550 -2198
rect 7434 -2982 7550 -2976
rect 7594 -2198 7710 -2194
rect 7594 -2976 7604 -2198
rect 7604 -2976 7700 -2198
rect 7700 -2976 7710 -2198
rect 7594 -2982 7710 -2976
rect 7752 -2198 7868 -2194
rect 7752 -2976 7762 -2198
rect 7762 -2976 7858 -2198
rect 7858 -2976 7868 -2198
rect 7752 -2982 7868 -2976
rect 7910 -2198 8026 -2194
rect 7910 -2976 7920 -2198
rect 7920 -2976 8016 -2198
rect 8016 -2976 8026 -2198
rect 7910 -2982 8026 -2976
rect 8068 -2198 8184 -2194
rect 8068 -2976 8078 -2198
rect 8078 -2976 8174 -2198
rect 8174 -2976 8184 -2198
rect 8068 -2982 8184 -2976
rect 8224 -2198 8340 -2192
rect 8224 -2976 8234 -2198
rect 8234 -2976 8330 -2198
rect 8330 -2976 8340 -2198
rect 8224 -2980 8340 -2976
rect 8382 -2198 8498 -2194
rect 8382 -2976 8392 -2198
rect 8392 -2976 8488 -2198
rect 8488 -2976 8498 -2198
rect 8382 -2982 8498 -2976
rect 8542 -2198 8658 -2192
rect 8542 -2976 8552 -2198
rect 8552 -2976 8648 -2198
rect 8648 -2976 8658 -2198
rect 8542 -2980 8658 -2976
rect 8698 -2198 8814 -2194
rect 8698 -2976 8708 -2198
rect 8708 -2976 8804 -2198
rect 8804 -2976 8814 -2198
rect 8698 -2982 8814 -2976
rect 8856 -2198 8972 -2194
rect 8856 -2976 8866 -2198
rect 8866 -2976 8962 -2198
rect 8962 -2976 8972 -2198
rect 8856 -2982 8972 -2976
rect 9014 -2198 9130 -2194
rect 9014 -2976 9024 -2198
rect 9024 -2976 9120 -2198
rect 9120 -2976 9130 -2198
rect 9014 -2982 9130 -2976
rect 9360 -2202 9476 -2198
rect 9360 -2980 9370 -2202
rect 9370 -2980 9466 -2202
rect 9466 -2980 9476 -2202
rect 9360 -2986 9476 -2980
rect 9518 -2202 9634 -2198
rect 9518 -2980 9528 -2202
rect 9528 -2980 9624 -2202
rect 9624 -2980 9634 -2202
rect 9518 -2986 9634 -2980
rect 9678 -2202 9794 -2198
rect 9678 -2980 9688 -2202
rect 9688 -2980 9784 -2202
rect 9784 -2980 9794 -2202
rect 9678 -2986 9794 -2980
rect 9836 -2202 9952 -2198
rect 9836 -2980 9846 -2202
rect 9846 -2980 9942 -2202
rect 9942 -2980 9952 -2202
rect 9836 -2986 9952 -2980
rect 9992 -2202 10108 -2198
rect 9992 -2980 10002 -2202
rect 10002 -2980 10098 -2202
rect 10098 -2980 10108 -2202
rect 9992 -2986 10108 -2980
rect 10152 -2202 10268 -2198
rect 10152 -2980 10162 -2202
rect 10162 -2980 10258 -2202
rect 10258 -2980 10268 -2202
rect 10152 -2986 10268 -2980
rect 10308 -2202 10424 -2198
rect 10308 -2980 10318 -2202
rect 10318 -2980 10414 -2202
rect 10414 -2980 10424 -2202
rect 10308 -2986 10424 -2980
rect 10466 -2202 10582 -2198
rect 10466 -2980 10476 -2202
rect 10476 -2980 10572 -2202
rect 10572 -2980 10582 -2202
rect 10466 -2986 10582 -2980
rect 10626 -2202 10742 -2198
rect 10626 -2980 10636 -2202
rect 10636 -2980 10732 -2202
rect 10732 -2980 10742 -2202
rect 10626 -2986 10742 -2980
rect 10782 -2202 10898 -2198
rect 10782 -2980 10792 -2202
rect 10792 -2980 10888 -2202
rect 10888 -2980 10898 -2202
rect 10782 -2986 10898 -2980
rect 10940 -2202 11056 -2198
rect 10940 -2980 10950 -2202
rect 10950 -2980 11046 -2202
rect 11046 -2980 11056 -2202
rect 10940 -2986 11056 -2980
rect 11310 -2180 11462 -2176
rect 11310 -2958 11462 -2180
rect 11310 -2964 11462 -2958
rect 13672 -1580 13852 -1576
rect 13672 -1752 13676 -1580
rect 13676 -1752 13848 -1580
rect 13848 -1752 13852 -1580
rect 13672 -1756 13852 -1752
rect 14082 -1538 14770 -1362
rect 11780 -3164 11972 -2980
rect 14202 -1960 14204 -1872
rect 14204 -1960 14242 -1872
rect 14242 -1960 14422 -1872
rect 14202 -1964 14422 -1960
rect 14738 -1924 14814 -1848
rect 14132 -2040 14238 -2024
rect 14132 -2074 14138 -2040
rect 14138 -2074 14230 -2040
rect 14230 -2074 14238 -2040
rect 14132 -2076 14238 -2074
rect 14132 -2156 14238 -2150
rect 14132 -2190 14136 -2156
rect 14136 -2190 14228 -2156
rect 14228 -2190 14238 -2156
rect 14132 -2202 14238 -2190
rect 15154 -1986 15226 -1982
rect 15154 -2066 15160 -1986
rect 15160 -2066 15200 -1986
rect 15200 -2066 15226 -1986
rect 15154 -2090 15226 -2066
rect 21962 -1966 22026 -1952
rect 21962 -2160 21974 -1966
rect 21974 -2160 22014 -1966
rect 22014 -2160 22026 -1966
rect 21962 -2174 22026 -2160
rect 14200 -2328 14204 -2258
rect 14204 -2328 14242 -2258
rect 14242 -2328 14420 -2258
rect 14200 -2350 14420 -2328
rect 14192 -2816 14260 -2748
rect 15154 -2522 15226 -2498
rect 15154 -2602 15160 -2522
rect 15160 -2602 15200 -2522
rect 15200 -2602 15226 -2522
rect 15154 -2606 15226 -2602
rect 21962 -2428 22026 -2414
rect 21962 -2622 21974 -2428
rect 21974 -2622 22014 -2428
rect 22014 -2622 22026 -2428
rect 21962 -2636 22026 -2622
rect 14738 -2740 14814 -2664
rect 22146 -2734 22288 -1854
rect 11426 -3386 11604 -3208
rect 1636 -5026 1920 -3600
rect 13942 -3128 14128 -3124
rect 13942 -3460 13950 -3128
rect 13950 -3460 14122 -3128
rect 14122 -3460 14128 -3128
rect 13942 -3470 14128 -3460
rect 15172 -3094 15938 -3048
rect 15172 -3126 15938 -3094
rect 14344 -3464 14520 -3152
rect 16124 -3514 16212 -3136
rect 16212 -3514 17524 -3136
rect 2668 -4088 2722 -4034
rect 2766 -4138 2950 -4134
rect 2766 -4714 2840 -4138
rect 2840 -4714 2874 -4138
rect 2874 -4714 2950 -4138
rect 2766 -4716 2950 -4714
rect 2668 -4818 2722 -4764
rect 3698 -4088 3752 -4034
rect 3472 -4138 3656 -4134
rect 3472 -4714 3546 -4138
rect 3546 -4714 3580 -4138
rect 3580 -4714 3656 -4138
rect 3472 -4716 3656 -4714
rect 3698 -4818 3752 -4764
rect 4584 -4088 4638 -4034
rect 4680 -4138 4864 -4134
rect 4680 -4714 4756 -4138
rect 4756 -4714 4790 -4138
rect 4790 -4714 4864 -4138
rect 4680 -4716 4864 -4714
rect 4584 -4818 4638 -4764
rect 5614 -4088 5668 -4034
rect 5386 -4138 5570 -4134
rect 5386 -4714 5462 -4138
rect 5462 -4714 5496 -4138
rect 5496 -4714 5570 -4138
rect 5386 -4716 5570 -4714
rect 5614 -4818 5668 -4764
rect 9146 -4152 9246 -4052
rect 11462 -4152 11562 -4052
rect 12112 -4316 15250 -4310
rect 2048 -5154 2454 -5122
rect 2048 -6772 2454 -5154
rect 3020 -5618 3400 -5438
rect 3622 -5441 3802 -5430
rect 3622 -5617 3656 -5441
rect 3656 -5617 3802 -5441
rect 3622 -5630 3802 -5617
rect 2620 -6045 2800 -6032
rect 2620 -6221 2764 -6045
rect 2764 -6221 2798 -6045
rect 2798 -6221 2800 -6045
rect 2620 -6232 2800 -6221
rect 3022 -6222 3402 -6042
rect 2048 -6798 2454 -6772
rect 3952 -6808 4374 -5116
rect 4534 -5441 4714 -5430
rect 4534 -5617 4680 -5441
rect 4680 -5617 4714 -5441
rect 4534 -5630 4714 -5617
rect 4936 -5618 5316 -5438
rect 4934 -6222 5314 -6042
rect 5536 -6045 5716 -6032
rect 5536 -6221 5538 -6045
rect 5538 -6221 5572 -6045
rect 5572 -6221 5716 -6045
rect 5536 -6232 5716 -6221
rect 9534 -4734 10888 -4324
rect 9534 -4970 10462 -4734
rect 10462 -4970 10476 -4734
rect 11780 -4810 11972 -4626
rect 12112 -4750 15250 -4316
rect 12112 -4760 15250 -4750
rect 9534 -5346 11224 -4970
rect 12122 -5346 12488 -4970
rect 12924 -5346 13168 -4970
rect 13276 -5346 13642 -4970
rect 14538 -5346 15284 -4970
rect 17508 -4750 17702 -4742
rect 17508 -5526 17514 -4750
rect 17514 -5004 17702 -4750
rect 17514 -5526 18002 -5004
rect 17508 -5530 18002 -5526
rect 3370 -7222 3478 -6962
rect 3620 -7214 3728 -6954
rect 2412 -7266 2520 -7254
rect 2412 -8042 2420 -7266
rect 2420 -8042 2512 -7266
rect 2512 -8042 2520 -7266
rect 2412 -8054 2520 -8042
rect 2570 -7266 2678 -7254
rect 2570 -8042 2578 -7266
rect 2578 -8042 2670 -7266
rect 2670 -8042 2678 -7266
rect 2570 -8054 2678 -8042
rect 2728 -7266 2836 -7254
rect 2728 -8042 2736 -7266
rect 2736 -8042 2828 -7266
rect 2828 -8042 2836 -7266
rect 2728 -8054 2836 -8042
rect 2886 -7266 2994 -7254
rect 2886 -8042 2894 -7266
rect 2894 -8042 2986 -7266
rect 2986 -8042 2994 -7266
rect 2886 -8054 2994 -8042
rect 3042 -7266 3150 -7254
rect 3042 -8042 3050 -7266
rect 3050 -8042 3142 -7266
rect 3142 -8042 3150 -7266
rect 3042 -8054 3150 -8042
rect 3202 -7266 3310 -7254
rect 3202 -8042 3210 -7266
rect 3210 -8042 3302 -7266
rect 3302 -8042 3310 -7266
rect 3202 -8054 3310 -8042
rect 3370 -8078 3478 -7906
rect 3620 -8078 3728 -7916
rect 3790 -7266 3894 -7254
rect 3790 -8044 3796 -7266
rect 3796 -8044 3888 -7266
rect 3888 -8044 3894 -7266
rect 3790 -8054 3894 -8044
rect 3946 -7266 4054 -7254
rect 3946 -8044 3954 -7266
rect 3954 -8044 4046 -7266
rect 4046 -8044 4054 -7266
rect 3946 -8054 4054 -8044
rect 4104 -7266 4212 -7254
rect 4104 -8044 4112 -7266
rect 4112 -8044 4204 -7266
rect 4204 -8044 4212 -7266
rect 4104 -8054 4212 -8044
rect 4262 -7266 4370 -7254
rect 4262 -8044 4270 -7266
rect 4270 -8044 4362 -7266
rect 4362 -8044 4370 -7266
rect 4262 -8054 4370 -8044
rect 4420 -7266 4528 -7254
rect 4420 -8044 4428 -7266
rect 4428 -8044 4520 -7266
rect 4520 -8044 4528 -7266
rect 4420 -8054 4528 -8044
rect 4578 -7266 4686 -7254
rect 4578 -8044 4586 -7266
rect 4586 -8044 4678 -7266
rect 4678 -8044 4686 -7266
rect 4578 -8054 4686 -8044
rect 7604 -5640 8962 -5608
rect 7604 -7366 8878 -5640
rect 8878 -7366 8962 -5640
rect 11666 -6000 11814 -5990
rect 11666 -6378 11814 -6000
rect 11666 -6388 11814 -6378
rect 11666 -6528 11814 -6518
rect 11666 -6906 11814 -6528
rect 11666 -6916 11814 -6906
rect 12924 -6392 13250 -5982
rect 12924 -6436 13250 -6392
rect 12924 -6468 13023 -6436
rect 13023 -6468 13250 -6436
rect 12810 -6528 12958 -6518
rect 12810 -6906 12958 -6528
rect 12810 -6916 12958 -6906
rect 13954 -6000 14102 -5990
rect 13954 -6378 14102 -6000
rect 13954 -6388 14102 -6378
rect 13954 -6528 14102 -6518
rect 13954 -6906 14102 -6528
rect 13954 -6916 14102 -6906
rect 16044 -7036 16148 -6554
rect 17014 -6890 17280 -6106
rect 19090 -5496 19230 -5466
rect 19090 -5672 19230 -5496
rect 19090 -5706 19230 -5672
rect 17528 -6108 17782 -6100
rect 17528 -6886 17532 -6108
rect 17532 -6886 17782 -6108
rect 17528 -6894 17782 -6886
rect 18146 -7036 18250 -6554
rect 21468 -5368 21556 -5334
rect 21468 -5544 21556 -5368
rect 21468 -5578 21556 -5544
rect 20580 -6104 20668 -6016
rect 19092 -6500 19232 -6474
rect 19092 -6694 19232 -6500
rect 19092 -6714 19232 -6694
rect 21468 -5754 21556 -5578
rect 21468 -5788 21556 -5754
rect 23006 -5246 23868 -4406
rect 22006 -6124 22302 -5996
rect 21470 -6364 21560 -6330
rect 21470 -6558 21560 -6364
rect 21470 -6592 21560 -6558
rect 21470 -6786 21560 -6592
rect 21470 -6820 21560 -6786
rect 22726 -6132 23002 -5852
rect 24796 -5830 25120 -4334
rect 24010 -6130 24210 -5930
rect 22262 -7202 24596 -6846
rect 7604 -7438 8962 -7366
rect 24230 -7454 24644 -7402
rect 24230 -7492 24237 -7454
rect 24237 -7492 24634 -7454
rect 24634 -7492 24644 -7454
rect 24230 -7540 24644 -7492
rect 9636 -9408 10048 -9406
rect 9636 -9922 10048 -9408
rect 24792 -10142 25112 -7416
rect 24792 -10144 25112 -10142
rect 15988 -11130 16648 -10464
rect 17142 -10898 18052 -10464
rect 2030 -11824 3298 -11314
rect 15036 -11798 15812 -11484
rect 17714 -11798 18284 -11310
rect 2030 -11974 3298 -11824
rect 2032 -12806 3288 -11974
rect 2032 -13766 2930 -12806
rect 15036 -12058 15812 -11798
rect 17714 -12066 18284 -11798
rect 7542 -12430 7572 -12270
rect 7572 -12430 7704 -12270
rect 9998 -12272 11440 -12268
rect 9998 -12432 11440 -12272
rect 11662 -12272 13104 -12268
rect 9998 -12434 11440 -12432
rect 11662 -12432 13104 -12272
rect 11662 -12434 13104 -12432
rect 20292 -12468 20464 -12298
rect 7346 -12910 7506 -12620
rect 16050 -14472 16548 -13980
rect 18384 -14042 19346 -13994
rect 18384 -14080 18949 -14042
rect 18949 -14080 19346 -14042
rect 18384 -14132 19346 -14080
rect 18384 -14456 18848 -14132
rect 19712 -14762 19844 -13440
rect 20214 -14482 20590 -13716
rect 20882 -14052 21736 -14030
rect 20882 -14306 20916 -14052
rect 20916 -14306 21698 -14052
rect 21698 -14306 21736 -14052
rect 18420 -15530 18784 -15164
rect 2148 -22284 2654 -22232
rect 2148 -22322 2545 -22284
rect 2545 -22322 2654 -22284
rect 2148 -22372 2654 -22322
rect 19884 -17992 20222 -16020
rect 20476 -16268 21250 -16010
rect 20474 -16332 21252 -16324
rect 20474 -16424 20476 -16332
rect 20476 -16424 21252 -16332
rect 20474 -16430 21252 -16424
rect 22612 -13924 23390 -13716
rect 23540 -13716 24316 -13714
rect 24316 -13716 24318 -13714
rect 23540 -13922 24318 -13716
rect 23628 -15592 24228 -14938
rect 20474 -16490 21252 -16482
rect 20474 -16582 20476 -16490
rect 20476 -16582 21252 -16490
rect 20474 -16588 21252 -16582
rect 20474 -16648 21252 -16640
rect 20474 -16740 20476 -16648
rect 20476 -16740 21252 -16648
rect 20474 -16746 21252 -16740
rect 20474 -16806 21252 -16798
rect 20474 -16898 20476 -16806
rect 20476 -16898 21252 -16806
rect 20474 -16904 21252 -16898
rect 20474 -16964 21252 -16956
rect 20474 -17056 20476 -16964
rect 20476 -17056 21252 -16964
rect 20474 -17062 21252 -17056
rect 20476 -17122 21254 -17114
rect 20476 -17214 21252 -17122
rect 21252 -17214 21254 -17122
rect 20476 -17220 21254 -17214
rect 21718 -17098 22090 -16590
rect 20474 -17280 21252 -17272
rect 20474 -17372 20476 -17280
rect 20476 -17372 21252 -17280
rect 20474 -17378 21252 -17372
rect 20474 -17438 21252 -17430
rect 20474 -17530 20476 -17438
rect 20476 -17530 21252 -17438
rect 20474 -17536 21252 -17530
rect 20474 -17596 21252 -17588
rect 20474 -17688 20476 -17596
rect 20476 -17688 21252 -17596
rect 20474 -17694 21252 -17688
rect 20476 -17756 21250 -17750
rect 20476 -18008 21250 -17756
rect 17768 -19030 19592 -18590
rect 22610 -16812 23388 -16604
rect 23540 -16606 24316 -16604
rect 24316 -16606 24318 -16604
rect 23540 -16812 24318 -16606
rect 23114 -20260 23386 -19984
rect 20718 -20882 20990 -20606
rect 20720 -22440 20992 -22168
rect 20664 -23696 21048 -23312
rect 23070 -23690 23440 -23316
<< metal2 >>
rect 1626 -826 2026 -812
rect 1626 -1200 1638 -826
rect 2012 -1200 2026 -826
rect 1626 -1212 2026 -1200
rect 2178 -826 2578 -812
rect 2178 -1200 2190 -826
rect 2564 -1200 2578 -826
rect 2178 -1212 2578 -1200
rect 3592 -826 3992 -812
rect 3592 -1200 3606 -826
rect 3980 -1200 3992 -826
rect 3592 -1212 3992 -1200
rect 4338 -824 4738 -812
rect 4338 -1198 4350 -824
rect 4724 -1198 4738 -824
rect 4338 -1212 4738 -1198
rect 8076 -822 8476 -812
rect 8076 -1200 8088 -822
rect 8464 -1200 8476 -822
rect 8076 -1210 8476 -1200
rect 9976 -818 10376 -812
rect 9976 -1206 9982 -818
rect 10370 -1206 10376 -818
rect 9976 -1210 10376 -1206
rect 11192 -822 11592 -812
rect 11192 -1204 11200 -822
rect 11580 -1204 11592 -822
rect 23912 -820 24312 -812
rect 14082 -936 23806 -852
rect 1626 -3600 1926 -1212
rect 2226 -1362 2526 -1212
rect 7542 -1220 9136 -1210
rect 1626 -7264 1636 -3600
rect 1920 -5026 1926 -3600
rect 1830 -6974 1926 -5026
rect 2026 -1662 2526 -1362
rect 6632 -1444 7372 -1344
rect 7472 -1444 7478 -1344
rect 2026 -5102 2326 -1662
rect 6632 -1672 6732 -1444
rect 3038 -1690 4632 -1680
rect 3038 -1772 3046 -1690
rect 3414 -1772 4632 -1690
rect 4904 -1682 6732 -1672
rect 4904 -1764 4912 -1682
rect 5280 -1764 6732 -1682
rect 4904 -1772 6732 -1764
rect 6812 -1600 7378 -1500
rect 7478 -1600 7484 -1500
rect 7542 -1562 7548 -1220
rect 9128 -1562 9136 -1220
rect 3038 -1780 4632 -1772
rect 4532 -1864 4632 -1780
rect 6812 -1864 6912 -1600
rect 4532 -1964 6912 -1864
rect 6974 -1784 7378 -1684
rect 7478 -1784 7484 -1684
rect 6974 -2026 7074 -1784
rect 7542 -1854 9136 -1562
rect 3772 -2044 4562 -2026
rect 3772 -2272 3788 -2044
rect 3162 -2350 3262 -2342
rect 3162 -2656 3168 -2350
rect 3256 -2656 3262 -2350
rect 3162 -3012 3262 -2656
rect 2622 -3264 3262 -3012
rect 3462 -2370 3562 -2356
rect 3462 -2654 3468 -2370
rect 3556 -2654 3562 -2370
rect 3462 -3044 3562 -2654
rect 3770 -2726 3788 -2272
rect 4544 -2726 4562 -2044
rect 6042 -2126 7074 -2026
rect 7428 -2084 9136 -1854
rect 5074 -2350 5174 -2342
rect 3770 -2742 4562 -2726
rect 4774 -2370 4874 -2356
rect 4774 -2654 4780 -2370
rect 4868 -2654 4874 -2370
rect 3864 -2870 4470 -2854
rect 3462 -3144 3798 -3044
rect 2622 -4034 2728 -3264
rect 2622 -4088 2668 -4034
rect 2722 -4088 2728 -4034
rect 2622 -4764 2728 -4088
rect 3692 -4034 3798 -3144
rect 3864 -3308 3880 -2870
rect 4452 -3308 4470 -2870
rect 4774 -3044 4874 -2654
rect 3864 -3324 4470 -3308
rect 4538 -3144 4874 -3044
rect 5074 -2656 5080 -2350
rect 5168 -2656 5174 -2350
rect 5074 -3012 5174 -2656
rect 5074 -3082 5714 -3012
rect 6042 -3082 6142 -2126
rect 7428 -2194 7556 -2084
rect 7428 -2982 7434 -2194
rect 7550 -2982 7556 -2194
rect 7428 -2992 7556 -2982
rect 7588 -2194 7716 -2184
rect 7588 -2982 7594 -2194
rect 7710 -2982 7716 -2194
rect 3692 -4088 3698 -4034
rect 3752 -4088 3798 -4034
rect 2756 -4134 2958 -4126
rect 2756 -4716 2766 -4134
rect 2950 -4716 2958 -4134
rect 2756 -4724 2958 -4716
rect 2622 -4818 2668 -4764
rect 2722 -4818 2728 -4764
rect 2622 -4824 2728 -4818
rect 2758 -4932 2958 -4724
rect 2026 -5122 2480 -5102
rect 2026 -6798 2048 -5122
rect 2454 -6798 2480 -5122
rect 2026 -6822 2480 -6798
rect 2610 -5132 2958 -4932
rect 3462 -4134 3664 -4126
rect 3462 -4716 3472 -4134
rect 3656 -4716 3664 -4134
rect 3462 -4724 3664 -4716
rect 3462 -4932 3662 -4724
rect 3692 -4764 3798 -4088
rect 3692 -4818 3698 -4764
rect 3752 -4818 3798 -4764
rect 3692 -4824 3798 -4818
rect 4538 -4034 4644 -3144
rect 5074 -3182 6142 -3082
rect 7588 -3092 7716 -2982
rect 7746 -2194 7874 -2084
rect 7746 -2982 7752 -2194
rect 7868 -2982 7874 -2194
rect 7746 -2992 7874 -2982
rect 7904 -2194 8032 -2184
rect 7904 -2982 7910 -2194
rect 8026 -2982 8032 -2194
rect 7904 -3092 8032 -2982
rect 8062 -2194 8190 -2084
rect 8062 -2982 8068 -2194
rect 8184 -2982 8190 -2194
rect 8062 -2992 8190 -2982
rect 8218 -2192 8346 -2184
rect 8218 -2980 8224 -2192
rect 8340 -2980 8346 -2192
rect 8218 -3092 8346 -2980
rect 8376 -2194 8504 -2084
rect 8376 -2982 8382 -2194
rect 8498 -2982 8504 -2194
rect 8376 -2992 8504 -2982
rect 8536 -2192 8664 -2184
rect 8536 -2980 8542 -2192
rect 8658 -2980 8664 -2192
rect 8536 -3092 8664 -2980
rect 8692 -2194 8820 -2084
rect 8692 -2982 8698 -2194
rect 8814 -2982 8820 -2194
rect 8692 -2992 8820 -2982
rect 8850 -2194 8978 -2184
rect 8850 -2982 8856 -2194
rect 8972 -2982 8978 -2194
rect 8850 -3092 8978 -2982
rect 9008 -2194 9136 -2084
rect 9008 -2982 9014 -2194
rect 9130 -2982 9136 -2194
rect 9008 -2992 9136 -2982
rect 9354 -1238 11062 -1210
rect 11192 -1212 11592 -1204
rect 12712 -960 13510 -946
rect 9354 -1640 9390 -1238
rect 11028 -1640 11062 -1238
rect 9354 -2088 11062 -1640
rect 9354 -2198 9482 -2088
rect 9354 -2986 9360 -2198
rect 9476 -2986 9482 -2198
rect 9354 -2996 9482 -2986
rect 9512 -2198 9640 -2188
rect 9512 -2986 9518 -2198
rect 9634 -2986 9640 -2198
rect 5074 -3264 5714 -3182
rect 4538 -4088 4584 -4034
rect 4638 -4088 4644 -4034
rect 4538 -4764 4644 -4088
rect 5608 -4034 5714 -3264
rect 5608 -4088 5614 -4034
rect 5668 -4088 5714 -4034
rect 4672 -4134 4874 -4126
rect 4672 -4716 4680 -4134
rect 4864 -4716 4874 -4134
rect 4672 -4724 4874 -4716
rect 4538 -4818 4584 -4764
rect 4638 -4818 4644 -4764
rect 4538 -4824 4644 -4818
rect 4674 -4932 4874 -4724
rect 3462 -5132 3812 -4932
rect 2610 -5430 2810 -5132
rect 3612 -5430 3812 -5132
rect 2610 -5438 3410 -5430
rect 2610 -5618 3020 -5438
rect 3400 -5618 3410 -5438
rect 2610 -5628 3410 -5618
rect 2610 -6032 2810 -5628
rect 2610 -6232 2620 -6032
rect 2800 -6232 2810 -6032
rect 3612 -5630 3622 -5430
rect 3802 -5630 3812 -5430
rect 3612 -6034 3812 -5630
rect 3012 -6042 3812 -6034
rect 3012 -6222 3022 -6042
rect 3402 -6222 3812 -6042
rect 3012 -6232 3812 -6222
rect 2610 -6740 2810 -6232
rect 2610 -6860 3484 -6740
rect 3612 -6860 3812 -6232
rect 3940 -5116 4386 -5102
rect 3940 -6808 3952 -5116
rect 4374 -6808 4386 -5116
rect 3364 -6962 3484 -6860
rect 1830 -7174 3158 -6974
rect 1830 -7254 2526 -7174
rect 2722 -7254 2842 -7174
rect 3036 -7254 3158 -7174
rect 3364 -7222 3370 -6962
rect 3478 -7222 3484 -6962
rect 1830 -7264 2412 -7254
rect 1626 -7274 2412 -7264
rect 2406 -8054 2412 -7274
rect 2520 -8054 2526 -7254
rect 2564 -8054 2570 -7254
rect 2678 -8054 2684 -7254
rect 2722 -8054 2728 -7254
rect 2836 -8054 2842 -7254
rect 2880 -8054 2886 -7254
rect 2994 -8054 3000 -7254
rect 3036 -8054 3042 -7254
rect 3150 -7554 3158 -7254
rect 3150 -8054 3156 -7554
rect 3196 -8054 3202 -7254
rect 3310 -8054 3316 -7254
rect 2564 -8134 2684 -8054
rect 2880 -8134 3000 -8054
rect 3196 -8134 3316 -8054
rect 3364 -7906 3484 -7222
rect 3364 -8078 3370 -7906
rect 3478 -8078 3484 -7906
rect 3614 -6954 3734 -6860
rect 3614 -7214 3620 -6954
rect 3728 -7214 3734 -6954
rect 3614 -7916 3734 -7214
rect 3940 -7014 4000 -6808
rect 4308 -6974 4386 -6808
rect 4524 -5132 4874 -4932
rect 5378 -4134 5580 -4126
rect 5378 -4716 5386 -4134
rect 5570 -4716 5580 -4134
rect 5378 -4724 5580 -4716
rect 5378 -4932 5578 -4724
rect 5608 -4764 5714 -4088
rect 5608 -4818 5614 -4764
rect 5668 -4818 5714 -4764
rect 5608 -4824 5714 -4818
rect 5378 -5132 5726 -4932
rect 4524 -5430 4724 -5132
rect 5526 -5430 5726 -5132
rect 4524 -5630 4534 -5430
rect 4714 -5630 4724 -5430
rect 4926 -5438 5726 -5430
rect 4926 -5618 4936 -5438
rect 5316 -5618 5726 -5438
rect 4926 -5628 5726 -5618
rect 4524 -6034 4724 -5630
rect 5526 -6032 5726 -5628
rect 4524 -6042 5324 -6034
rect 4524 -6222 4934 -6042
rect 5314 -6222 5324 -6042
rect 4524 -6232 5324 -6222
rect 5526 -6232 5536 -6032
rect 5716 -6232 5726 -6032
rect 4524 -6860 4724 -6232
rect 5526 -6860 5726 -6232
rect 7588 -5608 8978 -3092
rect 9512 -3096 9640 -2986
rect 9672 -2198 9800 -2088
rect 9672 -2986 9678 -2198
rect 9794 -2986 9800 -2198
rect 9672 -2996 9800 -2986
rect 9830 -2198 9958 -2188
rect 9830 -2986 9836 -2198
rect 9952 -2986 9958 -2198
rect 9830 -3096 9958 -2986
rect 9986 -2198 10114 -2088
rect 9986 -2986 9992 -2198
rect 10108 -2986 10114 -2198
rect 9986 -2996 10114 -2986
rect 10146 -2198 10274 -2188
rect 10146 -2986 10152 -2198
rect 10268 -2986 10274 -2198
rect 10146 -3096 10274 -2986
rect 10302 -2198 10430 -2088
rect 10302 -2986 10308 -2198
rect 10424 -2986 10430 -2198
rect 10302 -2996 10430 -2986
rect 10460 -2198 10588 -2188
rect 10460 -2986 10466 -2198
rect 10582 -2986 10588 -2198
rect 10460 -3096 10588 -2986
rect 10620 -2198 10748 -2088
rect 10620 -2986 10626 -2198
rect 10742 -2986 10748 -2198
rect 10620 -2996 10748 -2986
rect 10776 -2198 10904 -2188
rect 10776 -2986 10782 -2198
rect 10898 -2986 10904 -2198
rect 10776 -3096 10904 -2986
rect 10934 -2198 11062 -2088
rect 10934 -2986 10940 -2198
rect 11056 -2986 11062 -2198
rect 11300 -2176 11474 -1212
rect 12358 -1344 12458 -1338
rect 12184 -1500 12284 -1494
rect 12006 -1684 12106 -1678
rect 12006 -1874 12106 -1784
rect 12184 -1736 12284 -1600
rect 12358 -1586 12458 -1444
rect 12712 -1490 12730 -960
rect 13494 -1490 13510 -960
rect 14082 -1350 15334 -936
rect 12712 -1504 13510 -1490
rect 14070 -1362 15334 -1350
rect 14070 -1538 14082 -1362
rect 14770 -1508 15334 -1362
rect 15922 -1508 23806 -936
rect 23912 -1200 23924 -820
rect 24302 -1200 24312 -820
rect 23912 -1212 24312 -1200
rect 14770 -1532 23806 -1508
rect 14770 -1538 14782 -1532
rect 14070 -1542 14782 -1538
rect 13662 -1576 13862 -1566
rect 13662 -1586 13672 -1576
rect 12358 -1686 13672 -1586
rect 12184 -1836 13542 -1736
rect 13662 -1756 13672 -1686
rect 13852 -1756 13862 -1576
rect 13662 -1766 13862 -1756
rect 14356 -1702 15244 -1602
rect 12006 -1974 13372 -1874
rect 11300 -2964 11310 -2176
rect 11462 -2964 11474 -2176
rect 13272 -2204 13372 -1974
rect 13442 -1926 13542 -1836
rect 14356 -1858 14436 -1702
rect 14188 -1872 14436 -1858
rect 13662 -1926 13862 -1890
rect 13442 -2010 13862 -1926
rect 14188 -1964 14202 -1872
rect 14422 -1964 14436 -1872
rect 14188 -1978 14436 -1964
rect 14726 -1848 14826 -1836
rect 14726 -1924 14738 -1848
rect 14814 -1924 14826 -1848
rect 14726 -1936 14826 -1924
rect 14726 -2010 14806 -1936
rect 13442 -2024 14806 -2010
rect 13442 -2026 14132 -2024
rect 13662 -2076 14132 -2026
rect 14238 -2076 14806 -2024
rect 13662 -2090 14806 -2076
rect 15144 -1982 15244 -1702
rect 15144 -2090 15154 -1982
rect 15226 -2090 15244 -1982
rect 15402 -1838 23806 -1532
rect 15402 -2058 21844 -1838
rect 22136 -1854 23806 -1838
rect 21954 -1952 22034 -1942
rect 13662 -2150 14806 -2136
rect 13662 -2202 14132 -2150
rect 14238 -2202 14806 -2150
rect 13662 -2204 14806 -2202
rect 13272 -2216 14806 -2204
rect 15144 -2152 15244 -2090
rect 21954 -2152 21962 -1952
rect 15144 -2174 21962 -2152
rect 22026 -2174 22034 -1952
rect 15144 -2212 22034 -2174
rect 13272 -2304 13862 -2216
rect 13662 -2336 13862 -2304
rect 14186 -2258 14434 -2244
rect 14186 -2350 14200 -2258
rect 14420 -2350 14434 -2258
rect 14186 -2364 14434 -2350
rect 11300 -2974 11474 -2964
rect 14186 -2748 14266 -2742
rect 14186 -2816 14192 -2748
rect 14260 -2816 14266 -2748
rect 10934 -2996 11062 -2986
rect 11772 -2980 11980 -2972
rect 4308 -7014 4692 -6974
rect 3940 -7174 4692 -7014
rect 3940 -7254 4060 -7174
rect 4256 -7254 4376 -7174
rect 4572 -7254 4692 -7174
rect 3614 -8078 3620 -7916
rect 3728 -8078 3734 -7916
rect 3782 -8054 3790 -7254
rect 3894 -8054 3902 -7254
rect 3940 -8054 3946 -7254
rect 4054 -8054 4060 -7254
rect 4098 -8054 4104 -7254
rect 4212 -8054 4218 -7254
rect 4256 -8054 4262 -7254
rect 4370 -8054 4376 -7254
rect 4414 -8054 4420 -7254
rect 4528 -8054 4534 -7254
rect 4572 -8054 4578 -7254
rect 4686 -8054 4692 -7254
rect 5592 -7536 5692 -6860
rect 7588 -7438 7604 -5608
rect 8962 -7438 8978 -5608
rect 7588 -7454 8978 -7438
rect 9146 -4052 9246 -4046
rect 9146 -7536 9246 -4152
rect 9512 -4324 10904 -3096
rect 11772 -3164 11780 -2980
rect 11972 -3164 11980 -2980
rect 14186 -3038 14266 -2816
rect 14354 -2886 14434 -2364
rect 14726 -2652 14806 -2216
rect 15144 -2414 22034 -2376
rect 15144 -2436 21962 -2414
rect 15144 -2498 15244 -2436
rect 15144 -2606 15154 -2498
rect 15226 -2606 15244 -2498
rect 14726 -2664 14826 -2652
rect 14726 -2740 14738 -2664
rect 14814 -2740 14826 -2664
rect 14726 -2752 14826 -2740
rect 15144 -2886 15244 -2606
rect 14354 -2986 15244 -2886
rect 16192 -2550 21842 -2532
rect 16192 -3006 16208 -2550
rect 17532 -2752 21842 -2550
rect 21954 -2636 21962 -2436
rect 22026 -2636 22034 -2414
rect 21954 -2646 22034 -2636
rect 22136 -2734 22146 -1854
rect 22288 -2734 23806 -1854
rect 22136 -2752 23806 -2734
rect 17532 -3006 23812 -2752
rect 16192 -3022 23812 -3006
rect 14186 -3048 15950 -3038
rect 14186 -3098 15172 -3048
rect 11772 -3172 11980 -3164
rect 13934 -3124 14136 -3116
rect 11416 -3208 11616 -3198
rect 11416 -3386 11426 -3208
rect 11604 -3386 11616 -3208
rect 11416 -3398 11616 -3386
rect 11462 -4052 11568 -3398
rect 11562 -4152 11568 -4052
rect 11462 -4156 11568 -4152
rect 11462 -4158 11562 -4156
rect 9512 -5346 9534 -4324
rect 10888 -4734 10904 -4324
rect 11826 -4616 11926 -3172
rect 13934 -3470 13942 -3124
rect 14128 -3470 14136 -3124
rect 15160 -3126 15172 -3098
rect 15938 -3126 15950 -3048
rect 15160 -3134 15950 -3126
rect 16104 -3136 17546 -3120
rect 13934 -3476 14136 -3470
rect 14332 -3152 14532 -3140
rect 14332 -3464 14344 -3152
rect 14520 -3464 14532 -3152
rect 14332 -3476 14532 -3464
rect 13962 -3882 14102 -3476
rect 14360 -3640 14500 -3476
rect 16104 -3514 16124 -3136
rect 17524 -3514 17546 -3136
rect 16104 -3534 17546 -3514
rect 17668 -3530 23812 -3022
rect 14360 -3780 22856 -3640
rect 13962 -4022 22308 -3882
rect 12104 -4310 15264 -4298
rect 10476 -4958 10904 -4734
rect 11772 -4626 11980 -4616
rect 11772 -4810 11780 -4626
rect 11972 -4810 11980 -4626
rect 11772 -4816 11980 -4810
rect 12104 -4760 12112 -4310
rect 15250 -4760 15264 -4310
rect 12104 -4768 15264 -4760
rect 17500 -4742 17712 -4734
rect 12104 -4958 12504 -4768
rect 13260 -4958 13660 -4768
rect 10476 -4970 12504 -4958
rect 11224 -5346 12122 -4970
rect 12488 -5346 12504 -4970
rect 9512 -5358 12504 -5346
rect 12918 -4970 13178 -4958
rect 12918 -5346 12924 -4970
rect 13168 -5346 13178 -4970
rect 12918 -5358 13178 -5346
rect 13260 -4970 15296 -4958
rect 13260 -5346 13276 -4970
rect 13642 -5346 14538 -4970
rect 15284 -5346 15296 -4970
rect 17500 -4994 17508 -4742
rect 13260 -5358 15296 -5346
rect 17212 -5014 17508 -4994
rect 17702 -4994 17712 -4742
rect 17702 -5004 18012 -4994
rect 5592 -7636 9246 -7536
rect 2564 -8280 3316 -8134
rect 3782 -8134 3902 -8054
rect 4098 -8134 4218 -8054
rect 4414 -8134 4534 -8054
rect 2018 -10686 3318 -8280
rect 3782 -8282 4534 -8134
rect 2016 -11314 3318 -10686
rect 3780 -10450 5080 -8282
rect 9616 -9406 10068 -5358
rect 12998 -5896 13098 -5358
rect 17212 -5772 17232 -5014
rect 18002 -5530 18012 -5004
rect 21462 -5334 21562 -5328
rect 17990 -5772 18012 -5530
rect 17212 -5794 18012 -5772
rect 19082 -5466 19242 -5462
rect 19082 -5706 19090 -5466
rect 19230 -5706 19242 -5466
rect 12912 -5982 13260 -5896
rect 11660 -5990 11820 -5984
rect 11660 -6388 11666 -5990
rect 11814 -6388 11820 -5990
rect 11660 -6512 11820 -6388
rect 12912 -6468 12924 -5982
rect 13250 -6468 13260 -5982
rect 12912 -6482 13260 -6468
rect 13948 -5990 14108 -5984
rect 13948 -6388 13954 -5990
rect 14102 -6388 14108 -5990
rect 17500 -6092 17712 -5794
rect 19082 -6036 19242 -5706
rect 21462 -5788 21468 -5334
rect 21556 -5788 21562 -5334
rect 21462 -5794 21562 -5788
rect 21466 -6010 21562 -5794
rect 22168 -5990 22308 -4022
rect 22716 -5842 22856 -3780
rect 22972 -4394 23904 -4378
rect 22972 -4406 23036 -4394
rect 23488 -4406 23904 -4394
rect 22972 -5246 23006 -4406
rect 23868 -5246 23904 -4406
rect 22972 -5266 23036 -5246
rect 23488 -5266 23904 -5246
rect 22972 -5276 23904 -5266
rect 13948 -6402 14108 -6388
rect 16998 -6106 17298 -6092
rect 16998 -6402 17014 -6106
rect 13948 -6502 17014 -6402
rect 13948 -6512 14108 -6502
rect 11660 -6518 14108 -6512
rect 11660 -6916 11666 -6518
rect 11814 -6916 12810 -6518
rect 12958 -6916 13954 -6518
rect 14102 -6916 14108 -6518
rect 11660 -6922 14108 -6916
rect 16036 -6554 16156 -6544
rect 16036 -7036 16044 -6554
rect 16148 -7036 16156 -6554
rect 16998 -6890 17014 -6502
rect 17280 -6890 17298 -6106
rect 16998 -6902 17298 -6890
rect 17500 -6100 17790 -6092
rect 17500 -6894 17528 -6100
rect 17782 -6894 17790 -6100
rect 17500 -6902 17790 -6894
rect 17854 -6196 19242 -6036
rect 20574 -6016 21562 -6010
rect 20574 -6104 20580 -6016
rect 20668 -6104 21562 -6016
rect 20574 -6110 21562 -6104
rect 16036 -7424 16156 -7036
rect 16036 -7544 16904 -7424
rect 9616 -9922 9636 -9406
rect 10048 -9922 10068 -9406
rect 9616 -9948 10068 -9922
rect 3780 -10464 16668 -10450
rect 3780 -10468 15988 -10464
rect 3780 -11132 5904 -10468
rect 7226 -11124 12774 -10468
rect 13664 -11124 15988 -10468
rect 7226 -11130 15988 -11124
rect 16648 -11130 16668 -10464
rect 7226 -11132 16668 -11130
rect 3780 -11150 16668 -11132
rect 2016 -11974 2030 -11314
rect 3298 -11974 3318 -11314
rect 15028 -11482 15826 -11470
rect 15028 -11484 15304 -11482
rect 15554 -11484 15826 -11482
rect 2016 -13536 2032 -11974
rect 3288 -11990 3318 -11974
rect 5808 -11778 7106 -11760
rect 5808 -11790 7984 -11778
rect 3288 -12806 3304 -11990
rect 5808 -12116 5830 -11790
rect 7082 -11968 7984 -11790
rect 7082 -12116 7106 -11968
rect 5808 -12148 7106 -12116
rect 7534 -12270 7714 -12260
rect 7534 -12430 7542 -12270
rect 7704 -12272 7714 -12270
rect 7816 -12272 7984 -11968
rect 15028 -12058 15036 -11484
rect 15812 -12058 15826 -11484
rect 9978 -12268 13126 -12252
rect 9978 -12272 9998 -12268
rect 7704 -12428 9998 -12272
rect 7704 -12430 7714 -12428
rect 7534 -12440 7714 -12430
rect 9978 -12434 9998 -12428
rect 11440 -12434 11662 -12268
rect 13104 -12434 13126 -12268
rect 15028 -12262 15304 -12058
rect 15554 -12262 15826 -12058
rect 15028 -12272 15826 -12262
rect 9978 -12452 13126 -12434
rect 1900 -13570 2032 -13536
rect 2930 -13536 3304 -12806
rect 7334 -12620 7520 -12612
rect 7334 -12910 7346 -12620
rect 7506 -12910 7520 -12620
rect 2930 -13570 3682 -13536
rect 1900 -14770 1946 -13570
rect 3638 -14770 3682 -13570
rect 7334 -13976 7520 -12910
rect 7334 -13978 9618 -13976
rect 16042 -13978 16556 -13972
rect 7334 -13980 16556 -13978
rect 7334 -14146 16050 -13980
rect 7334 -14148 9618 -14146
rect 7334 -14154 7520 -14148
rect 16042 -14472 16050 -14146
rect 16548 -14472 16556 -13980
rect 16042 -14480 16556 -14472
rect 1900 -14810 3682 -14770
rect 16784 -20684 16904 -7544
rect 17854 -7546 18014 -6196
rect 19082 -6474 19242 -6196
rect 21466 -6324 21562 -6110
rect 22000 -5996 22308 -5990
rect 22000 -6124 22006 -5996
rect 22302 -6124 22308 -5996
rect 22000 -6130 22308 -6124
rect 22714 -5852 23014 -5842
rect 22714 -6132 22726 -5852
rect 23002 -6132 23014 -5852
rect 24010 -5930 24210 -1212
rect 24762 -4334 25158 -4298
rect 24762 -5830 24796 -4334
rect 25120 -5830 25158 -4334
rect 24004 -6130 24010 -5930
rect 24210 -6130 24216 -5930
rect 22714 -6142 23014 -6132
rect 17214 -7568 18014 -7546
rect 17214 -8326 17236 -7568
rect 17994 -8326 18014 -7568
rect 17214 -8346 18014 -8326
rect 18138 -6554 18258 -6546
rect 18138 -7036 18146 -6554
rect 18250 -7036 18258 -6554
rect 17112 -10446 18066 -10434
rect 17112 -10904 17124 -10446
rect 17812 -10464 18066 -10446
rect 18052 -10898 18066 -10464
rect 17812 -10904 18066 -10898
rect 17112 -10906 18066 -10904
rect 18138 -10970 18258 -7036
rect 19082 -6714 19092 -6474
rect 19232 -6714 19242 -6474
rect 19082 -7390 19242 -6714
rect 21464 -6330 21564 -6324
rect 21464 -6820 21470 -6330
rect 21560 -6820 21564 -6330
rect 21464 -6826 21564 -6820
rect 22244 -6836 24622 -6828
rect 22244 -6846 22880 -6836
rect 23376 -6846 24622 -6836
rect 22244 -7202 22262 -6846
rect 24596 -7202 24622 -6846
rect 22244 -7224 24622 -7202
rect 19082 -7402 24654 -7390
rect 19082 -7540 24230 -7402
rect 24644 -7540 24654 -7402
rect 19082 -7550 24654 -7540
rect 24762 -7416 25158 -5830
rect 24762 -10144 24792 -7416
rect 25112 -10144 25158 -7416
rect 24762 -10176 25158 -10144
rect 17400 -11090 18258 -10970
rect 17400 -20062 17520 -11090
rect 17700 -11310 18300 -11292
rect 17700 -12066 17714 -11310
rect 18284 -12066 18300 -11310
rect 17700 -15994 18300 -12066
rect 20278 -12298 20478 -12284
rect 20278 -12468 20292 -12298
rect 20464 -12468 20478 -12298
rect 20278 -12484 20478 -12468
rect 19698 -13440 19858 -13426
rect 19698 -13978 19712 -13440
rect 18372 -13994 19712 -13978
rect 18372 -14456 18384 -13994
rect 19346 -14132 19712 -13994
rect 18848 -14146 19712 -14132
rect 18848 -14456 18870 -14146
rect 18372 -14466 18870 -14456
rect 19698 -14762 19712 -14146
rect 19844 -14762 19858 -13440
rect 20328 -13702 20478 -12484
rect 20200 -13716 20600 -13702
rect 20200 -14482 20214 -13716
rect 20590 -14482 20600 -13716
rect 22596 -13714 24330 -13688
rect 22596 -13716 23540 -13714
rect 22596 -13924 22612 -13716
rect 23390 -13922 23540 -13716
rect 24318 -13922 24330 -13714
rect 23390 -13924 24330 -13922
rect 22596 -13956 24330 -13924
rect 20200 -14496 20600 -14482
rect 20856 -14030 21760 -14010
rect 20856 -14306 20882 -14030
rect 21736 -14306 21760 -14030
rect 20856 -14328 21760 -14306
rect 19698 -14776 19858 -14762
rect 20856 -15148 21256 -14328
rect 18402 -15164 21256 -15148
rect 18402 -15530 18420 -15164
rect 18784 -15530 21256 -15164
rect 18402 -15546 21256 -15530
rect 23584 -14938 24274 -13956
rect 18402 -15548 21222 -15546
rect 23584 -15592 23628 -14938
rect 24228 -15592 24274 -14938
rect 17700 -16010 21264 -15994
rect 17700 -16020 20476 -16010
rect 17700 -16410 19884 -16020
rect 17700 -16810 18944 -16410
rect 19854 -16810 19884 -16410
rect 17700 -17210 19884 -16810
rect 17700 -17610 18944 -17210
rect 19854 -17610 19884 -17210
rect 17700 -17992 19884 -17610
rect 20222 -16268 20476 -16020
rect 21250 -16268 21264 -16010
rect 20222 -16284 21264 -16268
rect 20222 -16470 20432 -16284
rect 20464 -16324 21704 -16312
rect 20464 -16430 20474 -16324
rect 21252 -16430 21704 -16324
rect 20464 -16442 21704 -16430
rect 20222 -16482 21264 -16470
rect 20222 -16588 20474 -16482
rect 21252 -16588 21264 -16482
rect 20222 -16600 21264 -16588
rect 21296 -16576 21704 -16442
rect 23584 -16576 24274 -15592
rect 21296 -16590 24330 -16576
rect 20222 -16786 20432 -16600
rect 21296 -16628 21718 -16590
rect 20464 -16640 21718 -16628
rect 20464 -16746 20474 -16640
rect 21252 -16746 21718 -16640
rect 20464 -16758 21718 -16746
rect 20222 -16798 21264 -16786
rect 20222 -16904 20474 -16798
rect 21252 -16904 21264 -16798
rect 20222 -16916 21264 -16904
rect 20222 -17102 20432 -16916
rect 21296 -16944 21718 -16758
rect 20464 -16956 21718 -16944
rect 20464 -17062 20474 -16956
rect 21252 -17062 21718 -16956
rect 20464 -17074 21718 -17062
rect 21296 -17098 21718 -17074
rect 22090 -16604 24330 -16590
rect 22090 -16812 22610 -16604
rect 23388 -16812 23540 -16604
rect 24318 -16812 24330 -16604
rect 22090 -16844 24330 -16812
rect 22090 -17098 22104 -16844
rect 20222 -17114 21264 -17102
rect 20222 -17220 20476 -17114
rect 21254 -17220 21264 -17114
rect 20222 -17232 21264 -17220
rect 21296 -17112 22104 -17098
rect 20222 -17418 20432 -17232
rect 21296 -17260 21704 -17112
rect 20464 -17272 21704 -17260
rect 20464 -17378 20474 -17272
rect 21252 -17378 21704 -17272
rect 20464 -17390 21704 -17378
rect 20222 -17430 21264 -17418
rect 20222 -17536 20474 -17430
rect 21252 -17536 21264 -17430
rect 20222 -17548 21264 -17536
rect 20222 -17734 20432 -17548
rect 21296 -17576 21704 -17390
rect 20464 -17588 21704 -17576
rect 20464 -17694 20474 -17588
rect 21252 -17694 21704 -17588
rect 20464 -17706 21704 -17694
rect 20222 -17750 21264 -17734
rect 20222 -17992 20476 -17750
rect 17700 -18008 20476 -17992
rect 21250 -18008 21264 -17750
rect 17700 -18010 21264 -18008
rect 17700 -18012 18300 -18010
rect 19854 -18022 21264 -18010
rect 17556 -18474 19806 -18462
rect 17556 -18744 17574 -18474
rect 19792 -18744 19806 -18474
rect 17556 -18758 17768 -18744
rect 17680 -19030 17768 -18758
rect 19592 -18758 19806 -18744
rect 19592 -19030 19684 -18758
rect 17680 -19098 19684 -19030
rect 23102 -19984 23402 -19970
rect 23102 -20062 23114 -19984
rect 17400 -20182 23114 -20062
rect 23102 -20260 23114 -20182
rect 23386 -20260 23402 -19984
rect 23102 -20270 23402 -20260
rect 20704 -20606 21004 -20592
rect 20704 -20684 20718 -20606
rect 16784 -20804 20718 -20684
rect 20704 -20882 20718 -20804
rect 20990 -20882 21004 -20606
rect 20704 -20892 21004 -20882
rect 6298 -21038 6540 -21026
rect 6298 -22222 6310 -21038
rect 2136 -22232 6310 -22222
rect 2136 -22372 2148 -22232
rect 2654 -22372 6310 -22232
rect 2136 -22382 6310 -22372
rect 6298 -23318 6310 -22382
rect 6530 -22222 6540 -21038
rect 11016 -21038 11258 -21024
rect 11016 -22222 11030 -21038
rect 6530 -22382 11030 -22222
rect 6530 -23318 6540 -22382
rect 6298 -23330 6540 -23318
rect 11016 -23318 11030 -22382
rect 11250 -22222 11258 -21038
rect 15738 -21036 15980 -21026
rect 15738 -22222 15744 -21036
rect 11250 -22382 15744 -22222
rect 11250 -23318 11258 -22382
rect 11016 -23328 11258 -23318
rect 15738 -23316 15744 -22382
rect 15970 -22222 15980 -21036
rect 20706 -22168 21006 -22154
rect 20706 -22222 20720 -22168
rect 15970 -22382 20720 -22222
rect 15970 -23316 15980 -22382
rect 20706 -22440 20720 -22382
rect 20992 -22440 21006 -22168
rect 20706 -22454 21006 -22440
rect 15738 -23330 15980 -23316
rect 20656 -23312 21056 -23304
rect 20656 -23696 20664 -23312
rect 21048 -23696 21056 -23312
rect 20656 -23704 21056 -23696
rect 23054 -23316 23454 -23304
rect 23054 -23690 23070 -23316
rect 23440 -23690 23454 -23316
rect 23054 -23704 23454 -23690
<< via2 >>
rect 1636 -5026 1830 -3912
rect 1636 -7264 1830 -5026
rect 7548 -1562 9128 -1220
rect 3788 -2726 4544 -2044
rect 3880 -3308 4452 -2870
rect 9390 -1640 11028 -1238
rect 4000 -5886 4308 -5136
rect 3956 -6210 4358 -5886
rect 4000 -6808 4308 -6210
rect 4000 -7014 4308 -6808
rect 12730 -1490 13494 -960
rect 15334 -1508 15922 -936
rect 16208 -3006 17532 -2550
rect 16124 -3514 17524 -3136
rect 17232 -5530 17508 -5014
rect 17508 -5530 17990 -5014
rect 17232 -5772 17990 -5530
rect 23036 -4406 23488 -4394
rect 23036 -5246 23488 -4406
rect 23036 -5266 23488 -5246
rect 5904 -11132 7226 -10468
rect 12774 -11124 13664 -10468
rect 15304 -11484 15554 -11482
rect 5830 -12116 7082 -11790
rect 15304 -11764 15554 -11484
rect 15038 -12026 15810 -11764
rect 15304 -12058 15554 -12026
rect 15304 -12262 15554 -12058
rect 1946 -13766 2032 -13570
rect 2032 -13766 2930 -13570
rect 2930 -13766 3638 -13570
rect 1946 -14770 3638 -13766
rect 16050 -14470 16546 -13980
rect 17236 -8326 17994 -7568
rect 17124 -10464 17812 -10446
rect 17124 -10898 17142 -10464
rect 17142 -10898 17812 -10464
rect 17124 -10904 17812 -10898
rect 22880 -6846 23376 -6836
rect 22880 -7182 23376 -6846
rect 17574 -18590 19792 -18474
rect 17574 -18744 17768 -18590
rect 17768 -18744 19592 -18590
rect 19592 -18744 19792 -18590
rect 6310 -23318 6530 -21038
rect 11030 -23318 11250 -21038
rect 15744 -23316 15970 -21036
<< metal3 >>
rect 15322 -936 15936 -922
rect 12712 -960 13510 -946
rect 7540 -1216 9136 -1210
rect 7540 -1562 7548 -1216
rect 9128 -1562 9136 -1216
rect 7540 -1570 9136 -1562
rect 9356 -1238 11066 -1212
rect 9356 -1640 9390 -1238
rect 11028 -1640 11066 -1238
rect 9356 -1654 11066 -1640
rect 12712 -1490 12730 -960
rect 13494 -1490 13510 -960
rect 12712 -1654 13510 -1490
rect 15322 -1508 15334 -936
rect 15922 -1508 15936 -936
rect 15322 -1520 15936 -1508
rect 3772 -2044 4562 -2026
rect 3772 -2272 3788 -2044
rect 3770 -2726 3788 -2272
rect 4544 -2726 4562 -2044
rect 3770 -2742 4562 -2726
rect 6984 -2454 9064 -1654
rect 9304 -2454 11384 -1654
rect 11624 -2454 13704 -1654
rect 13944 -2454 16024 -1654
rect 6984 -2854 16024 -2454
rect 3864 -2870 16024 -2854
rect 3864 -3308 3880 -2870
rect 4452 -2944 16024 -2870
rect 4452 -3308 9064 -2944
rect 3864 -3324 9064 -3308
rect 6984 -3730 9064 -3324
rect 9304 -3730 11384 -2944
rect 11624 -3730 13704 -2944
rect 13944 -3120 16024 -2944
rect 16192 -2550 17548 -2532
rect 16192 -3006 16208 -2550
rect 17532 -3006 17548 -2550
rect 16192 -3022 17548 -3006
rect 18342 -2652 20424 -1794
rect 20702 -2652 22784 -1798
rect 23468 -2652 25560 -1798
rect 18342 -3052 25560 -2652
rect 13944 -3136 17546 -3120
rect 13944 -3514 16124 -3136
rect 17524 -3514 17546 -3136
rect 13944 -3534 17546 -3514
rect 13944 -3730 16024 -3534
rect 1626 -3906 1842 -3900
rect 1626 -7268 1632 -3906
rect 1836 -7268 1842 -3906
rect 1932 -5120 4012 -3820
rect 4288 -5120 6372 -3818
rect 18342 -3874 20424 -3052
rect 19154 -4114 19556 -3874
rect 20702 -3878 22784 -3052
rect 23468 -3878 25560 -3052
rect 1932 -5136 6372 -5120
rect 1932 -5886 4000 -5136
rect 4308 -5886 6372 -5136
rect 1932 -5900 3956 -5886
rect 3886 -6194 3956 -5900
rect 1626 -7274 1842 -7268
rect 1934 -6210 3956 -6194
rect 4358 -5898 6372 -5886
rect 7792 -5266 9872 -4384
rect 10112 -5266 12192 -4384
rect 12432 -5266 14512 -4384
rect 14752 -5238 16832 -4384
rect 18342 -4906 20424 -4114
rect 21512 -4118 21914 -3878
rect 24304 -4118 24706 -3878
rect 20702 -4906 22784 -4118
rect 23468 -4378 25560 -4118
rect 23024 -4394 25560 -4378
rect 23024 -4906 23036 -4394
rect 17212 -5014 18012 -4994
rect 17212 -5238 17232 -5014
rect 14752 -5266 17232 -5238
rect 7792 -5538 17232 -5266
rect 7792 -5564 16832 -5538
rect 4358 -6192 4460 -5898
rect 4358 -6210 6374 -6192
rect 1934 -7014 4000 -6210
rect 4308 -7014 6374 -6210
rect 7792 -6466 9872 -5564
rect 10112 -6466 12192 -5564
rect 12432 -6466 14512 -5564
rect 14752 -6466 16832 -5564
rect 17212 -5772 17232 -5538
rect 17990 -5772 18012 -5014
rect 17212 -5794 18012 -5772
rect 18342 -5266 23036 -4906
rect 23488 -5266 25560 -4394
rect 18342 -5306 25560 -5266
rect 18342 -6194 20424 -5306
rect 19154 -6434 19556 -6194
rect 20702 -6198 22784 -5306
rect 23468 -6198 25560 -5306
rect 8690 -6996 8988 -6466
rect 11026 -6996 11324 -6466
rect 13324 -6996 13624 -6466
rect 15622 -6996 15922 -6466
rect 1934 -7028 6374 -7014
rect 1934 -8274 4014 -7028
rect 4290 -8272 6374 -7028
rect 7792 -7878 9872 -6996
rect 10112 -7878 12192 -6996
rect 12432 -7878 14512 -6996
rect 14752 -7878 16832 -6996
rect 18342 -7252 20424 -6434
rect 21512 -6438 21914 -6198
rect 24304 -6438 24706 -6198
rect 20702 -7252 22784 -6438
rect 22870 -6836 23384 -6830
rect 22870 -7182 22880 -6836
rect 23376 -7182 23384 -6836
rect 22870 -7190 23384 -7182
rect 23468 -7252 25560 -6438
rect 7792 -8176 16832 -7878
rect 7792 -9076 9872 -8176
rect 10112 -9076 12192 -8176
rect 12432 -9076 14512 -8176
rect 14752 -9076 16832 -8176
rect 17214 -7568 18014 -7546
rect 17214 -8326 17236 -7568
rect 17994 -8326 18014 -7568
rect 17214 -8346 18014 -8326
rect 18342 -7652 25560 -7252
rect 18342 -8514 20424 -7652
rect 19154 -8754 19556 -8514
rect 20702 -8518 22784 -7652
rect 23468 -8518 25560 -7652
rect 1706 -11760 5774 -9330
rect 8690 -9608 8988 -9076
rect 11026 -9608 11324 -9076
rect 18342 -9574 20424 -8754
rect 21512 -8758 21914 -8518
rect 24304 -8758 24706 -8518
rect 20702 -9574 22784 -8758
rect 23468 -9574 25560 -8758
rect 5864 -10412 7262 -10390
rect 5864 -11184 5884 -10412
rect 7244 -11184 7262 -10412
rect 5864 -11204 7262 -11184
rect 7792 -10476 9872 -9608
rect 10112 -10476 12192 -9608
rect 18342 -9974 25560 -9574
rect 7792 -10774 12192 -10476
rect 7792 -11688 9872 -10774
rect 10112 -11688 12192 -10774
rect 12752 -10430 13730 -10410
rect 12752 -11172 12774 -10430
rect 13704 -11172 13730 -10430
rect 12752 -11190 13730 -11172
rect 13824 -11470 15304 -10276
rect 15544 -11470 17024 -10276
rect 17112 -10446 17824 -10432
rect 17112 -10904 17124 -10446
rect 17812 -10904 17824 -10446
rect 18342 -10834 20424 -9974
rect 17112 -11156 17128 -10904
rect 17808 -11156 17824 -10904
rect 19154 -11074 19556 -10834
rect 20702 -10838 22784 -9974
rect 23468 -10838 25560 -9974
rect 17112 -11168 17824 -11156
rect 13824 -11482 17024 -11470
rect 1706 -11790 7106 -11760
rect 1706 -12116 5830 -11790
rect 7082 -12116 7106 -11790
rect 1706 -12148 7106 -12116
rect 1706 -13410 5774 -12148
rect 8690 -12168 8988 -11688
rect 7790 -13056 9870 -12168
rect 11026 -12172 11324 -11688
rect 13824 -11764 15304 -11482
rect 15554 -11764 17024 -11482
rect 13824 -11774 15038 -11764
rect 15026 -12018 15038 -11774
rect 13834 -12026 15038 -12018
rect 15810 -11774 17024 -11764
rect 15810 -12018 15830 -11774
rect 18342 -11958 20424 -11074
rect 21512 -11078 21914 -10838
rect 24304 -11078 24706 -10838
rect 20702 -11958 22784 -11078
rect 23468 -11958 25560 -11078
rect 15810 -12026 17034 -12018
rect 10116 -13056 12196 -12172
rect 7790 -13354 12196 -13056
rect 1898 -13570 3682 -13536
rect 1898 -13572 1946 -13570
rect 3638 -13572 3682 -13570
rect 1898 -14772 1932 -13572
rect 3642 -14772 3682 -13572
rect 7790 -14248 9870 -13354
rect 10116 -14252 12196 -13354
rect 13834 -12262 15304 -12026
rect 15554 -12262 17034 -12026
rect 13834 -12272 17034 -12262
rect 13834 -13504 15314 -12272
rect 15554 -13504 17034 -12272
rect 18342 -12358 25560 -11958
rect 18342 -13154 20424 -12358
rect 19154 -13394 19556 -13154
rect 20702 -13158 22784 -12358
rect 23468 -13158 25560 -12358
rect 16042 -13980 16556 -13972
rect 1898 -14810 3682 -14772
rect 16042 -14470 16050 -13980
rect 16546 -14470 16556 -13980
rect 16042 -14920 16556 -14470
rect 18342 -14194 20424 -13394
rect 21512 -13398 21914 -13158
rect 24304 -13398 24706 -13158
rect 20702 -14194 22784 -13398
rect 23468 -14194 25560 -13398
rect 18342 -14594 25560 -14194
rect 1808 -16466 5488 -14920
rect 5728 -16466 9408 -14920
rect 9648 -16466 13328 -14920
rect 13568 -16466 17248 -14920
rect 18342 -15474 20424 -14594
rect 19154 -15714 19556 -15474
rect 20702 -15478 22784 -14594
rect 23468 -15478 25560 -14594
rect 1808 -17098 17248 -16466
rect 1808 -18606 5488 -17098
rect 5728 -18606 9408 -17098
rect 9648 -18606 13328 -17098
rect 13568 -18606 17248 -17098
rect 18342 -16576 20424 -15714
rect 21512 -15718 21914 -15478
rect 24304 -15718 24706 -15478
rect 20702 -16576 22784 -15718
rect 23468 -16576 25560 -15718
rect 18342 -16976 25560 -16576
rect 18342 -17794 20424 -16976
rect 20702 -17798 22784 -16976
rect 23468 -17798 25560 -16976
rect 17544 -18462 19818 -18448
rect 17544 -18758 17556 -18462
rect 19806 -18758 19818 -18462
rect 17544 -18770 19818 -18758
rect 1818 -20952 6298 -18852
rect 1820 -21016 6298 -20952
rect 6538 -21016 11018 -18852
rect 11258 -21016 15738 -18852
rect 15978 -21016 20458 -18852
rect 20698 -21016 25178 -18852
rect 1820 -21036 25178 -21016
rect 1820 -21038 15744 -21036
rect 1820 -21250 6310 -21038
rect 1818 -23318 6310 -21250
rect 6530 -23318 11030 -21038
rect 11250 -23316 15744 -21038
rect 15970 -21412 25178 -21036
rect 15970 -23316 20458 -21412
rect 11250 -23318 20458 -23316
rect 1818 -23326 20458 -23318
rect 1818 -23330 11018 -23326
rect 11258 -23328 20458 -23326
rect 11258 -23330 15738 -23328
rect 15978 -23330 20458 -23328
rect 20698 -23330 25178 -21412
<< via3 >>
rect 7548 -1220 9128 -1216
rect 7548 -1562 9128 -1220
rect 15334 -1508 15922 -936
rect 3788 -2726 4544 -2044
rect 16208 -3006 17532 -2550
rect 1632 -3912 1836 -3906
rect 1632 -7264 1636 -3912
rect 1636 -7264 1830 -3912
rect 1830 -7264 1836 -3912
rect 1632 -7268 1836 -7264
rect 22880 -7182 23376 -6836
rect 17236 -8326 17994 -7568
rect 5884 -10468 7244 -10412
rect 5884 -11132 5904 -10468
rect 5904 -11132 7226 -10468
rect 7226 -11132 7244 -10468
rect 5884 -11184 7244 -11132
rect 12774 -10468 13704 -10430
rect 12774 -11124 13664 -10468
rect 13664 -11124 13704 -10468
rect 12774 -11172 13704 -11124
rect 17128 -10904 17808 -10448
rect 17128 -11156 17808 -10904
rect 1932 -14770 1946 -13572
rect 1946 -14770 3638 -13572
rect 3638 -14770 3642 -13572
rect 1932 -14772 3642 -14770
rect 17556 -18474 19806 -18462
rect 17556 -18744 17574 -18474
rect 17574 -18744 19792 -18474
rect 19792 -18744 19806 -18474
rect 17556 -18758 19806 -18744
<< mimcap >>
rect 7024 -1730 9024 -1690
rect 7024 -3650 7064 -1730
rect 8984 -3650 9024 -1730
rect 7024 -3690 9024 -3650
rect 9344 -1730 11344 -1690
rect 9344 -3650 9384 -1730
rect 11304 -3650 11344 -1730
rect 9344 -3690 11344 -3650
rect 11664 -1730 13664 -1690
rect 11664 -3650 11704 -1730
rect 13624 -3650 13664 -1730
rect 11664 -3690 13664 -3650
rect 13984 -1730 15984 -1690
rect 13984 -3650 14024 -1730
rect 15944 -3650 15984 -1730
rect 13984 -3690 15984 -3650
rect 18382 -1874 20382 -1834
rect 18382 -3794 18422 -1874
rect 20342 -3794 20382 -1874
rect 18382 -3834 20382 -3794
rect 20742 -1878 22742 -1838
rect 20742 -3798 20782 -1878
rect 22702 -3798 22742 -1878
rect 20742 -3838 22742 -3798
rect 23508 -1878 25508 -1838
rect 23508 -3798 23548 -1878
rect 25468 -3798 25508 -1878
rect 23508 -3838 25508 -3798
rect 1972 -3900 3972 -3860
rect 1972 -5820 2012 -3900
rect 3932 -5820 3972 -3900
rect 1972 -5860 3972 -5820
rect 4328 -3898 6328 -3858
rect 4328 -5818 4368 -3898
rect 6288 -5818 6328 -3898
rect 18382 -4194 20382 -4154
rect 4328 -5858 6328 -5818
rect 7832 -4464 9832 -4424
rect 1974 -6274 3974 -6234
rect 1974 -8194 2014 -6274
rect 3934 -8194 3974 -6274
rect 1974 -8234 3974 -8194
rect 4330 -6272 6330 -6232
rect 4330 -8192 4370 -6272
rect 6290 -8192 6330 -6272
rect 7832 -6384 7872 -4464
rect 9792 -6384 9832 -4464
rect 7832 -6424 9832 -6384
rect 10152 -4464 12152 -4424
rect 10152 -6384 10192 -4464
rect 12112 -6384 12152 -4464
rect 10152 -6424 12152 -6384
rect 12472 -4464 14472 -4424
rect 12472 -6384 12512 -4464
rect 14432 -6384 14472 -4464
rect 12472 -6424 14472 -6384
rect 14792 -4464 16792 -4424
rect 14792 -6384 14832 -4464
rect 16752 -6384 16792 -4464
rect 18382 -6114 18422 -4194
rect 20342 -6114 20382 -4194
rect 18382 -6154 20382 -6114
rect 20742 -4198 22742 -4158
rect 20742 -6118 20782 -4198
rect 22702 -6118 22742 -4198
rect 20742 -6158 22742 -6118
rect 23508 -4198 25508 -4158
rect 23508 -6118 23548 -4198
rect 25468 -6118 25508 -4198
rect 23508 -6158 25508 -6118
rect 14792 -6424 16792 -6384
rect 18382 -6514 20382 -6474
rect 4330 -8232 6330 -8192
rect 7832 -7076 9832 -7036
rect 7832 -8996 7872 -7076
rect 9792 -8996 9832 -7076
rect 7832 -9036 9832 -8996
rect 10152 -7076 12152 -7036
rect 10152 -8996 10192 -7076
rect 12112 -8996 12152 -7076
rect 10152 -9036 12152 -8996
rect 12472 -7076 14472 -7036
rect 12472 -8996 12512 -7076
rect 14432 -8996 14472 -7076
rect 12472 -9036 14472 -8996
rect 14792 -7076 16792 -7036
rect 14792 -8996 14832 -7076
rect 16752 -8996 16792 -7076
rect 18382 -8434 18422 -6514
rect 20342 -8434 20382 -6514
rect 18382 -8474 20382 -8434
rect 20742 -6518 22742 -6478
rect 20742 -8438 20782 -6518
rect 22702 -8438 22742 -6518
rect 20742 -8478 22742 -8438
rect 23508 -6518 25508 -6478
rect 23508 -8438 23548 -6518
rect 25468 -8438 25508 -6518
rect 23508 -8478 25508 -8438
rect 14792 -9036 16792 -8996
rect 18382 -8834 20382 -8794
rect 1734 -9410 5734 -9370
rect 1734 -13330 1774 -9410
rect 5694 -13330 5734 -9410
rect 7832 -9688 9832 -9648
rect 7832 -11608 7872 -9688
rect 9792 -11608 9832 -9688
rect 7832 -11648 9832 -11608
rect 10152 -9688 12152 -9648
rect 10152 -11608 10192 -9688
rect 12112 -11608 12152 -9688
rect 10152 -11648 12152 -11608
rect 13864 -10356 15264 -10316
rect 13864 -11676 13904 -10356
rect 15224 -11676 15264 -10356
rect 13864 -11716 15264 -11676
rect 15584 -10356 16984 -10316
rect 15584 -11676 15624 -10356
rect 16944 -11676 16984 -10356
rect 18382 -10754 18422 -8834
rect 20342 -10754 20382 -8834
rect 18382 -10794 20382 -10754
rect 20742 -8838 22742 -8798
rect 20742 -10758 20782 -8838
rect 22702 -10758 22742 -8838
rect 20742 -10798 22742 -10758
rect 23508 -8838 25508 -8798
rect 23508 -10758 23548 -8838
rect 25468 -10758 25508 -8838
rect 23508 -10798 25508 -10758
rect 15584 -11716 16984 -11676
rect 18382 -11154 20382 -11114
rect 13874 -12098 15274 -12058
rect 1734 -13370 5734 -13330
rect 7836 -12252 9836 -12212
rect 7836 -14172 7876 -12252
rect 9796 -14172 9836 -12252
rect 7836 -14212 9836 -14172
rect 10156 -12252 12156 -12212
rect 10156 -14172 10196 -12252
rect 12116 -14172 12156 -12252
rect 13874 -13418 13914 -12098
rect 15234 -13418 15274 -12098
rect 13874 -13458 15274 -13418
rect 15594 -12098 16994 -12058
rect 15594 -13418 15634 -12098
rect 16954 -13418 16994 -12098
rect 18382 -13074 18422 -11154
rect 20342 -13074 20382 -11154
rect 18382 -13114 20382 -13074
rect 20742 -11158 22742 -11118
rect 20742 -13078 20782 -11158
rect 22702 -13078 22742 -11158
rect 20742 -13118 22742 -13078
rect 23508 -11158 25508 -11118
rect 23508 -13078 23548 -11158
rect 25468 -13078 25508 -11158
rect 23508 -13118 25508 -13078
rect 15594 -13458 16994 -13418
rect 10156 -14212 12156 -14172
rect 18382 -13474 20382 -13434
rect 1848 -15006 5448 -14966
rect 1848 -18526 1888 -15006
rect 5408 -18526 5448 -15006
rect 1848 -18566 5448 -18526
rect 5768 -15006 9368 -14966
rect 5768 -18526 5808 -15006
rect 9328 -18526 9368 -15006
rect 5768 -18566 9368 -18526
rect 9688 -15006 13288 -14966
rect 9688 -18526 9728 -15006
rect 13248 -18526 13288 -15006
rect 9688 -18566 13288 -18526
rect 13608 -15006 17208 -14966
rect 13608 -18526 13648 -15006
rect 17168 -18526 17208 -15006
rect 18382 -15394 18422 -13474
rect 20342 -15394 20382 -13474
rect 18382 -15434 20382 -15394
rect 20742 -13478 22742 -13438
rect 20742 -15398 20782 -13478
rect 22702 -15398 22742 -13478
rect 20742 -15438 22742 -15398
rect 23508 -13478 25508 -13438
rect 23508 -15398 23548 -13478
rect 25468 -15398 25508 -13478
rect 23508 -15438 25508 -15398
rect 18382 -15794 20382 -15754
rect 18382 -17714 18422 -15794
rect 20342 -17714 20382 -15794
rect 18382 -17754 20382 -17714
rect 20742 -15798 22742 -15758
rect 20742 -17718 20782 -15798
rect 22702 -17718 22742 -15798
rect 20742 -17758 22742 -17718
rect 23508 -15798 25508 -15758
rect 23508 -17718 23548 -15798
rect 25468 -17718 25508 -15798
rect 23508 -17758 25508 -17718
rect 13608 -18566 17208 -18526
rect 1858 -18932 6258 -18892
rect 1858 -23252 1898 -18932
rect 6218 -23252 6258 -18932
rect 1858 -23292 6258 -23252
rect 6578 -18932 10978 -18892
rect 6578 -23252 6618 -18932
rect 10938 -23252 10978 -18932
rect 6578 -23292 10978 -23252
rect 11298 -18932 15698 -18892
rect 11298 -23252 11338 -18932
rect 15658 -23252 15698 -18932
rect 11298 -23292 15698 -23252
rect 16018 -18932 20418 -18892
rect 16018 -23252 16058 -18932
rect 20378 -23252 20418 -18932
rect 16018 -23292 20418 -23252
rect 20738 -18932 25138 -18892
rect 20738 -23252 20778 -18932
rect 25098 -23252 25138 -18932
rect 20738 -23292 25138 -23252
<< mimcapcontact >>
rect 7064 -3650 8984 -1730
rect 9384 -3650 11304 -1730
rect 11704 -3650 13624 -1730
rect 14024 -3650 15944 -1730
rect 18422 -3794 20342 -1874
rect 20782 -3798 22702 -1878
rect 23548 -3798 25468 -1878
rect 2012 -5820 3932 -3900
rect 4368 -5818 6288 -3898
rect 2014 -8194 3934 -6274
rect 4370 -8192 6290 -6272
rect 7872 -6384 9792 -4464
rect 10192 -6384 12112 -4464
rect 12512 -6384 14432 -4464
rect 14832 -6384 16752 -4464
rect 18422 -6114 20342 -4194
rect 20782 -6118 22702 -4198
rect 23548 -6118 25468 -4198
rect 7872 -8996 9792 -7076
rect 10192 -8996 12112 -7076
rect 12512 -8996 14432 -7076
rect 14832 -8996 16752 -7076
rect 18422 -8434 20342 -6514
rect 20782 -8438 22702 -6518
rect 23548 -8438 25468 -6518
rect 1774 -13330 5694 -9410
rect 7872 -11608 9792 -9688
rect 10192 -11608 12112 -9688
rect 13904 -11676 15224 -10356
rect 15624 -11676 16944 -10356
rect 18422 -10754 20342 -8834
rect 20782 -10758 22702 -8838
rect 23548 -10758 25468 -8838
rect 7876 -14172 9796 -12252
rect 10196 -14172 12116 -12252
rect 13914 -13418 15234 -12098
rect 15634 -13418 16954 -12098
rect 18422 -13074 20342 -11154
rect 20782 -13078 22702 -11158
rect 23548 -13078 25468 -11158
rect 1888 -18526 5408 -15006
rect 5808 -18526 9328 -15006
rect 9728 -18526 13248 -15006
rect 13648 -18526 17168 -15006
rect 18422 -15394 20342 -13474
rect 20782 -15398 22702 -13478
rect 23548 -15398 25468 -13478
rect 18422 -17714 20342 -15794
rect 20782 -17718 22702 -15798
rect 23548 -17718 25468 -15798
rect 1898 -23252 6218 -18932
rect 6618 -23252 10938 -18932
rect 11338 -23252 15658 -18932
rect 16058 -23252 20378 -18932
rect 20778 -23252 25098 -18932
<< metal4 >>
rect 15322 -936 15936 -922
rect 7540 -1216 9136 -1210
rect 7540 -1562 7548 -1216
rect 9128 -1562 9136 -1216
rect 7540 -1729 9136 -1562
rect 15322 -1508 15334 -936
rect 15922 -1508 15936 -936
rect 15322 -1729 15936 -1508
rect 7063 -1730 9136 -1729
rect 3772 -2044 4562 -2026
rect 3772 -2726 3788 -2044
rect 4544 -2272 4562 -2044
rect 7063 -2272 7064 -1730
rect 4544 -2726 7064 -2272
rect 3772 -2742 7064 -2726
rect 7063 -3650 7064 -2742
rect 8984 -1758 9136 -1730
rect 9383 -1730 11305 -1729
rect 8984 -2454 8985 -1758
rect 9383 -2454 9384 -1730
rect 8984 -2944 9384 -2454
rect 8984 -3650 8985 -2944
rect 7063 -3651 8985 -3650
rect 9383 -3650 9384 -2944
rect 11304 -2454 11305 -1730
rect 11703 -1730 13625 -1729
rect 11703 -2454 11704 -1730
rect 11304 -2944 11704 -2454
rect 11304 -3650 11305 -2944
rect 9383 -3651 11305 -3650
rect 11703 -3650 11704 -2944
rect 13624 -2454 13625 -1730
rect 14023 -1730 15945 -1729
rect 14023 -2454 14024 -1730
rect 13624 -2944 14024 -2454
rect 13624 -3650 13625 -2944
rect 11703 -3651 13625 -3650
rect 14023 -3650 14024 -2944
rect 15944 -2532 15945 -1730
rect 19330 -1873 19434 -1778
rect 18421 -1874 20343 -1873
rect 15944 -2550 17548 -2532
rect 15944 -3006 16208 -2550
rect 17532 -3006 17548 -2550
rect 15944 -3022 17548 -3006
rect 15944 -3650 15945 -3022
rect 14023 -3651 15945 -3650
rect 18421 -3794 18422 -1874
rect 20342 -2652 20343 -1874
rect 21690 -1877 21794 -1782
rect 24456 -1877 24560 -1782
rect 20781 -1878 22703 -1877
rect 20781 -2652 20782 -1878
rect 20342 -3052 20782 -2652
rect 20342 -3794 20343 -3052
rect 18421 -3795 20343 -3794
rect 2920 -3899 3024 -3800
rect 5276 -3897 5380 -3798
rect 4367 -3898 6289 -3897
rect 2011 -3900 3933 -3899
rect 1626 -3906 2012 -3900
rect 1626 -7268 1632 -3906
rect 1836 -5820 2012 -3906
rect 3932 -4072 3933 -3900
rect 4367 -4072 4368 -3898
rect 3932 -4398 4368 -4072
rect 3932 -5820 3933 -4398
rect 4367 -5818 4368 -4398
rect 6288 -5818 6289 -3898
rect 19154 -4193 19556 -3795
rect 20781 -3798 20782 -3052
rect 22702 -2652 22703 -1878
rect 23547 -1878 25469 -1877
rect 23547 -2652 23548 -1878
rect 22702 -3052 23548 -2652
rect 22702 -3798 22703 -3052
rect 20781 -3799 22703 -3798
rect 23547 -3798 23548 -3052
rect 25468 -3798 25469 -1878
rect 23547 -3799 25469 -3798
rect 18421 -4194 20343 -4193
rect 7871 -4464 9793 -4463
rect 7871 -5372 7872 -4464
rect 7780 -5476 7872 -5372
rect 4367 -5819 6289 -5818
rect 1836 -5821 3933 -5820
rect 1836 -6273 2088 -5821
rect 2794 -6273 3160 -5821
rect 5138 -6271 5504 -5819
rect 4369 -6272 6291 -6271
rect 1836 -6274 3935 -6273
rect 1836 -7268 2014 -6274
rect 1626 -7274 2014 -7268
rect 2013 -8194 2014 -7274
rect 3934 -7480 3935 -6274
rect 4369 -7480 4370 -6272
rect 3934 -7806 4370 -7480
rect 3934 -8194 3935 -7806
rect 4369 -8192 4370 -7806
rect 6290 -8192 6291 -6272
rect 7871 -6384 7872 -5476
rect 9792 -5266 9793 -4464
rect 10191 -4464 12113 -4463
rect 10191 -5266 10192 -4464
rect 9792 -5564 10192 -5266
rect 9792 -6384 9793 -5564
rect 7871 -6385 9793 -6384
rect 10191 -6384 10192 -5564
rect 12112 -5266 12113 -4464
rect 12511 -4464 14433 -4463
rect 12511 -5266 12512 -4464
rect 12112 -5564 12512 -5266
rect 12112 -6384 12113 -5564
rect 10191 -6385 12113 -6384
rect 12511 -6384 12512 -5564
rect 14432 -5266 14433 -4464
rect 14831 -4464 16753 -4463
rect 14831 -5266 14832 -4464
rect 14432 -5564 14832 -5266
rect 14432 -6384 14433 -5564
rect 12511 -6385 14433 -6384
rect 14831 -6384 14832 -5564
rect 16752 -5372 16753 -4464
rect 16752 -5476 16846 -5372
rect 16752 -6384 16753 -5476
rect 18421 -6114 18422 -4194
rect 20342 -4906 20343 -4194
rect 21512 -4197 21914 -3799
rect 24304 -4197 24706 -3799
rect 20781 -4198 22703 -4197
rect 20781 -4906 20782 -4198
rect 20342 -5306 20782 -4906
rect 20342 -6114 20343 -5306
rect 18421 -6115 20343 -6114
rect 14831 -6385 16753 -6384
rect 8690 -7075 8988 -6385
rect 11026 -7075 11324 -6385
rect 13324 -7075 13624 -6385
rect 15622 -7075 15922 -6385
rect 19154 -6513 19556 -6115
rect 20781 -6118 20782 -5306
rect 22702 -4906 22703 -4198
rect 23547 -4198 25469 -4197
rect 23547 -4906 23548 -4198
rect 22702 -5306 23548 -4906
rect 22702 -6118 22703 -5306
rect 20781 -6119 22703 -6118
rect 23547 -6118 23548 -5306
rect 25468 -6118 25469 -4198
rect 23547 -6119 25469 -6118
rect 18421 -6514 20343 -6513
rect 7871 -7076 9793 -7075
rect 7871 -7984 7872 -7076
rect 7780 -8088 7872 -7984
rect 4369 -8193 6291 -8192
rect 2013 -8195 3935 -8194
rect 2922 -8288 3026 -8195
rect 5278 -8286 5382 -8193
rect 7871 -8996 7872 -8088
rect 9792 -7878 9793 -7076
rect 10191 -7076 12113 -7075
rect 10191 -7878 10192 -7076
rect 9792 -8176 10192 -7878
rect 9792 -8996 9793 -8176
rect 7871 -8997 9793 -8996
rect 10191 -8996 10192 -8176
rect 12112 -7878 12113 -7076
rect 12511 -7076 14433 -7075
rect 12511 -7878 12512 -7076
rect 12112 -8176 12512 -7878
rect 12112 -8996 12113 -8176
rect 10191 -8997 12113 -8996
rect 12511 -8996 12512 -8176
rect 14432 -7878 14433 -7076
rect 14831 -7076 16753 -7075
rect 14831 -7878 14832 -7076
rect 14432 -8176 14832 -7878
rect 14432 -8996 14433 -8176
rect 12511 -8997 14433 -8996
rect 14831 -8996 14832 -8176
rect 16752 -7802 16753 -7076
rect 17214 -7568 18014 -7546
rect 17214 -7802 17236 -7568
rect 16752 -8102 17236 -7802
rect 16752 -8996 16753 -8102
rect 17214 -8326 17236 -8102
rect 17994 -8326 18014 -7568
rect 17214 -8346 18014 -8326
rect 18421 -8434 18422 -6514
rect 20342 -7252 20343 -6514
rect 21512 -6517 21914 -6119
rect 24304 -6517 24706 -6119
rect 20781 -6518 22703 -6517
rect 20781 -7252 20782 -6518
rect 20342 -7652 20782 -7252
rect 20342 -8434 20343 -7652
rect 18421 -8435 20343 -8434
rect 19154 -8833 19556 -8435
rect 20781 -8438 20782 -7652
rect 22702 -6828 22703 -6518
rect 23547 -6518 25469 -6517
rect 23547 -6828 23548 -6518
rect 22702 -6836 23548 -6828
rect 22702 -7182 22880 -6836
rect 23376 -7182 23548 -6836
rect 22702 -7652 23548 -7182
rect 22702 -8438 22703 -7652
rect 20781 -8439 22703 -8438
rect 23547 -8438 23548 -7652
rect 25468 -8438 25469 -6518
rect 23547 -8439 25469 -8438
rect 14831 -8997 16753 -8996
rect 18421 -8834 20343 -8833
rect 1773 -9410 5695 -9409
rect 1773 -13330 1774 -9410
rect 5694 -10390 5695 -9410
rect 8690 -9687 8988 -8997
rect 11026 -9687 11324 -8997
rect 7871 -9688 9793 -9687
rect 5694 -10412 7262 -10390
rect 5694 -11184 5884 -10412
rect 7244 -11184 7262 -10412
rect 7871 -10596 7872 -9688
rect 7780 -10700 7872 -10596
rect 5694 -11204 7262 -11184
rect 5694 -13330 5695 -11204
rect 7871 -11608 7872 -10700
rect 9792 -10476 9793 -9688
rect 10191 -9688 12113 -9687
rect 10191 -10476 10192 -9688
rect 9792 -10774 10192 -10476
rect 9792 -11608 9793 -10774
rect 7871 -11609 9793 -11608
rect 10191 -11608 10192 -10774
rect 12112 -10596 12113 -9688
rect 13903 -10356 15225 -10355
rect 13903 -10410 13904 -10356
rect 12752 -10430 13904 -10410
rect 12112 -10700 12198 -10596
rect 12112 -11608 12113 -10700
rect 12752 -11172 12774 -10430
rect 13704 -11172 13904 -10430
rect 12752 -11190 13904 -11172
rect 10191 -11609 12113 -11608
rect 8690 -12251 8988 -11609
rect 11026 -12251 11324 -11609
rect 13903 -11676 13904 -11190
rect 15224 -10396 15225 -10356
rect 15623 -10356 16945 -10355
rect 15623 -10396 15624 -10356
rect 15224 -10608 15624 -10396
rect 15224 -10964 15225 -10608
rect 15623 -10964 15624 -10608
rect 15224 -11068 15624 -10964
rect 15224 -11676 15225 -11068
rect 13903 -11677 15225 -11676
rect 15623 -11676 15624 -11068
rect 16944 -10434 16945 -10356
rect 16944 -10448 17824 -10434
rect 16944 -11156 17128 -10448
rect 17808 -11156 17824 -10448
rect 18421 -10754 18422 -8834
rect 20342 -9574 20343 -8834
rect 21512 -8837 21914 -8439
rect 24304 -8837 24706 -8439
rect 20781 -8838 22703 -8837
rect 20781 -9574 20782 -8838
rect 20342 -9974 20782 -9574
rect 20342 -10754 20343 -9974
rect 18421 -10755 20343 -10754
rect 19154 -11153 19556 -10755
rect 20781 -10758 20782 -9974
rect 22702 -9574 22703 -8838
rect 23547 -8838 25469 -8837
rect 23547 -9574 23548 -8838
rect 22702 -9974 23548 -9574
rect 22702 -10758 22703 -9974
rect 20781 -10759 22703 -10758
rect 23547 -10758 23548 -9974
rect 25468 -10758 25469 -8838
rect 23547 -10759 25469 -10758
rect 16944 -11168 17824 -11156
rect 18421 -11154 20343 -11153
rect 16944 -11676 16945 -11168
rect 15623 -11677 16945 -11676
rect 14052 -12097 14260 -11677
rect 16656 -12097 16864 -11677
rect 13913 -12098 15235 -12097
rect 7875 -12252 9797 -12251
rect 7875 -13160 7876 -12252
rect 7790 -13264 7876 -13160
rect 1773 -13331 5695 -13330
rect 1900 -13572 3680 -13538
rect 1900 -14772 1932 -13572
rect 3642 -14772 3680 -13572
rect 7875 -14172 7876 -13264
rect 9796 -13056 9797 -12252
rect 10195 -12252 12117 -12251
rect 10195 -13056 10196 -12252
rect 9796 -13354 10196 -13056
rect 9796 -14172 9797 -13354
rect 7875 -14173 9797 -14172
rect 10195 -14172 10196 -13354
rect 12116 -13160 12117 -12252
rect 13913 -12706 13914 -12098
rect 13820 -12810 13914 -12706
rect 12116 -13264 12210 -13160
rect 12116 -14172 12117 -13264
rect 13913 -13418 13914 -12810
rect 15234 -12706 15235 -12098
rect 15633 -12098 16955 -12097
rect 15633 -12706 15634 -12098
rect 15234 -12810 15634 -12706
rect 15234 -13142 15235 -12810
rect 15633 -13142 15634 -12810
rect 15234 -13354 15634 -13142
rect 15234 -13418 15235 -13354
rect 13913 -13419 15235 -13418
rect 15633 -13418 15634 -13354
rect 16954 -12706 16955 -12098
rect 16954 -12810 17048 -12706
rect 16954 -13418 16955 -12810
rect 18421 -13074 18422 -11154
rect 20342 -11958 20343 -11154
rect 21512 -11157 21914 -10759
rect 24304 -11157 24706 -10759
rect 20781 -11158 22703 -11157
rect 20781 -11958 20782 -11158
rect 20342 -12358 20782 -11958
rect 20342 -13074 20343 -12358
rect 18421 -13075 20343 -13074
rect 15633 -13419 16955 -13418
rect 19154 -13473 19556 -13075
rect 20781 -13078 20782 -12358
rect 22702 -11958 22703 -11158
rect 23547 -11158 25469 -11157
rect 23547 -11958 23548 -11158
rect 22702 -12358 23548 -11958
rect 22702 -13078 22703 -12358
rect 20781 -13079 22703 -13078
rect 23547 -13078 23548 -12358
rect 25468 -13078 25469 -11158
rect 23547 -13079 25469 -13078
rect 10195 -14173 12117 -14172
rect 18421 -13474 20343 -13473
rect 1900 -15005 3680 -14772
rect 1887 -15006 5409 -15005
rect 1887 -16714 1888 -15006
rect 1804 -16818 1888 -16714
rect 1887 -18526 1888 -16818
rect 5408 -16466 5409 -15006
rect 5807 -15006 9329 -15005
rect 5807 -16466 5808 -15006
rect 5408 -17098 5808 -16466
rect 5408 -18526 5409 -17098
rect 1887 -18527 5409 -18526
rect 5807 -18526 5808 -17098
rect 9328 -16466 9329 -15006
rect 9727 -15006 13249 -15005
rect 9727 -16466 9728 -15006
rect 9328 -17098 9728 -16466
rect 9328 -18526 9329 -17098
rect 5807 -18527 9329 -18526
rect 9727 -18526 9728 -17098
rect 13248 -16466 13249 -15006
rect 13647 -15006 17169 -15005
rect 13647 -16466 13648 -15006
rect 13248 -17098 13648 -16466
rect 13248 -18526 13249 -17098
rect 9727 -18527 13249 -18526
rect 13647 -18526 13648 -17098
rect 17168 -16714 17169 -15006
rect 18421 -15394 18422 -13474
rect 20342 -14194 20343 -13474
rect 21512 -13477 21914 -13079
rect 24304 -13477 24706 -13079
rect 20781 -13478 22703 -13477
rect 20781 -14194 20782 -13478
rect 20342 -14594 20782 -14194
rect 20342 -15394 20343 -14594
rect 18421 -15395 20343 -15394
rect 19154 -15793 19556 -15395
rect 20781 -15398 20782 -14594
rect 22702 -14194 22703 -13478
rect 23547 -13478 25469 -13477
rect 23547 -14194 23548 -13478
rect 22702 -14594 23548 -14194
rect 22702 -15398 22703 -14594
rect 20781 -15399 22703 -15398
rect 23547 -15398 23548 -14594
rect 25468 -15398 25469 -13478
rect 23547 -15399 25469 -15398
rect 18421 -15794 20343 -15793
rect 17168 -16818 17250 -16714
rect 17168 -18526 17169 -16818
rect 18421 -17714 18422 -15794
rect 20342 -16576 20343 -15794
rect 21512 -15797 21914 -15399
rect 24304 -15797 24706 -15399
rect 20781 -15798 22703 -15797
rect 20781 -16576 20782 -15798
rect 20342 -16976 20782 -16576
rect 20342 -17714 20343 -16976
rect 18421 -17715 20343 -17714
rect 19330 -17802 19434 -17715
rect 20781 -17718 20782 -16976
rect 22702 -16576 22703 -15798
rect 23547 -15798 25469 -15797
rect 23547 -16576 23548 -15798
rect 22702 -16976 23548 -16576
rect 22702 -17718 22703 -16976
rect 20781 -17719 22703 -17718
rect 23547 -17718 23548 -16976
rect 25468 -17718 25469 -15798
rect 23547 -17719 25469 -17718
rect 21690 -17806 21794 -17719
rect 24456 -17806 24560 -17719
rect 13647 -18527 17169 -18526
rect 17542 -18462 19822 -18442
rect 17542 -18758 17556 -18462
rect 19806 -18758 19822 -18462
rect 17542 -18931 19822 -18758
rect 1897 -18932 6219 -18931
rect 1897 -21040 1898 -18932
rect 1820 -21144 1898 -21040
rect 1897 -23252 1898 -21144
rect 6218 -20766 6219 -18932
rect 6617 -18932 10939 -18931
rect 6617 -20766 6618 -18932
rect 6218 -21440 6618 -20766
rect 6218 -23252 6219 -21440
rect 1897 -23253 6219 -23252
rect 6617 -23252 6618 -21440
rect 10938 -20766 10939 -18932
rect 11337 -18932 15659 -18931
rect 11337 -20766 11338 -18932
rect 10938 -21440 11338 -20766
rect 10938 -23252 10939 -21440
rect 6617 -23253 10939 -23252
rect 11337 -23252 11338 -21440
rect 15658 -20766 15659 -18932
rect 16057 -18932 20379 -18931
rect 16057 -20766 16058 -18932
rect 15658 -21440 16058 -20766
rect 15658 -23252 15659 -21440
rect 11337 -23253 15659 -23252
rect 16057 -23252 16058 -21440
rect 20378 -20766 20379 -18932
rect 20777 -18932 25099 -18931
rect 20777 -20766 20778 -18932
rect 20378 -21440 20778 -20766
rect 20378 -23252 20379 -21440
rect 16057 -23253 20379 -23252
rect 20777 -23252 20778 -21440
rect 25098 -21040 25099 -18932
rect 25098 -21144 25182 -21040
rect 25098 -23252 25099 -21144
rect 20777 -23253 25099 -23252
<< labels >>
flabel metal2 2178 -1212 2578 -812 0 FreeSans 1200 0 0 0 avdd
port 1 nsew
flabel metal2 1626 -1212 2026 -812 0 FreeSans 1200 0 0 0 avss
port 2 nsew
flabel metal2 8076 -1212 8476 -812 0 FreeSans 1200 0 0 0 dvdd
port 3 nsew
flabel metal2 9976 -1212 10376 -812 0 FreeSans 1200 0 0 0 dvss
port 4 nsew
flabel metal2 11192 -1212 11592 -812 0 FreeSans 1200 0 0 0 ibias
port 5 nsew
flabel metal2 3592 -1212 3992 -812 0 FreeSans 1200 0 0 0 ena
port 6 nsew
flabel metal2 4338 -1212 4738 -812 0 FreeSans 1200 0 0 0 standby
port 7 nsew
flabel metal2 23912 -1212 24312 -812 0 FreeSans 1200 0 0 0 dout
port 8 nsew
flabel metal1 23054 -23704 23454 -23304 0 FreeSans 1200 0 0 0 xout
port 9 nsew
flabel metal1 20656 -23704 21056 -23304 0 FreeSans 1200 0 0 0 xin
port 10 nsew
flabel metal1 19460 -14978 19640 -13228 0 FreeSans 400 0 0 0 vrb
flabel metal1 22240 -14982 22400 -14170 0 FreeSans 400 0 0 0 vg1
flabel metal1 22120 -11668 25450 -10450 0 FreeSans 3200 0 0 0 avdd_ip
flabel metal1 18284 -11798 21916 -11292 0 FreeSans 3200 0 0 0 avss_ip
flabel metal2 18932 -14146 19712 -13978 0 FreeSans 400 0 0 0 vg2
flabel metal1 21956 -15750 22156 -14384 0 FreeSans 400 0 0 0 vbreg
flabel metal2 7082 -11968 7984 -11778 0 FreeSans 800 0 0 0 icnode
flabel metal2 5592 -7636 9246 -7536 0 FreeSans 800 0 0 0 standby_33
flabel metal2 6632 -1444 7372 -1344 0 FreeSans 800 0 0 0 standby_ip
flabel metal2 6812 -1600 7378 -1500 0 FreeSans 800 0 0 0 ena_ip
flabel metal2 6974 -1784 7378 -1684 0 FreeSans 800 0 0 0 standby_b
flabel viali 8878 -7250 10492 -5640 0 FreeSans 3200 0 0 0 dvdd_ip
flabel viali 8900 -5476 10462 -4316 0 FreeSans 3200 0 0 0 dvss_ip
flabel metal2 13962 -4022 22308 -3882 0 FreeSans 800 0 0 0 dout_ip
flabel metal2 14360 -3780 22856 -3640 0 FreeSans 800 0 0 0 dout_filt
flabel metal2 11826 -4626 11926 -3164 0 FreeSans 800 0 0 0 ibias_ip
flabel metal2 12998 -5906 13098 -5346 0 FreeSans 800 0 0 0 vbp
flabel metal2 13948 -6502 17014 -6402 0 FreeSans 800 0 0 0 tail
flabel metal1 16648 -6108 16728 -5530 0 FreeSans 800 0 0 0 vn
flabel metal2 17500 -6100 17712 -5772 0 FreeSans 800 0 0 0 xin_buf
flabel metal2 19082 -6474 19242 -5706 0 FreeSans 800 0 0 0 inv_in
flabel metal2 20668 -6110 21562 -6010 0 FreeSans 800 0 0 0 inv_m1
flabel metal1 21718 -6828 21818 -5328 0 FreeSans 800 0 0 0 inv_m2
flabel metal1 3772 -2624 4122 -1842 0 FreeSans 1600 0 0 0 x3.dvdd
flabel metal1 2300 -2608 2652 -1842 0 FreeSans 1600 0 0 0 x3.dvss
flabel metal1 3872 -6560 4122 -5102 0 FreeSans 1600 0 0 0 x3.avdd
flabel metal1 2300 -5042 2456 -3770 0 FreeSans 1200 0 0 0 x3.avss
flabel metal1 2894 -2090 3278 -1842 0 FreeSans 1200 0 0 0 x3.in
flabel metal2 2622 -3264 3262 -3012 0 FreeSans 800 0 0 0 x3.in_b
flabel metal2 3612 -6860 3812 -5630 0 FreeSans 1200 0 0 0 x3.out_b
flabel metal2 2610 -6860 2810 -6232 0 FreeSans 1200 0 0 0 x3.out
flabel metal1 4214 -2624 4564 -1842 0 FreeSans 1600 0 0 0 x4.dvdd
flabel metal1 5684 -2608 6036 -1842 0 FreeSans 1600 0 0 0 x4.dvss
flabel metal1 4214 -6560 4464 -5102 0 FreeSans 1600 0 0 0 x4.avdd
flabel metal1 5880 -5042 6036 -3770 0 FreeSans 1200 0 0 0 x4.avss
flabel metal1 5058 -2090 5442 -1842 0 FreeSans 1200 0 0 0 x4.in
flabel metal2 5074 -3264 5714 -3012 0 FreeSans 800 0 0 0 x4.in_b
flabel metal2 4524 -6860 4724 -5630 0 FreeSans 1200 0 0 0 x4.out_b
flabel metal2 5526 -6860 5726 -6232 0 FreeSans 1200 0 0 0 x4.out
flabel space 14070 -1550 14782 -1350 0 FreeSans 800 0 0 0 x7.dvdd
flabel metal1 13936 -3476 14136 -3116 0 FreeSans 800 0 0 0 x7.clkin
flabel metal1 14332 -3476 14532 -3266 0 FreeSans 800 0 0 0 x7.clkout
flabel metal2 13662 -2090 13862 -1890 0 FreeSans 800 0 0 0 x7.ena
flabel metal2 13662 -1766 13862 -1566 0 FreeSans 800 0 0 0 x7.stby
flabel metal2 13662 -2336 13862 -2136 0 FreeSans 800 0 0 0 x7.stby_b
flabel metal2 14186 -3098 15172 -3038 0 FreeSans 400 0 0 0 x7.clk_disable
flabel metal1 13940 -1280 14916 -1180 0 FreeSans 800 0 0 0 x7.dvss
flabel metal2 14356 -1702 15244 -1602 0 FreeSans 400 0 0 0 x7.ena_done_b
flabel metal2 14354 -2986 15244 -2886 0 FreeSans 400 0 0 0 x7.stby_done_b
flabel locali 14345 -2825 14379 -2791 0 FreeSans 200 0 0 0 x7.x5.A
flabel locali 14277 -2825 14311 -2791 0 FreeSans 200 0 0 0 x7.x5.A
flabel locali 14209 -2549 14243 -2515 0 FreeSans 200 0 0 0 x7.x5.TE_B
flabel locali 14277 -2549 14311 -2515 0 FreeSans 200 0 0 0 x7.x5.TE_B
flabel locali 14209 -2825 14243 -2791 0 FreeSans 200 0 0 0 x7.x5.A
flabel locali 14141 -2825 14175 -2791 0 FreeSans 200 0 0 0 x7.x5.A
flabel locali 14413 -2825 14447 -2791 0 FreeSans 200 0 0 0 x7.x5.Z
flabel locali 14073 -2825 14107 -2791 0 FreeSans 200 0 0 0 x7.x5.Z
flabel metal1 14515 -2549 14549 -2515 0 FreeSans 200 0 0 0 x7.x5.VPWR
flabel metal1 13971 -2549 14005 -2515 0 FreeSans 200 0 0 0 x7.x5.VGND
flabel nwell 14515 -2549 14549 -2515 0 FreeSans 200 0 0 0 x7.x5.VPB
flabel pwell 13971 -2549 14005 -2515 0 FreeSans 200 0 0 0 x7.x5.VNB
rlabel comment 13988 -2486 13988 -2486 6 x7.x5.einvn_0
rlabel metal1 13940 -2854 14036 -2486 3 x7.x5.VGND
rlabel metal1 14484 -2854 14580 -2486 3 x7.x5.VPWR
flabel locali 14073 -2462 14107 -2428 0 FreeSans 200 0 0 0 x7.x3.X
flabel locali 14141 -2090 14175 -2056 0 FreeSans 200 0 0 0 x7.x3.B1
flabel locali 14141 -2186 14175 -2152 0 FreeSans 200 0 0 0 x7.x3.A1
flabel locali 14209 -2090 14243 -2056 0 FreeSans 200 0 0 0 x7.x3.B1
flabel locali 14209 -1906 14243 -1872 0 FreeSans 200 0 0 0 x7.x3.B2
flabel locali 14413 -2462 14447 -2428 0 FreeSans 200 0 0 0 x7.x3.X
flabel locali 14209 -2278 14243 -2244 0 FreeSans 200 0 0 0 x7.x3.A2
flabel locali 14209 -2186 14243 -2152 0 FreeSans 200 0 0 0 x7.x3.A1
flabel locali 13971 -1906 14005 -1872 0 FreeSans 200 0 0 0 x7.x3.VGND
flabel locali 14515 -1906 14549 -1872 0 FreeSans 200 0 0 0 x7.x3.VPWR
flabel locali 14209 -1814 14243 -1780 0 FreeSans 200 0 0 0 x7.x3.C1
flabel metal1 14515 -1814 14549 -1780 0 FreeSans 200 0 0 0 x7.x3.VPWR
flabel metal1 13971 -1814 14005 -1780 0 FreeSans 200 0 0 0 x7.x3.VGND
flabel nwell 14515 -1814 14549 -1780 0 FreeSans 200 0 0 0 x7.x3.VPB
flabel pwell 13971 -1814 14005 -1780 0 FreeSans 200 0 0 0 x7.x3.VNB
rlabel comment 13988 -1750 13988 -1750 6 x7.x3.a221o_1
rlabel metal1 13940 -2486 14036 -1750 3 x7.x3.VGND
rlabel metal1 14484 -2486 14580 -1750 3 x7.x3.VPWR
flabel metal1 14512 -1733 14541 -1680 0 FreeSans 200 0 0 0 x7.sky130_fd_sc_hd__tapvpwrvgnd_1_3.VPWR
flabel metal1 13970 -1730 14008 -1679 0 FreeSans 200 0 0 0 x7.sky130_fd_sc_hd__tapvpwrvgnd_1_3.VGND
rlabel comment 13988 -1658 13988 -1658 6 x7.sky130_fd_sc_hd__tapvpwrvgnd_1_3.tapvpwrvgnd_1
rlabel metal1 13940 -1750 14036 -1658 3 x7.sky130_fd_sc_hd__tapvpwrvgnd_1_3.VGND
rlabel metal1 14484 -1750 14580 -1658 3 x7.sky130_fd_sc_hd__tapvpwrvgnd_1_3.VPWR
flabel metal1 15220 -2324 16926 -2260 0 FreeSans 800 0 0 0 x7.x2.dvdd
flabel metal1 15202 -2872 16908 -2808 0 FreeSans 800 0 0 0 x7.x2.dvss
flabel metal1 14726 -2576 14826 -2476 0 FreeSans 800 0 0 0 x7.x2.clkin
flabel metal1 14726 -2752 14826 -2652 0 FreeSans 800 0 0 0 x7.x2.ena
flabel space 15350 -2634 15544 -2584 0 FreeSans 400 0 0 0 x7.x2.gated_clk
flabel metal1 15854 -2548 17556 -2516 0 FreeSans 400 0 0 0 x7.x2.Qb1
flabel metal1 18062 -2548 19766 -2516 0 FreeSans 400 0 0 0 x7.x2.Qb2
flabel space 21663 -2741 21729 -2522 0 FreeSans 400 0 0 0 x7.x2.done
flabel metal2 15144 -2616 15244 -2376 0 FreeSans 800 0 0 0 x7.x2.doneb
flabel locali 17266 -2620 17295 -2585 0 FreeSans 200 0 0 0 x7.x2.x2.Q
flabel locali 17568 -2617 17590 -2584 0 FreeSans 200 0 0 0 x7.x2.x2.Q_N
flabel locali 16993 -2685 17027 -2651 0 FreeSans 400 0 0 0 x7.x2.x2.RESET_B
flabel locali 15817 -2549 15851 -2515 0 FreeSans 400 0 0 0 x7.x2.x2.D
flabel locali 15542 -2549 15576 -2515 0 FreeSans 400 0 0 0 x7.x2.x2.CLK
flabel locali 15542 -2617 15576 -2583 0 FreeSans 400 0 0 0 x7.x2.x2.CLK
flabel locali 16993 -2617 17027 -2583 0 FreeSans 400 0 0 0 x7.x2.x2.RESET_B
flabel metal1 15541 -2855 15575 -2821 0 FreeSans 200 0 0 0 x7.x2.x2.VGND
flabel metal1 15541 -2311 15575 -2277 0 FreeSans 200 0 0 0 x7.x2.x2.VPWR
flabel nwell 15541 -2311 15575 -2277 0 FreeSans 200 0 0 0 x7.x2.x2.VPB
flabel pwell 15541 -2855 15575 -2821 0 FreeSans 200 0 0 0 x7.x2.x2.VNB
rlabel comment 15512 -2838 15512 -2838 4 x7.x2.x2.dfrbp_1
rlabel locali 16993 -2711 17041 -2631 1 x7.x2.x2.RESET_B
rlabel locali 16933 -2631 17041 -2557 1 x7.x2.x2.RESET_B
rlabel metal1 16981 -2691 17039 -2682 1 x7.x2.x2.RESET_B
rlabel metal1 16921 -2645 16979 -2582 1 x7.x2.x2.RESET_B
rlabel metal1 16921 -2654 17039 -2645 1 x7.x2.x2.RESET_B
rlabel metal1 16261 -2654 16391 -2645 1 x7.x2.x2.RESET_B
rlabel metal1 16261 -2682 17039 -2654 1 x7.x2.x2.RESET_B
rlabel metal1 16261 -2691 16391 -2682 1 x7.x2.x2.RESET_B
rlabel metal1 15512 -2886 17628 -2790 1 x7.x2.x2.VGND
rlabel metal1 15512 -2342 17628 -2246 1 x7.x2.x2.VPWR
flabel locali 19474 -2620 19503 -2585 0 FreeSans 200 0 0 0 x7.x2.x3.Q
flabel locali 19776 -2617 19798 -2584 0 FreeSans 200 0 0 0 x7.x2.x3.Q_N
flabel locali 19201 -2685 19235 -2651 0 FreeSans 400 0 0 0 x7.x2.x3.RESET_B
flabel locali 18025 -2549 18059 -2515 0 FreeSans 400 0 0 0 x7.x2.x3.D
flabel locali 17750 -2549 17784 -2515 0 FreeSans 400 0 0 0 x7.x2.x3.CLK
flabel locali 17750 -2617 17784 -2583 0 FreeSans 400 0 0 0 x7.x2.x3.CLK
flabel locali 19201 -2617 19235 -2583 0 FreeSans 400 0 0 0 x7.x2.x3.RESET_B
flabel metal1 17749 -2855 17783 -2821 0 FreeSans 200 0 0 0 x7.x2.x3.VGND
flabel metal1 17749 -2311 17783 -2277 0 FreeSans 200 0 0 0 x7.x2.x3.VPWR
flabel nwell 17749 -2311 17783 -2277 0 FreeSans 200 0 0 0 x7.x2.x3.VPB
flabel pwell 17749 -2855 17783 -2821 0 FreeSans 200 0 0 0 x7.x2.x3.VNB
rlabel comment 17720 -2838 17720 -2838 4 x7.x2.x3.dfrbp_1
rlabel locali 19201 -2711 19249 -2631 1 x7.x2.x3.RESET_B
rlabel locali 19141 -2631 19249 -2557 1 x7.x2.x3.RESET_B
rlabel metal1 19189 -2691 19247 -2682 1 x7.x2.x3.RESET_B
rlabel metal1 19129 -2645 19187 -2582 1 x7.x2.x3.RESET_B
rlabel metal1 19129 -2654 19247 -2645 1 x7.x2.x3.RESET_B
rlabel metal1 18469 -2654 18599 -2645 1 x7.x2.x3.RESET_B
rlabel metal1 18469 -2682 19247 -2654 1 x7.x2.x3.RESET_B
rlabel metal1 18469 -2691 18599 -2682 1 x7.x2.x3.RESET_B
rlabel metal1 17720 -2886 19836 -2790 1 x7.x2.x3.VGND
rlabel metal1 17720 -2342 19836 -2246 1 x7.x2.x3.VPWR
flabel locali 21682 -2620 21711 -2585 0 FreeSans 200 0 0 0 x7.x2.x4.Q
flabel locali 21984 -2617 22006 -2584 0 FreeSans 200 0 0 0 x7.x2.x4.Q_N
flabel locali 21409 -2685 21443 -2651 0 FreeSans 400 0 0 0 x7.x2.x4.RESET_B
flabel locali 20233 -2549 20267 -2515 0 FreeSans 400 0 0 0 x7.x2.x4.D
flabel locali 19958 -2549 19992 -2515 0 FreeSans 400 0 0 0 x7.x2.x4.CLK
flabel locali 19958 -2617 19992 -2583 0 FreeSans 400 0 0 0 x7.x2.x4.CLK
flabel locali 21409 -2617 21443 -2583 0 FreeSans 400 0 0 0 x7.x2.x4.RESET_B
flabel metal1 19957 -2855 19991 -2821 0 FreeSans 200 0 0 0 x7.x2.x4.VGND
flabel metal1 19957 -2311 19991 -2277 0 FreeSans 200 0 0 0 x7.x2.x4.VPWR
flabel nwell 19957 -2311 19991 -2277 0 FreeSans 200 0 0 0 x7.x2.x4.VPB
flabel pwell 19957 -2855 19991 -2821 0 FreeSans 200 0 0 0 x7.x2.x4.VNB
rlabel comment 19928 -2838 19928 -2838 4 x7.x2.x4.dfrbp_1
rlabel locali 21409 -2711 21457 -2631 1 x7.x2.x4.RESET_B
rlabel locali 21349 -2631 21457 -2557 1 x7.x2.x4.RESET_B
rlabel metal1 21397 -2691 21455 -2682 1 x7.x2.x4.RESET_B
rlabel metal1 21337 -2645 21395 -2582 1 x7.x2.x4.RESET_B
rlabel metal1 21337 -2654 21455 -2645 1 x7.x2.x4.RESET_B
rlabel metal1 20677 -2654 20807 -2645 1 x7.x2.x4.RESET_B
rlabel metal1 20677 -2682 21455 -2654 1 x7.x2.x4.RESET_B
rlabel metal1 20677 -2691 20807 -2682 1 x7.x2.x4.RESET_B
rlabel metal1 19928 -2886 22044 -2790 1 x7.x2.x4.VGND
rlabel metal1 19928 -2342 22044 -2246 1 x7.x2.x4.VPWR
flabel pwell 14989 -2855 15023 -2821 0 FreeSans 200 0 0 0 x7.x2.x1.VNB
flabel nwell 14989 -2311 15023 -2277 0 FreeSans 200 0 0 0 x7.x2.x1.VPB
flabel metal1 14989 -2311 15023 -2277 0 FreeSans 200 0 0 0 x7.x2.x1.VPWR
flabel metal1 14989 -2855 15023 -2821 0 FreeSans 200 0 0 0 x7.x2.x1.VGND
flabel locali 15357 -2413 15391 -2379 0 FreeSans 340 0 0 0 x7.x2.x1.X
flabel locali 15173 -2549 15207 -2515 0 FreeSans 340 0 0 0 x7.x2.x1.B
flabel locali 14989 -2481 15023 -2447 0 FreeSans 340 0 0 0 x7.x2.x1.A
rlabel comment 14960 -2838 14960 -2838 4 x7.x2.x1.and2_0
rlabel metal1 14960 -2886 15420 -2790 1 x7.x2.x1.VGND
rlabel metal1 14960 -2342 15420 -2246 1 x7.x2.x1.VPWR
flabel metal1 17650 -2314 17703 -2285 0 FreeSans 200 0 0 0 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_0.VPWR
flabel metal1 17649 -2856 17700 -2818 0 FreeSans 200 0 0 0 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_0.VGND
rlabel comment 17628 -2838 17628 -2838 4 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_0.tapvpwrvgnd_1
rlabel metal1 17628 -2886 17720 -2790 1 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_0.VGND
rlabel metal1 17628 -2342 17720 -2246 1 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_0.VPWR
flabel metal1 14890 -2314 14943 -2285 0 FreeSans 200 0 0 0 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_1.VPWR
flabel metal1 14889 -2856 14940 -2818 0 FreeSans 200 0 0 0 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_1.VGND
rlabel comment 14868 -2838 14868 -2838 4 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_1.tapvpwrvgnd_1
rlabel metal1 14868 -2886 14960 -2790 1 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_1.VGND
rlabel metal1 14868 -2342 14960 -2246 1 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_1.VPWR
flabel metal1 15442 -2314 15495 -2285 0 FreeSans 200 0 0 0 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_2.VPWR
flabel metal1 15441 -2856 15492 -2818 0 FreeSans 200 0 0 0 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_2.VGND
rlabel comment 15420 -2838 15420 -2838 4 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_2.tapvpwrvgnd_1
rlabel metal1 15420 -2886 15512 -2790 1 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_2.VGND
rlabel metal1 15420 -2342 15512 -2246 1 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_2.VPWR
flabel metal1 19858 -2314 19911 -2285 0 FreeSans 200 0 0 0 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_3.VPWR
flabel metal1 19857 -2856 19908 -2818 0 FreeSans 200 0 0 0 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_3.VGND
rlabel comment 19836 -2838 19836 -2838 4 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_3.tapvpwrvgnd_1
rlabel metal1 19836 -2886 19928 -2790 1 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_3.VGND
rlabel metal1 19836 -2342 19928 -2246 1 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_3.VPWR
flabel metal1 22066 -2314 22119 -2285 0 FreeSans 200 0 0 0 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_4.VPWR
flabel metal1 22065 -2856 22116 -2818 0 FreeSans 200 0 0 0 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_4.VGND
rlabel comment 22044 -2838 22044 -2838 4 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_4.tapvpwrvgnd_1
rlabel metal1 22044 -2886 22136 -2790 1 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_4.VGND
rlabel metal1 22044 -2342 22136 -2246 1 x7.x2.sky130_fd_sc_hd__tapvpwrvgnd_1_4.VPWR
flabel metal1 15220 -2328 16926 -2264 0 FreeSans 800 0 0 0 x7.x1.dvdd
flabel metal1 15202 -1780 16908 -1716 0 FreeSans 800 0 0 0 x7.x1.dvss
flabel metal1 14726 -2112 14826 -2012 0 FreeSans 800 0 0 0 x7.x1.clkin
flabel metal1 14726 -1936 14826 -1836 0 FreeSans 800 0 0 0 x7.x1.ena
flabel space 15350 -2004 15544 -1954 0 FreeSans 400 0 0 0 x7.x1.gated_clk
flabel metal1 15854 -2072 17556 -2040 0 FreeSans 400 0 0 0 x7.x1.Qb1
flabel metal1 18062 -2072 19766 -2040 0 FreeSans 400 0 0 0 x7.x1.Qb2
flabel space 21663 -2066 21729 -1847 0 FreeSans 400 0 0 0 x7.x1.done
flabel metal2 15144 -2212 15244 -1972 0 FreeSans 800 0 0 0 x7.x1.doneb
flabel locali 17266 -2003 17295 -1968 0 FreeSans 200 0 0 0 x7.x1.x2.Q
flabel locali 17568 -2004 17590 -1971 0 FreeSans 200 0 0 0 x7.x1.x2.Q_N
flabel locali 16993 -1937 17027 -1903 0 FreeSans 400 0 0 0 x7.x1.x2.RESET_B
flabel locali 15817 -2073 15851 -2039 0 FreeSans 400 0 0 0 x7.x1.x2.D
flabel locali 15542 -2073 15576 -2039 0 FreeSans 400 0 0 0 x7.x1.x2.CLK
flabel locali 15542 -2005 15576 -1971 0 FreeSans 400 0 0 0 x7.x1.x2.CLK
flabel locali 16993 -2005 17027 -1971 0 FreeSans 400 0 0 0 x7.x1.x2.RESET_B
flabel metal1 15541 -1767 15575 -1733 0 FreeSans 200 0 0 0 x7.x1.x2.VGND
flabel metal1 15541 -2311 15575 -2277 0 FreeSans 200 0 0 0 x7.x1.x2.VPWR
flabel nwell 15541 -2311 15575 -2277 0 FreeSans 200 0 0 0 x7.x1.x2.VPB
flabel pwell 15541 -1767 15575 -1733 0 FreeSans 200 0 0 0 x7.x1.x2.VNB
rlabel comment 15512 -1750 15512 -1750 2 x7.x1.x2.dfrbp_1
rlabel locali 16993 -1957 17041 -1877 5 x7.x1.x2.RESET_B
rlabel locali 16933 -2031 17041 -1957 5 x7.x1.x2.RESET_B
rlabel metal1 16981 -1906 17039 -1897 5 x7.x1.x2.RESET_B
rlabel metal1 16921 -2006 16979 -1943 5 x7.x1.x2.RESET_B
rlabel metal1 16921 -1943 17039 -1934 5 x7.x1.x2.RESET_B
rlabel metal1 16261 -1943 16391 -1934 5 x7.x1.x2.RESET_B
rlabel metal1 16261 -1934 17039 -1906 5 x7.x1.x2.RESET_B
rlabel metal1 16261 -1906 16391 -1897 5 x7.x1.x2.RESET_B
rlabel metal1 15512 -1798 17628 -1702 5 x7.x1.x2.VGND
rlabel metal1 15512 -2342 17628 -2246 5 x7.x1.x2.VPWR
flabel locali 19474 -2003 19503 -1968 0 FreeSans 200 0 0 0 x7.x1.x3.Q
flabel locali 19776 -2004 19798 -1971 0 FreeSans 200 0 0 0 x7.x1.x3.Q_N
flabel locali 19201 -1937 19235 -1903 0 FreeSans 400 0 0 0 x7.x1.x3.RESET_B
flabel locali 18025 -2073 18059 -2039 0 FreeSans 400 0 0 0 x7.x1.x3.D
flabel locali 17750 -2073 17784 -2039 0 FreeSans 400 0 0 0 x7.x1.x3.CLK
flabel locali 17750 -2005 17784 -1971 0 FreeSans 400 0 0 0 x7.x1.x3.CLK
flabel locali 19201 -2005 19235 -1971 0 FreeSans 400 0 0 0 x7.x1.x3.RESET_B
flabel metal1 17749 -1767 17783 -1733 0 FreeSans 200 0 0 0 x7.x1.x3.VGND
flabel metal1 17749 -2311 17783 -2277 0 FreeSans 200 0 0 0 x7.x1.x3.VPWR
flabel nwell 17749 -2311 17783 -2277 0 FreeSans 200 0 0 0 x7.x1.x3.VPB
flabel pwell 17749 -1767 17783 -1733 0 FreeSans 200 0 0 0 x7.x1.x3.VNB
rlabel comment 17720 -1750 17720 -1750 2 x7.x1.x3.dfrbp_1
rlabel locali 19201 -1957 19249 -1877 5 x7.x1.x3.RESET_B
rlabel locali 19141 -2031 19249 -1957 5 x7.x1.x3.RESET_B
rlabel metal1 19189 -1906 19247 -1897 5 x7.x1.x3.RESET_B
rlabel metal1 19129 -2006 19187 -1943 5 x7.x1.x3.RESET_B
rlabel metal1 19129 -1943 19247 -1934 5 x7.x1.x3.RESET_B
rlabel metal1 18469 -1943 18599 -1934 5 x7.x1.x3.RESET_B
rlabel metal1 18469 -1934 19247 -1906 5 x7.x1.x3.RESET_B
rlabel metal1 18469 -1906 18599 -1897 5 x7.x1.x3.RESET_B
rlabel metal1 17720 -1798 19836 -1702 5 x7.x1.x3.VGND
rlabel metal1 17720 -2342 19836 -2246 5 x7.x1.x3.VPWR
flabel locali 21682 -2003 21711 -1968 0 FreeSans 200 0 0 0 x7.x1.x4.Q
flabel locali 21984 -2004 22006 -1971 0 FreeSans 200 0 0 0 x7.x1.x4.Q_N
flabel locali 21409 -1937 21443 -1903 0 FreeSans 400 0 0 0 x7.x1.x4.RESET_B
flabel locali 20233 -2073 20267 -2039 0 FreeSans 400 0 0 0 x7.x1.x4.D
flabel locali 19958 -2073 19992 -2039 0 FreeSans 400 0 0 0 x7.x1.x4.CLK
flabel locali 19958 -2005 19992 -1971 0 FreeSans 400 0 0 0 x7.x1.x4.CLK
flabel locali 21409 -2005 21443 -1971 0 FreeSans 400 0 0 0 x7.x1.x4.RESET_B
flabel metal1 19957 -1767 19991 -1733 0 FreeSans 200 0 0 0 x7.x1.x4.VGND
flabel metal1 19957 -2311 19991 -2277 0 FreeSans 200 0 0 0 x7.x1.x4.VPWR
flabel nwell 19957 -2311 19991 -2277 0 FreeSans 200 0 0 0 x7.x1.x4.VPB
flabel pwell 19957 -1767 19991 -1733 0 FreeSans 200 0 0 0 x7.x1.x4.VNB
rlabel comment 19928 -1750 19928 -1750 2 x7.x1.x4.dfrbp_1
rlabel locali 21409 -1957 21457 -1877 5 x7.x1.x4.RESET_B
rlabel locali 21349 -2031 21457 -1957 5 x7.x1.x4.RESET_B
rlabel metal1 21397 -1906 21455 -1897 5 x7.x1.x4.RESET_B
rlabel metal1 21337 -2006 21395 -1943 5 x7.x1.x4.RESET_B
rlabel metal1 21337 -1943 21455 -1934 5 x7.x1.x4.RESET_B
rlabel metal1 20677 -1943 20807 -1934 5 x7.x1.x4.RESET_B
rlabel metal1 20677 -1934 21455 -1906 5 x7.x1.x4.RESET_B
rlabel metal1 20677 -1906 20807 -1897 5 x7.x1.x4.RESET_B
rlabel metal1 19928 -1798 22044 -1702 5 x7.x1.x4.VGND
rlabel metal1 19928 -2342 22044 -2246 5 x7.x1.x4.VPWR
flabel pwell 14989 -1767 15023 -1733 0 FreeSans 200 0 0 0 x7.x1.x1.VNB
flabel nwell 14989 -2311 15023 -2277 0 FreeSans 200 0 0 0 x7.x1.x1.VPB
flabel metal1 14989 -2311 15023 -2277 0 FreeSans 200 0 0 0 x7.x1.x1.VPWR
flabel metal1 14989 -1767 15023 -1733 0 FreeSans 200 0 0 0 x7.x1.x1.VGND
flabel locali 15357 -2209 15391 -2175 0 FreeSans 340 0 0 0 x7.x1.x1.X
flabel locali 15173 -2073 15207 -2039 0 FreeSans 340 0 0 0 x7.x1.x1.B
flabel locali 14989 -2141 15023 -2107 0 FreeSans 340 0 0 0 x7.x1.x1.A
rlabel comment 14960 -1750 14960 -1750 2 x7.x1.x1.and2_0
rlabel metal1 14960 -1798 15420 -1702 5 x7.x1.x1.VGND
rlabel metal1 14960 -2342 15420 -2246 5 x7.x1.x1.VPWR
flabel metal1 17650 -2303 17703 -2274 0 FreeSans 200 0 0 0 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_0.VPWR
flabel metal1 17649 -1770 17700 -1732 0 FreeSans 200 0 0 0 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_0.VGND
rlabel comment 17628 -1750 17628 -1750 2 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_0.tapvpwrvgnd_1
rlabel metal1 17628 -1798 17720 -1702 5 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_0.VGND
rlabel metal1 17628 -2342 17720 -2246 5 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_0.VPWR
flabel metal1 14890 -2303 14943 -2274 0 FreeSans 200 0 0 0 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_1.VPWR
flabel metal1 14889 -1770 14940 -1732 0 FreeSans 200 0 0 0 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_1.VGND
rlabel comment 14868 -1750 14868 -1750 2 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_1.tapvpwrvgnd_1
rlabel metal1 14868 -1798 14960 -1702 5 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_1.VGND
rlabel metal1 14868 -2342 14960 -2246 5 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_1.VPWR
flabel metal1 15442 -2303 15495 -2274 0 FreeSans 200 0 0 0 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_2.VPWR
flabel metal1 15441 -1770 15492 -1732 0 FreeSans 200 0 0 0 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_2.VGND
rlabel comment 15420 -1750 15420 -1750 2 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_2.tapvpwrvgnd_1
rlabel metal1 15420 -1798 15512 -1702 5 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_2.VGND
rlabel metal1 15420 -2342 15512 -2246 5 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_2.VPWR
flabel metal1 19858 -2303 19911 -2274 0 FreeSans 200 0 0 0 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_3.VPWR
flabel metal1 19857 -1770 19908 -1732 0 FreeSans 200 0 0 0 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_3.VGND
rlabel comment 19836 -1750 19836 -1750 2 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_3.tapvpwrvgnd_1
rlabel metal1 19836 -1798 19928 -1702 5 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_3.VGND
rlabel metal1 19836 -2342 19928 -2246 5 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_3.VPWR
flabel metal1 22066 -2303 22119 -2274 0 FreeSans 200 0 0 0 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_4.VPWR
flabel metal1 22065 -1770 22116 -1732 0 FreeSans 200 0 0 0 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_4.VGND
rlabel comment 22044 -1750 22044 -1750 2 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_4.tapvpwrvgnd_1
rlabel metal1 22044 -1798 22136 -1702 5 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_4.VGND
rlabel metal1 22044 -2342 22136 -2246 5 x7.x1.sky130_fd_sc_hd__tapvpwrvgnd_1_4.VPWR
flabel metal1 3474 -1307 3503 -1254 0 FreeSans 200 0 0 0 ena_buf_tap.VPWR
flabel metal1 2932 -1304 2970 -1253 0 FreeSans 200 0 0 0 ena_buf_tap.VGND
rlabel comment 2950 -1232 2950 -1232 6 ena_buf_tap.tapvpwrvgnd_1
rlabel metal1 2902 -1324 2998 -1232 3 ena_buf_tap.VGND
rlabel metal1 3446 -1324 3542 -1232 3 ena_buf_tap.VPWR
flabel metal1 4827 -1302 4856 -1249 0 FreeSans 200 0 0 0 standby_buf_tap.VPWR
flabel metal1 5360 -1303 5398 -1252 0 FreeSans 200 0 0 0 standby_buf_tap.VGND
rlabel comment 5380 -1324 5380 -1324 2 standby_buf_tap.tapvpwrvgnd_1
rlabel metal1 5332 -1324 5428 -1232 7 standby_buf_tap.VGND
rlabel metal1 4788 -1324 4884 -1232 7 standby_buf_tap.VPWR
flabel metal1 2933 -1389 2967 -1355 0 FreeSans 200 0 0 0 x1.VGND
flabel metal1 3477 -1387 3511 -1353 0 FreeSans 200 0 0 0 x1.VPWR
flabel locali 3477 -1387 3511 -1353 0 FreeSans 200 0 0 0 x1.VPWR
flabel locali 2933 -1389 2967 -1355 0 FreeSans 200 0 0 0 x1.VGND
flabel locali 3035 -1569 3069 -1535 0 FreeSans 200 0 0 0 x1.X
flabel locali 3307 -1569 3341 -1535 0 FreeSans 200 0 0 0 x1.X
flabel locali 3375 -1569 3409 -1535 0 FreeSans 200 0 0 0 x1.X
flabel locali 3171 -1387 3205 -1353 0 FreeSans 200 0 0 0 x1.A
flabel nwell 3477 -1387 3511 -1353 0 FreeSans 200 0 0 0 x1.VPB
flabel pwell 2933 -1389 2967 -1355 0 FreeSans 200 0 0 0 x1.VNB
rlabel comment 2950 -1324 2950 -1324 6 x1.buf_1
rlabel metal1 2902 -1600 2998 -1324 3 x1.VGND
rlabel metal1 3446 -1600 3542 -1324 3 x1.VPWR
flabel metal1 5363 -1389 5397 -1355 0 FreeSans 200 0 0 0 x2.VGND
flabel metal1 4819 -1387 4853 -1353 0 FreeSans 200 0 0 0 x2.VPWR
flabel locali 4819 -1387 4853 -1353 0 FreeSans 200 0 0 0 x2.VPWR
flabel locali 5363 -1389 5397 -1355 0 FreeSans 200 0 0 0 x2.VGND
flabel locali 5261 -1569 5295 -1535 0 FreeSans 200 0 0 0 x2.X
flabel locali 4989 -1569 5023 -1535 0 FreeSans 200 0 0 0 x2.X
flabel locali 4921 -1569 4955 -1535 0 FreeSans 200 0 0 0 x2.X
flabel locali 5125 -1387 5159 -1353 0 FreeSans 200 0 0 0 x2.A
flabel nwell 4819 -1387 4853 -1353 0 FreeSans 200 0 0 0 x2.VPB
flabel pwell 5363 -1389 5397 -1355 0 FreeSans 200 0 0 0 x2.VNB
rlabel comment 5380 -1324 5380 -1324 4 x2.buf_1
rlabel metal1 5332 -1600 5428 -1324 7 x2.VGND
rlabel metal1 4788 -1600 4884 -1324 7 x2.VPWR
<< end >>
