magic
tech sky130A
magscale 1 2
timestamp 1713362978
<< dnwell >>
rect 1926 -9006 6422 -3446
rect 8780 -10312 25248 -4220
rect 1706 -23624 25490 -11618
<< nwell >>
rect 1846 -3652 6502 -3366
rect 1846 -8800 2132 -3652
rect 6216 -8800 6502 -3652
rect 1846 -9086 6502 -8800
rect 8700 -4426 25328 -4140
rect 8700 -10106 8986 -4426
rect 25042 -10106 25328 -4426
rect 8700 -10392 25328 -10106
rect 1626 -11824 25570 -11538
rect 1626 -23418 1912 -11824
rect 25284 -23418 25570 -11824
rect 1626 -23704 25570 -23418
<< pwell >>
rect 10652 -5358 11064 -4958
rect 12592 -5420 12844 -4896
rect 14698 -5358 15110 -4958
<< psubdiff >>
rect 6058 -862 6672 -858
rect 6058 -874 7112 -862
rect 6058 -882 7024 -874
rect 13398 -878 13422 -874
rect 22618 -878 25234 -854
rect 6672 -886 7024 -882
rect 1716 -914 2190 -890
rect 13398 -1614 13422 -1162
rect 1694 -3228 1716 -2904
rect 1694 -3270 1718 -3228
rect 12228 -3358 12252 -3356
rect 6578 -3496 6586 -3472
rect 13778 -3634 13802 -3358
rect 25260 -4056 25284 -3634
rect 12228 -4068 12252 -4056
rect 1668 -11496 1692 -9154
rect 8614 -9164 8626 -9154
rect 8606 -9242 8626 -9164
rect 8602 -10436 8626 -9242
rect 8524 -11500 8548 -11496
rect 25508 -11500 25532 -10436
<< nsubdiff >>
rect 1883 -3423 6465 -3403
rect 1883 -3457 1963 -3423
rect 6385 -3457 6465 -3423
rect 1883 -3477 6465 -3457
rect 1883 -3483 1957 -3477
rect 1883 -8969 1903 -3483
rect 1937 -8969 1957 -3483
rect 1883 -8975 1957 -8969
rect 6391 -3483 6465 -3477
rect 6391 -8969 6411 -3483
rect 6445 -8969 6465 -3483
rect 6391 -8975 6465 -8969
rect 1883 -8995 6465 -8975
rect 1883 -9029 1963 -8995
rect 6385 -9029 6465 -8995
rect 1883 -9049 6465 -9029
rect 8737 -4197 25291 -4177
rect 8737 -4231 8817 -4197
rect 25211 -4231 25291 -4197
rect 8737 -4251 25291 -4231
rect 8737 -4257 8811 -4251
rect 8737 -10275 8757 -4257
rect 8791 -10275 8811 -4257
rect 8737 -10281 8811 -10275
rect 25217 -4257 25291 -4251
rect 25217 -10275 25237 -4257
rect 25271 -10275 25291 -4257
rect 25217 -10281 25291 -10275
rect 8737 -10301 25291 -10281
rect 8737 -10335 8817 -10301
rect 25211 -10335 25291 -10301
rect 8737 -10355 25291 -10335
rect 1663 -11595 25533 -11575
rect 1663 -11629 1743 -11595
rect 25453 -11629 25533 -11595
rect 1663 -11649 25533 -11629
rect 1663 -11655 1737 -11649
rect 1663 -23587 1683 -11655
rect 1717 -23587 1737 -11655
rect 1663 -23593 1737 -23587
rect 25459 -11655 25533 -11649
rect 25459 -23587 25479 -11655
rect 25513 -23587 25533 -11655
rect 25459 -23593 25533 -23587
rect 1663 -23613 25533 -23593
rect 1663 -23647 1743 -23613
rect 25453 -23647 25533 -23613
rect 1663 -23667 25533 -23647
<< psubdiffcont >>
rect 7024 -878 13398 -874
rect 6058 -886 6672 -882
rect 7024 -886 25234 -878
rect 1716 -2904 2190 -914
rect 6058 -1162 25234 -886
rect 6058 -1614 13398 -1162
rect 6058 -2904 7112 -1614
rect 1716 -3228 7112 -2904
rect 1718 -3270 7112 -3228
rect 6578 -3356 7112 -3270
rect 6578 -3358 12228 -3356
rect 6578 -3472 13778 -3358
rect 6586 -3634 13778 -3472
rect 22618 -3634 25234 -1162
rect 6586 -4056 25260 -3634
rect 6586 -4068 12228 -4056
rect 6586 -9154 8614 -4068
rect 1692 -9164 8614 -9154
rect 1692 -9242 8606 -9164
rect 1692 -10436 8602 -9242
rect 1692 -11496 25508 -10436
rect 8548 -11500 25508 -11496
<< nsubdiffcont >>
rect 1963 -3457 6385 -3423
rect 1903 -8969 1937 -3483
rect 6411 -8969 6445 -3483
rect 1963 -9029 6385 -8995
rect 8817 -4231 25211 -4197
rect 8757 -10275 8791 -4257
rect 25237 -10275 25271 -4257
rect 8817 -10335 25211 -10301
rect 1743 -11629 25453 -11595
rect 1683 -23587 1717 -11655
rect 25479 -23587 25513 -11655
rect 1743 -23647 25453 -23613
<< locali >>
rect 2748 -864 2806 -850
rect 1716 -914 2190 -898
rect 5530 -884 5586 -850
rect 3146 -956 3246 -946
rect 3018 -1182 3046 -1128
rect 3146 -1180 3156 -956
rect 3236 -1180 3246 -956
rect 3146 -1194 3246 -1180
rect 5086 -958 5186 -948
rect 5086 -1180 5096 -958
rect 5176 -1180 5186 -958
rect 5290 -1180 5316 -1126
rect 6058 -870 6672 -866
rect 6058 -874 7112 -870
rect 6058 -882 7024 -874
rect 13398 -878 13414 -874
rect 22618 -878 25234 -862
rect 6672 -886 7024 -882
rect 5086 -1192 5186 -1180
rect 3146 -1358 3210 -1194
rect 5120 -1350 5184 -1192
rect 1702 -3228 1716 -2904
rect 3038 -1694 3426 -1564
rect 3038 -1768 3050 -1694
rect 3412 -1768 3426 -1694
rect 3038 -1780 3426 -1768
rect 4904 -1686 5292 -1556
rect 4904 -1760 4916 -1686
rect 5278 -1760 5292 -1686
rect 4904 -1772 5292 -1760
rect 13398 -1614 13414 -1162
rect 1702 -3270 1718 -3228
rect 6406 -3417 6446 -3416
rect 1905 -3423 6446 -3417
rect 1903 -3457 1963 -3423
rect 6385 -3452 6446 -3423
rect 6385 -3457 6445 -3452
rect 1903 -3483 1943 -3457
rect 1937 -5100 1943 -3483
rect 6407 -3483 6445 -3457
rect 1937 -5154 2644 -5100
rect 6407 -5104 6411 -3483
rect 1937 -6772 1990 -5154
rect 2476 -6772 2644 -5154
rect 5692 -5156 6411 -5104
rect 5692 -6428 5838 -5156
rect 4762 -6434 5838 -6428
rect 3706 -6560 5838 -6434
rect 1937 -6822 2644 -6772
rect 3634 -6774 5838 -6560
rect 6324 -6774 6411 -5156
rect 1937 -8969 1943 -6822
rect 2128 -7064 3504 -6958
rect 2130 -7250 2336 -7064
rect 2496 -7126 3228 -7116
rect 2496 -7214 2510 -7126
rect 2130 -7254 2482 -7250
rect 2130 -7266 2526 -7254
rect 2130 -8042 2420 -7266
rect 2512 -8042 2526 -7266
rect 2130 -8054 2526 -8042
rect 2564 -7266 2684 -7254
rect 2564 -8042 2578 -7266
rect 2670 -8042 2684 -7266
rect 2564 -8054 2684 -8042
rect 2722 -7266 2842 -7254
rect 2722 -8042 2736 -7266
rect 2828 -8042 2842 -7266
rect 2722 -8054 2842 -8042
rect 2880 -7266 3000 -7254
rect 2880 -8042 2894 -7266
rect 2986 -8042 3000 -7266
rect 2880 -8054 3000 -8042
rect 3036 -7266 3156 -7254
rect 3036 -8042 3050 -7266
rect 3142 -8042 3156 -7266
rect 3036 -8054 3156 -8042
rect 3196 -7266 3316 -7254
rect 3196 -8042 3210 -7266
rect 3302 -8042 3316 -7266
rect 3196 -8054 3316 -8042
rect 2130 -8058 2482 -8054
rect 2130 -8250 2336 -8058
rect 2496 -8172 2512 -8092
rect 3212 -8172 3228 -8092
rect 2496 -8184 3228 -8172
rect 3408 -8250 3504 -7064
rect 2130 -8812 3504 -8250
rect 3634 -7050 6411 -6774
rect 3634 -8254 3708 -7050
rect 3872 -7120 4600 -7110
rect 3872 -7208 3888 -7120
rect 4588 -7208 4600 -7120
rect 4762 -7252 6411 -7050
rect 4616 -7254 6411 -7252
rect 3782 -7266 3902 -7254
rect 3782 -8044 3796 -7266
rect 3888 -8044 3902 -7266
rect 3782 -8054 3902 -8044
rect 3940 -7266 4060 -7254
rect 3940 -8044 3954 -7266
rect 4046 -8044 4060 -7266
rect 3940 -8054 4060 -8044
rect 4098 -7266 4218 -7254
rect 4098 -8044 4112 -7266
rect 4204 -8044 4218 -7266
rect 4098 -8054 4218 -8044
rect 4256 -7266 4376 -7254
rect 4256 -8044 4270 -7266
rect 4362 -8044 4376 -7266
rect 4256 -8054 4376 -8044
rect 4414 -7266 4534 -7254
rect 4414 -8044 4428 -7266
rect 4520 -8044 4534 -7266
rect 4414 -8054 4534 -8044
rect 4572 -7266 6411 -7254
rect 4572 -8044 4586 -7266
rect 4678 -8044 6411 -7266
rect 4572 -8054 6411 -8044
rect 4616 -8060 6411 -8054
rect 3872 -8188 3888 -8102
rect 4594 -8188 4608 -8102
rect 3872 -8196 4608 -8188
rect 4762 -8254 6411 -8060
rect 2130 -8814 3468 -8812
rect 1903 -8988 1943 -8969
rect 3634 -8969 6411 -8254
rect 7506 -2082 9044 -2072
rect 7506 -2128 7514 -2082
rect 9032 -2128 9044 -2082
rect 7506 -2140 9044 -2128
rect 9428 -2092 10970 -2086
rect 9428 -2140 9438 -2092
rect 10952 -2140 10970 -2092
rect 9428 -2154 10970 -2140
rect 12600 -2156 13048 -2092
rect 11300 -2180 11474 -2164
rect 7378 -2188 7492 -2184
rect 7378 -2198 7552 -2188
rect 7378 -2976 7444 -2198
rect 7540 -2976 7552 -2198
rect 7378 -2988 7552 -2976
rect 7592 -2198 7712 -2188
rect 7592 -2976 7604 -2198
rect 7700 -2976 7712 -2198
rect 7592 -2988 7712 -2976
rect 7750 -2198 7870 -2188
rect 7750 -2976 7762 -2198
rect 7858 -2976 7870 -2198
rect 7750 -2988 7870 -2976
rect 7908 -2198 8028 -2188
rect 7908 -2976 7920 -2198
rect 8016 -2976 8028 -2198
rect 7908 -2988 8028 -2976
rect 8066 -2198 8186 -2188
rect 8066 -2976 8078 -2198
rect 8174 -2976 8186 -2198
rect 8066 -2988 8186 -2976
rect 8222 -2198 8342 -2186
rect 8222 -2976 8234 -2198
rect 8330 -2976 8342 -2198
rect 8222 -2986 8342 -2976
rect 8380 -2198 8500 -2188
rect 8380 -2976 8392 -2198
rect 8488 -2976 8500 -2198
rect 8380 -2988 8500 -2976
rect 8540 -2198 8660 -2186
rect 9072 -2188 9186 -2186
rect 8540 -2976 8552 -2198
rect 8648 -2976 8660 -2198
rect 8540 -2986 8660 -2976
rect 8696 -2198 8816 -2188
rect 8696 -2976 8708 -2198
rect 8804 -2976 8816 -2198
rect 8696 -2988 8816 -2976
rect 8854 -2198 8974 -2188
rect 8854 -2976 8866 -2198
rect 8962 -2976 8974 -2198
rect 8854 -2988 8974 -2976
rect 9012 -2198 9186 -2188
rect 9012 -2976 9024 -2198
rect 9120 -2976 9186 -2198
rect 9012 -2988 9186 -2976
rect 9072 -2990 9186 -2988
rect 9306 -2192 9420 -2190
rect 11000 -2192 11114 -2190
rect 9306 -2202 9478 -2192
rect 9306 -2980 9370 -2202
rect 9466 -2980 9478 -2202
rect 9306 -2992 9478 -2980
rect 9516 -2202 9636 -2192
rect 9516 -2980 9528 -2202
rect 9624 -2980 9636 -2202
rect 9516 -2992 9636 -2980
rect 9676 -2202 9796 -2192
rect 9676 -2980 9688 -2202
rect 9784 -2980 9796 -2202
rect 9676 -2992 9796 -2980
rect 9834 -2202 9954 -2192
rect 9834 -2980 9846 -2202
rect 9942 -2980 9954 -2202
rect 9834 -2992 9954 -2980
rect 9990 -2202 10110 -2192
rect 9990 -2980 10002 -2202
rect 10098 -2980 10110 -2202
rect 9990 -2992 10110 -2980
rect 10150 -2202 10270 -2192
rect 10150 -2980 10162 -2202
rect 10258 -2980 10270 -2202
rect 10150 -2992 10270 -2980
rect 10306 -2202 10426 -2192
rect 10306 -2980 10318 -2202
rect 10414 -2980 10426 -2202
rect 10306 -2992 10426 -2980
rect 10464 -2202 10584 -2192
rect 10464 -2980 10476 -2202
rect 10572 -2980 10584 -2202
rect 10464 -2992 10584 -2980
rect 10624 -2202 10744 -2192
rect 10624 -2980 10636 -2202
rect 10732 -2980 10744 -2202
rect 10624 -2992 10744 -2980
rect 10780 -2202 10900 -2192
rect 10780 -2980 10792 -2202
rect 10888 -2980 10900 -2202
rect 10780 -2992 10900 -2980
rect 10938 -2202 11114 -2192
rect 10938 -2980 10950 -2202
rect 11046 -2980 11114 -2202
rect 11300 -2958 11310 -2180
rect 11468 -2958 11474 -2180
rect 11300 -2974 11474 -2958
rect 11592 -2182 11678 -2170
rect 11592 -2956 11606 -2182
rect 11666 -2956 11678 -2182
rect 12600 -2212 12634 -2156
rect 12770 -2212 12878 -2156
rect 13014 -2212 13048 -2156
rect 11592 -2968 11678 -2956
rect 13030 -2468 13668 -2446
rect 10938 -2992 11114 -2980
rect 9306 -2994 9420 -2992
rect 11000 -2994 11114 -2992
rect 13030 -3026 13052 -2468
rect 13648 -3026 13668 -2468
rect 7502 -3046 9044 -3034
rect 7502 -3092 7512 -3046
rect 9034 -3092 9044 -3046
rect 7502 -3102 9044 -3092
rect 9426 -3044 10970 -3030
rect 9426 -3092 9436 -3044
rect 10952 -3092 10970 -3044
rect 9426 -3098 10970 -3092
rect 13030 -3190 13668 -3026
rect 12440 -3216 13668 -3190
rect 12228 -3358 12244 -3356
rect 12440 -3358 12462 -3216
rect 12588 -3358 13668 -3216
rect 16104 -3004 16222 -2992
rect 6578 -3488 6586 -3472
rect 1902 -8989 1944 -8988
rect 3634 -8989 6445 -8969
rect 1902 -8995 6445 -8989
rect 1902 -9029 1963 -8995
rect 6385 -9029 6445 -8995
rect 1902 -9030 1944 -9029
rect 13778 -3634 13794 -3358
rect 16104 -3422 16120 -3004
rect 15008 -3442 16120 -3422
rect 16212 -3438 16222 -3004
rect 15008 -3516 15034 -3442
rect 16212 -3516 16220 -3438
rect 15008 -3534 16220 -3516
rect 25260 -4056 25276 -3634
rect 12228 -4068 12244 -4056
rect 1676 -11496 1692 -9154
rect 8757 -4231 8817 -4197
rect 25211 -4231 25271 -4197
rect 8757 -4257 8791 -4231
rect 8614 -9164 8618 -9154
rect 8606 -9242 8618 -9164
rect 8602 -10436 8618 -9242
rect 25237 -4257 25271 -4231
rect 8880 -4316 25158 -4298
rect 8791 -5608 8792 -5450
rect 8880 -5476 8900 -4316
rect 11694 -4734 12058 -4548
rect 10462 -4750 12058 -4734
rect 16094 -4556 16958 -4548
rect 17330 -4556 18192 -4548
rect 16094 -4582 18192 -4556
rect 10462 -4768 15282 -4750
rect 10462 -4958 10494 -4768
rect 11436 -4958 12014 -4818
rect 12592 -4958 12844 -4816
rect 13748 -4958 14326 -4818
rect 15264 -4958 15282 -4768
rect 10462 -4970 11230 -4958
rect 11224 -5346 11230 -4970
rect 10462 -5358 11230 -5346
rect 11436 -5354 11452 -4958
rect 11992 -5354 12014 -4958
rect 10462 -5476 10494 -5358
rect 8880 -5494 10494 -5476
rect 11436 -5500 12014 -5354
rect 12104 -4970 12504 -4958
rect 12104 -5346 12122 -4970
rect 12488 -5346 12504 -4970
rect 12104 -5358 12504 -5346
rect 12592 -5358 12604 -4958
rect 12826 -5358 12844 -4958
rect 12918 -4970 13178 -4958
rect 12918 -5346 12924 -4970
rect 13168 -5346 13178 -4970
rect 12918 -5358 13178 -5346
rect 13260 -4970 13660 -4958
rect 13260 -5346 13276 -4970
rect 13642 -5346 13660 -4970
rect 13260 -5358 13660 -5346
rect 13748 -5354 13768 -4958
rect 14308 -5354 14326 -4958
rect 12592 -5500 12844 -5358
rect 13748 -5500 14326 -5354
rect 14532 -4970 15282 -4958
rect 14532 -5346 14538 -4970
rect 14532 -5358 15282 -5346
rect 15264 -5530 15282 -5358
rect 16094 -5530 16118 -4582
rect 16260 -4700 18034 -4640
rect 16648 -4734 16924 -4700
rect 15264 -5548 16118 -5530
rect 16210 -4744 16924 -4734
rect 16210 -4794 16666 -4744
rect 16210 -5484 16228 -4794
rect 16210 -5530 16666 -5484
rect 16878 -5530 16924 -4744
rect 16210 -5542 16924 -5530
rect 17026 -4750 17266 -4734
rect 17026 -5526 17044 -4750
rect 17246 -5526 17266 -4750
rect 17026 -5542 17266 -5526
rect 17498 -4750 18082 -4734
rect 17498 -5526 17514 -4750
rect 18064 -5526 18082 -4750
rect 17498 -5542 18082 -5526
rect 16648 -5576 16924 -5542
rect 8791 -5636 16060 -5608
rect 16260 -5636 18034 -5576
rect 8791 -5640 15260 -5636
rect 8791 -7366 8878 -5640
rect 15938 -5752 16060 -5636
rect 18174 -5674 18192 -4582
rect 21246 -5244 22086 -5218
rect 18848 -5382 20732 -5352
rect 18848 -5530 18878 -5382
rect 18848 -5548 18904 -5530
rect 18174 -5694 18808 -5674
rect 15938 -5758 18742 -5752
rect 16602 -5762 18742 -5758
rect 10492 -5814 15260 -5776
rect 10492 -5988 10540 -5814
rect 10682 -5948 15086 -5888
rect 15230 -5894 15260 -5814
rect 16602 -5888 16776 -5762
rect 17510 -5886 17700 -5762
rect 18728 -5850 18742 -5762
rect 18788 -5790 18808 -5694
rect 18862 -5790 18904 -5548
rect 20690 -5776 20732 -5382
rect 21246 -5402 21272 -5244
rect 21246 -5486 21400 -5402
rect 21214 -5508 21400 -5486
rect 21214 -5776 21272 -5508
rect 20690 -5790 21272 -5776
rect 18788 -5808 18904 -5790
rect 18728 -5864 21204 -5850
rect 20504 -5870 21204 -5864
rect 17510 -5888 18330 -5886
rect 11088 -5988 11248 -5984
rect 10492 -6000 11248 -5988
rect 11242 -6378 11248 -6000
rect 10492 -6388 11248 -6378
rect 10492 -6518 10540 -6388
rect 11088 -6394 11248 -6388
rect 11362 -6430 11542 -5948
rect 11588 -6000 11892 -5984
rect 11588 -6378 11602 -6000
rect 11878 -6378 11892 -6000
rect 11588 -6394 11892 -6378
rect 11936 -6430 12116 -5948
rect 12912 -5982 13260 -5948
rect 12164 -6000 12850 -5984
rect 12164 -6378 12176 -6000
rect 12452 -6378 12850 -6000
rect 12164 -6394 12850 -6378
rect 12912 -6392 12924 -5982
rect 13252 -6392 13260 -5982
rect 12912 -6430 13260 -6392
rect 13300 -6000 13604 -5984
rect 13300 -6378 13316 -6000
rect 13592 -6378 13604 -6000
rect 13300 -6394 13604 -6378
rect 13650 -6430 13830 -5948
rect 13874 -6000 14178 -5984
rect 13874 -6378 13886 -6000
rect 14162 -6378 14178 -6000
rect 13874 -6394 14178 -6378
rect 14222 -6430 14402 -5948
rect 14520 -5988 14680 -5984
rect 15228 -5988 15260 -5894
rect 14520 -6000 15260 -5988
rect 15938 -5894 18330 -5888
rect 14520 -6378 14526 -6000
rect 14520 -6388 15260 -6378
rect 14520 -6394 14680 -6388
rect 10682 -6476 15086 -6430
rect 11088 -6518 11248 -6512
rect 10492 -6528 11248 -6518
rect 11242 -6906 11248 -6528
rect 10492 -6918 11248 -6906
rect 10492 -7080 10540 -6918
rect 11088 -6922 11248 -6918
rect 11362 -6958 11542 -6476
rect 11586 -6528 11890 -6512
rect 11586 -6906 11602 -6528
rect 11878 -6906 11890 -6528
rect 11586 -6922 11890 -6906
rect 11936 -6958 12116 -6476
rect 12160 -6528 12464 -6512
rect 12160 -6530 12238 -6528
rect 12388 -6530 12464 -6528
rect 12160 -6908 12174 -6530
rect 12450 -6908 12464 -6530
rect 12160 -6922 12464 -6908
rect 12508 -6958 12688 -6476
rect 12730 -6528 13034 -6512
rect 12730 -6906 12742 -6528
rect 13018 -6906 13034 -6528
rect 12730 -6922 13034 -6906
rect 13080 -6958 13260 -6476
rect 13304 -6528 13608 -6512
rect 13304 -6906 13316 -6528
rect 13592 -6906 13608 -6528
rect 13304 -6922 13608 -6906
rect 13650 -6958 13830 -6476
rect 13876 -6528 14180 -6512
rect 13876 -6906 13888 -6528
rect 14164 -6906 14180 -6528
rect 13876 -6922 14180 -6906
rect 14222 -6958 14402 -6476
rect 14522 -6518 14682 -6512
rect 15228 -6518 15260 -6388
rect 14522 -6528 15260 -6518
rect 14522 -6906 14526 -6528
rect 14522 -6918 15260 -6906
rect 14522 -6922 14682 -6918
rect 10682 -7018 15086 -6958
rect 10492 -7088 10764 -7080
rect 10492 -7096 10766 -7088
rect 15228 -7096 15260 -6918
rect 10492 -7114 15260 -7096
rect 15938 -7096 16104 -5894
rect 16156 -5956 17118 -5950
rect 16156 -5960 16770 -5956
rect 16156 -6050 16162 -5960
rect 16608 -6050 16770 -5960
rect 17066 -6050 17118 -5956
rect 17176 -5956 18138 -5950
rect 17176 -6050 17228 -5956
rect 17524 -5960 18138 -5956
rect 17524 -6050 17686 -5960
rect 18132 -6050 18138 -5960
rect 16208 -6108 16770 -6092
rect 16208 -6886 16224 -6108
rect 16758 -6886 16770 -6108
rect 16208 -6902 16770 -6886
rect 16998 -6106 17298 -6092
rect 16998 -6890 17014 -6106
rect 17280 -6890 17298 -6106
rect 16998 -6902 17298 -6890
rect 17520 -6108 18082 -6092
rect 17520 -6886 17532 -6108
rect 18066 -6886 18082 -6108
rect 17520 -6902 18082 -6886
rect 16156 -7034 16162 -6944
rect 17078 -7034 17118 -6944
rect 16156 -7044 17118 -7034
rect 17176 -7034 17216 -6944
rect 18132 -7034 18138 -6944
rect 17176 -7044 18138 -7034
rect 18200 -7096 18330 -5894
rect 20504 -6354 20736 -5870
rect 18834 -6382 20736 -6354
rect 18834 -6814 18892 -6382
rect 20670 -6814 20736 -6382
rect 21184 -5924 21204 -5870
rect 22012 -5852 22086 -5244
rect 23274 -5322 23778 -5298
rect 23274 -5404 23294 -5322
rect 23376 -5404 23642 -5322
rect 23724 -5404 23778 -5322
rect 23274 -5406 23278 -5404
rect 22816 -5758 23278 -5406
rect 23756 -5424 23778 -5404
rect 22638 -5788 23278 -5758
rect 23742 -5788 23778 -5424
rect 22638 -5834 23778 -5788
rect 25134 -5834 25158 -4316
rect 22638 -5852 25158 -5834
rect 22012 -5872 25158 -5852
rect 23754 -5874 25158 -5872
rect 21184 -5946 25237 -5924
rect 21184 -5948 24312 -5946
rect 21184 -6224 22398 -5948
rect 21184 -6242 22118 -6224
rect 21184 -6580 21272 -6242
rect 22012 -6308 22118 -6242
rect 18834 -6844 20736 -6814
rect 21202 -6636 21272 -6580
rect 21202 -6742 21400 -6636
rect 21202 -6902 21272 -6742
rect 22010 -6902 22118 -6308
rect 22620 -6246 24312 -5948
rect 22620 -6310 24114 -6246
rect 22620 -6694 22962 -6310
rect 24096 -6686 24114 -6310
rect 22930 -6760 22962 -6694
rect 22930 -6776 22982 -6760
rect 23332 -6774 23730 -6686
rect 24080 -6774 24114 -6686
rect 23332 -6776 24114 -6774
rect 22930 -6802 24114 -6776
rect 25178 -6802 25237 -5946
rect 21202 -6930 22118 -6902
rect 15938 -7114 18330 -7096
rect 25180 -7248 25237 -6802
rect 21202 -7250 25237 -7248
rect 10008 -7270 25237 -7250
rect 10008 -7366 10078 -7270
rect 8791 -7438 10078 -7366
rect 8791 -7454 9648 -7438
rect 9792 -7454 9902 -7438
rect 10046 -7454 10078 -7438
rect 9736 -7570 9952 -7552
rect 8920 -7608 9068 -7586
rect 8920 -10142 8940 -7608
rect 9046 -9422 9068 -7608
rect 9150 -7774 9366 -7684
rect 9150 -9240 9208 -7774
rect 9304 -9240 9366 -7774
rect 9736 -9050 9788 -7570
rect 9904 -9050 9952 -7570
rect 9736 -9136 9952 -9050
rect 10146 -9088 10510 -7380
rect 24760 -7404 25152 -7368
rect 10618 -7674 11048 -7438
rect 10620 -8006 11050 -7770
rect 24220 -7840 24650 -7604
rect 10620 -8338 11050 -8102
rect 24220 -8172 24650 -7936
rect 10620 -8670 11050 -8434
rect 24220 -8502 24650 -8266
rect 10620 -9002 11050 -8766
rect 24220 -8834 24650 -8598
rect 9150 -9268 9366 -9240
rect 10146 -9386 10162 -9088
rect 9208 -9388 9308 -9386
rect 9204 -9422 9312 -9388
rect 9448 -9408 10162 -9386
rect 9448 -9422 9466 -9408
rect 9046 -9442 9466 -9422
rect 10362 -9486 10510 -9088
rect 10620 -9334 11050 -9098
rect 24220 -9166 24650 -8930
rect 10362 -9940 10506 -9486
rect 10620 -9664 11050 -9428
rect 24220 -9500 24650 -9264
rect 24220 -9832 24650 -9596
rect 24760 -9940 24788 -7404
rect 10362 -9960 24788 -9940
rect 25116 -10142 25152 -7404
rect 8920 -10176 25152 -10142
rect 8757 -10301 8791 -10275
rect 25237 -10301 25271 -10275
rect 8757 -10335 8817 -10301
rect 25211 -10335 25271 -10301
rect 8532 -11500 8548 -11496
rect 25508 -11500 25524 -10436
rect 1662 -11588 1786 -11576
rect 1662 -23656 1674 -11588
rect 1772 -11595 1786 -11588
rect 25453 -11629 25513 -11595
rect 1772 -23544 1786 -11629
rect 22120 -11655 25513 -11629
rect 22120 -11668 25479 -11655
rect 1844 -11798 21916 -11756
rect 1844 -11824 7814 -11798
rect 1844 -13814 1996 -11824
rect 7070 -12034 7814 -11824
rect 7070 -12056 13436 -12034
rect 7070 -12246 7164 -12056
rect 7688 -12118 13436 -12056
rect 7070 -12454 7314 -12246
rect 7688 -12304 8232 -12118
rect 13348 -12194 13436 -12118
rect 7688 -12400 8256 -12304
rect 8336 -12322 9886 -12264
rect 8336 -12382 8348 -12322
rect 9840 -12382 9886 -12322
rect 7070 -12642 7164 -12454
rect 7688 -12584 8232 -12400
rect 8336 -12442 9886 -12382
rect 13348 -12510 20656 -12194
rect 13348 -12584 13436 -12510
rect 7688 -12642 13436 -12584
rect 7070 -12680 13436 -12642
rect 20150 -12646 20656 -12510
rect 21870 -12646 21916 -11798
rect 7070 -12862 7778 -12680
rect 20150 -12752 21916 -12646
rect 2982 -12898 7778 -12862
rect 2982 -12988 19070 -12898
rect 2982 -13422 3022 -12988
rect 18502 -13098 19070 -12988
rect 19808 -13098 21916 -12752
rect 3134 -13314 3566 -13098
rect 18502 -13154 21916 -13098
rect 19076 -13190 21916 -13154
rect 19076 -13422 19874 -13190
rect 19994 -13242 21712 -13228
rect 19994 -13244 20918 -13242
rect 19994 -13352 20008 -13244
rect 20788 -13286 20918 -13244
rect 20788 -13352 20802 -13286
rect 19994 -13368 20802 -13352
rect 20904 -13350 20918 -13286
rect 21698 -13350 21712 -13242
rect 20904 -13368 21712 -13350
rect 2982 -13538 19874 -13422
rect 19328 -13814 19874 -13538
rect 19924 -13452 21780 -13426
rect 19924 -13600 19998 -13452
rect 20798 -13600 20908 -13452
rect 21708 -13600 21780 -13452
rect 19924 -13626 21780 -13600
rect 1844 -13926 19874 -13814
rect 19994 -13702 20802 -13680
rect 19994 -13870 20010 -13702
rect 20786 -13760 20802 -13702
rect 20904 -13700 21712 -13680
rect 20904 -13760 20920 -13700
rect 20786 -13800 20920 -13760
rect 21696 -13800 21712 -13700
rect 20786 -13820 21712 -13800
rect 21816 -13746 21916 -13190
rect 22120 -12538 22152 -11668
rect 22120 -12714 24616 -12538
rect 21816 -13758 21956 -13746
rect 20786 -13870 20802 -13820
rect 19994 -13896 20204 -13870
rect 1844 -18014 2018 -13926
rect 2132 -14254 2564 -14038
rect 2134 -14584 2566 -14368
rect 18932 -14418 19364 -14202
rect 2132 -14916 2564 -14700
rect 18932 -14750 19364 -14534
rect 2132 -15248 2564 -15032
rect 18932 -15082 19364 -14866
rect 19474 -15014 19874 -13926
rect 20174 -14308 20204 -13896
rect 19994 -14336 20204 -14308
rect 20622 -13896 20802 -13870
rect 20622 -14308 20654 -13896
rect 20904 -13952 20920 -13856
rect 21696 -13952 21712 -13856
rect 20904 -13966 21712 -13952
rect 21816 -13874 21828 -13758
rect 21944 -13874 21956 -13758
rect 21816 -13886 21956 -13874
rect 20854 -14052 21764 -14008
rect 20854 -14308 20916 -14052
rect 21698 -14308 21764 -14052
rect 20622 -14336 20802 -14308
rect 20854 -14330 21764 -14308
rect 19994 -14500 20010 -14336
rect 20786 -14384 20802 -14336
rect 20786 -14404 21712 -14384
rect 20786 -14444 20920 -14404
rect 20786 -14500 20802 -14444
rect 19994 -14524 20802 -14500
rect 20904 -14504 20920 -14444
rect 21696 -14504 21712 -14404
rect 20904 -14524 21712 -14504
rect 19926 -14600 21782 -14576
rect 19926 -14602 20908 -14600
rect 19926 -14750 19998 -14602
rect 20798 -14748 20908 -14602
rect 21708 -14748 21782 -14600
rect 20798 -14750 21782 -14748
rect 19926 -14776 21782 -14750
rect 19994 -14854 20802 -14838
rect 19994 -14962 20008 -14854
rect 20788 -14920 20802 -14854
rect 20904 -14854 21712 -14838
rect 20904 -14920 20920 -14854
rect 20788 -14962 20920 -14920
rect 21700 -14962 21712 -14854
rect 19994 -14978 21712 -14962
rect 21816 -15014 21916 -13886
rect 2130 -15578 2562 -15362
rect 18932 -15414 19364 -15198
rect 2132 -15912 2564 -15696
rect 18932 -15746 19364 -15530
rect 19474 -15548 21914 -15014
rect 2132 -16242 2564 -16026
rect 18932 -16078 19364 -15862
rect 2132 -16576 2564 -16360
rect 18932 -16410 19364 -16194
rect 2130 -16908 2562 -16692
rect 18932 -16742 19364 -16526
rect 2130 -17240 2562 -17024
rect 18932 -17074 19364 -16858
rect 2132 -17570 2564 -17354
rect 18932 -17406 19364 -17190
rect 2132 -17904 2564 -17688
rect 18932 -17738 19364 -17522
rect 19474 -18014 19534 -15548
rect 20220 -15932 21532 -15878
rect 20220 -16020 20272 -15932
rect 20222 -17992 20272 -16020
rect 20462 -16008 21266 -15934
rect 20462 -16268 20474 -16008
rect 21252 -16268 21266 -16008
rect 20462 -16284 21266 -16268
rect 21474 -16254 21532 -15932
rect 21862 -16254 21914 -15548
rect 20464 -16332 21264 -16318
rect 20464 -16424 20476 -16332
rect 21252 -16424 21264 -16332
rect 20464 -16436 21264 -16424
rect 20464 -16490 21264 -16476
rect 20464 -16582 20476 -16490
rect 21252 -16582 21264 -16490
rect 20464 -16594 21264 -16582
rect 20464 -16648 21264 -16634
rect 20464 -16740 20476 -16648
rect 21252 -16740 21264 -16648
rect 20464 -16752 21264 -16740
rect 20464 -16806 21264 -16792
rect 20464 -16898 20476 -16806
rect 21252 -16898 21264 -16806
rect 20464 -16910 21264 -16898
rect 20464 -16964 21264 -16950
rect 20464 -17056 20476 -16964
rect 21252 -17056 21264 -16964
rect 20464 -17068 21264 -17056
rect 20464 -17122 21264 -17108
rect 20464 -17214 20476 -17122
rect 21252 -17214 21264 -17122
rect 20464 -17226 21264 -17214
rect 20464 -17280 21264 -17266
rect 20464 -17372 20476 -17280
rect 21252 -17372 21264 -17280
rect 20464 -17384 21264 -17372
rect 20464 -17438 21264 -17424
rect 20464 -17530 20476 -17438
rect 21252 -17530 21264 -17438
rect 20464 -17542 21264 -17530
rect 20464 -17596 21264 -17582
rect 20464 -17688 20476 -17596
rect 21252 -17688 21264 -17596
rect 20464 -17700 21264 -17688
rect 1844 -18128 19534 -18014
rect 20220 -18012 20272 -17992
rect 20462 -17756 21266 -17734
rect 20462 -17996 20472 -17756
rect 20462 -18010 20474 -17996
rect 21252 -18010 21266 -17756
rect 20462 -18012 21266 -18010
rect 21474 -18012 21914 -16254
rect 22120 -15876 22396 -12714
rect 22452 -13486 22554 -12794
rect 22596 -13092 23404 -12714
rect 22596 -13392 22608 -13092
rect 23388 -13138 23404 -13092
rect 23390 -13344 23404 -13138
rect 23388 -13392 23404 -13344
rect 22596 -13402 23404 -13392
rect 23448 -13486 23482 -12794
rect 23524 -13090 24332 -12714
rect 23524 -13390 23538 -13090
rect 24318 -13390 24332 -13090
rect 23524 -13402 24332 -13390
rect 24376 -13486 24478 -12794
rect 22452 -13586 24478 -13486
rect 22452 -14056 22554 -13586
rect 22594 -13668 23402 -13656
rect 22594 -13968 22610 -13668
rect 23390 -13702 23402 -13668
rect 23390 -13942 23404 -13702
rect 23390 -13968 23402 -13942
rect 22594 -13980 23402 -13968
rect 23448 -14056 23482 -13586
rect 23520 -13666 24328 -13656
rect 23520 -13966 23536 -13666
rect 24316 -13702 24328 -13666
rect 24316 -13716 24330 -13702
rect 24318 -13744 24330 -13716
rect 24318 -13898 24332 -13744
rect 24318 -13922 24330 -13898
rect 24316 -13942 24330 -13922
rect 24316 -13966 24328 -13942
rect 23520 -13980 24328 -13966
rect 24376 -14056 24478 -13586
rect 22452 -14156 24478 -14056
rect 22452 -14632 22554 -14156
rect 22596 -14242 23404 -14230
rect 22596 -14542 22608 -14242
rect 23388 -14298 23404 -14242
rect 23390 -14504 23404 -14298
rect 23388 -14542 23404 -14504
rect 22596 -14554 23404 -14542
rect 23448 -14632 23482 -14156
rect 23524 -14238 24332 -14230
rect 23524 -14538 23538 -14238
rect 24318 -14538 24332 -14238
rect 23524 -14554 24332 -14538
rect 24376 -14632 24478 -14156
rect 22452 -14732 24478 -14632
rect 22452 -15560 22554 -14732
rect 22596 -14814 23404 -14802
rect 22596 -14976 22610 -14814
rect 23390 -14976 23404 -14814
rect 22596 -14982 23404 -14976
rect 22598 -15512 23404 -15020
rect 23448 -15560 23482 -14732
rect 22452 -15598 23482 -15560
rect 22452 -15642 22612 -15598
rect 23390 -15642 23482 -15598
rect 23524 -14908 24332 -14894
rect 23524 -15622 23570 -14908
rect 24284 -15622 24332 -14908
rect 23524 -15638 24332 -15622
rect 22120 -16002 22400 -15876
rect 22452 -15914 22610 -15642
rect 23392 -15788 23482 -15642
rect 24376 -15788 24478 -14732
rect 23392 -15888 24478 -15788
rect 23392 -15914 23482 -15888
rect 22452 -15940 23482 -15914
rect 22120 -17820 22396 -16002
rect 22452 -16366 22554 -15940
rect 22596 -15988 23404 -15978
rect 22596 -16288 22610 -15988
rect 23390 -16288 23404 -15988
rect 22596 -16302 23404 -16288
rect 23448 -16366 23482 -15940
rect 23522 -15988 24330 -15978
rect 23522 -16288 23538 -15988
rect 24318 -16056 24330 -15988
rect 24318 -16210 24332 -16056
rect 24318 -16288 24330 -16210
rect 23522 -16302 24330 -16288
rect 24376 -16366 24478 -15888
rect 22452 -16466 24478 -16366
rect 22452 -16940 22554 -16466
rect 22596 -16552 23404 -16540
rect 22596 -16852 22610 -16552
rect 23390 -16852 23404 -16552
rect 22596 -16864 23404 -16852
rect 23448 -16940 23482 -16466
rect 23524 -16552 24332 -16540
rect 23524 -16852 23536 -16552
rect 24316 -16606 24332 -16552
rect 24318 -16812 24332 -16606
rect 24316 -16852 24332 -16812
rect 23524 -16864 24332 -16852
rect 24376 -16940 24478 -16466
rect 22452 -17040 24478 -16940
rect 22452 -17736 22554 -17040
rect 22596 -17138 23404 -17126
rect 22596 -17438 22610 -17138
rect 23390 -17438 23404 -17138
rect 22596 -17820 23404 -17438
rect 23448 -17736 23482 -17040
rect 23524 -17136 24332 -17126
rect 23524 -17436 23538 -17136
rect 24318 -17436 24332 -17136
rect 23524 -17820 24332 -17436
rect 24376 -17736 24478 -17040
rect 24524 -17820 24616 -12714
rect 22120 -17924 24616 -17820
rect 22120 -17984 25228 -17924
rect 1844 -18408 1996 -18128
rect 18346 -18408 18856 -18128
rect 20220 -18184 21914 -18012
rect 20220 -18342 24962 -18184
rect 1844 -18466 19534 -18408
rect 20220 -18466 25068 -18342
rect 1844 -18516 25068 -18466
rect 1844 -22518 2018 -18516
rect 2130 -18518 2564 -18516
rect 24528 -18520 24962 -18516
rect 2130 -18850 2564 -18616
rect 2130 -19184 2564 -18950
rect 24530 -19016 24964 -18782
rect 2130 -19514 2564 -19280
rect 24530 -19348 24964 -19114
rect 2130 -19846 2564 -19612
rect 24530 -19680 24964 -19446
rect 2130 -20180 2564 -19946
rect 24530 -20012 24964 -19778
rect 2130 -20510 2564 -20276
rect 24530 -20344 24964 -20110
rect 2130 -20842 2564 -20608
rect 24530 -20676 24964 -20442
rect 2128 -21174 2562 -20940
rect 24530 -21008 24964 -20774
rect 2130 -21506 2564 -21272
rect 24528 -21342 24962 -21108
rect 2130 -21838 2564 -21604
rect 24530 -21672 24964 -21438
rect 2128 -22170 2562 -21936
rect 24528 -22004 24962 -21770
rect 24528 -22338 24962 -22104
rect 2130 -22518 2564 -22444
rect 24530 -22518 24964 -22442
rect 1844 -22632 25076 -22518
rect 1844 -22708 23876 -22632
rect 25198 -22706 25228 -17984
rect 1844 -22710 21092 -22708
rect 1844 -23440 1890 -22710
rect 20268 -22858 21092 -22710
rect 20268 -23114 20374 -22858
rect 20632 -23114 21092 -22858
rect 21630 -22982 22518 -22708
rect 20268 -23440 21092 -23114
rect 21214 -23158 21226 -23096
rect 21744 -23090 22390 -23068
rect 21744 -23348 21764 -23090
rect 1844 -23486 21092 -23440
rect 1772 -23554 20612 -23544
rect 20600 -23613 20612 -23554
rect 21288 -23598 21764 -23348
rect 22366 -23348 22390 -23090
rect 23054 -22858 23876 -22708
rect 23054 -22982 23484 -22858
rect 23742 -22980 23876 -22858
rect 24040 -22730 25228 -22706
rect 22922 -23160 22928 -23098
rect 24040 -23206 24070 -22730
rect 23168 -23230 24070 -23206
rect 23168 -23348 23578 -23230
rect 22366 -23598 23578 -23348
rect 21288 -23613 23578 -23598
rect 25456 -23587 25479 -11668
rect 25456 -23630 25513 -23587
rect 25453 -23647 25513 -23630
rect 20600 -23656 20612 -23647
rect 1662 -23668 20612 -23656
<< viali >>
rect 2748 -1128 2806 -864
rect 2748 -1182 3018 -1128
rect 3156 -1180 3236 -956
rect 5096 -1180 5176 -958
rect 5530 -1126 5586 -884
rect 5316 -1180 5586 -1126
rect 1782 -2952 2162 -1378
rect 3050 -1768 3412 -1694
rect 4916 -1760 5278 -1686
rect 6110 -896 7000 -890
rect 6110 -1272 7934 -896
rect 8606 -1262 11080 -882
rect 11672 -1138 23756 -914
rect 11672 -1262 13372 -1138
rect 6110 -2952 7000 -1272
rect 12602 -1582 13370 -1262
rect 1782 -3222 7000 -2952
rect 1990 -6772 2476 -5154
rect 5838 -6774 6324 -5156
rect 2510 -7214 3230 -7126
rect 2420 -8042 2512 -7266
rect 2578 -8042 2670 -7266
rect 2736 -8042 2828 -7266
rect 2894 -8042 2986 -7266
rect 3050 -8042 3142 -7266
rect 3210 -8042 3302 -7266
rect 2512 -8172 3212 -8092
rect 3888 -7208 4588 -7120
rect 3796 -8044 3888 -7266
rect 3954 -8044 4046 -7266
rect 4112 -8044 4204 -7266
rect 4270 -8044 4362 -7266
rect 4428 -8044 4520 -7266
rect 4586 -8044 4678 -7266
rect 3888 -8188 4594 -8102
rect 6720 -3434 7000 -3222
rect 7514 -2128 9032 -2082
rect 9438 -2140 10952 -2092
rect 7444 -2976 7540 -2198
rect 7604 -2976 7700 -2198
rect 7762 -2976 7858 -2198
rect 7920 -2976 8016 -2198
rect 8078 -2976 8174 -2198
rect 8234 -2976 8330 -2198
rect 8392 -2976 8488 -2198
rect 8552 -2976 8648 -2198
rect 8708 -2976 8804 -2198
rect 8866 -2976 8962 -2198
rect 9024 -2976 9120 -2198
rect 9370 -2980 9466 -2202
rect 9528 -2980 9624 -2202
rect 9688 -2980 9784 -2202
rect 9846 -2980 9942 -2202
rect 10002 -2980 10098 -2202
rect 10162 -2980 10258 -2202
rect 10318 -2980 10414 -2202
rect 10476 -2980 10572 -2202
rect 10636 -2980 10732 -2202
rect 10792 -2980 10888 -2202
rect 10950 -2980 11046 -2202
rect 11310 -2958 11468 -2180
rect 11606 -2956 11666 -2182
rect 13052 -3026 13648 -2468
rect 7512 -3092 9034 -3046
rect 9436 -3092 10952 -3044
rect 12462 -3358 12588 -3216
rect 12462 -3380 12588 -3358
rect 12222 -3414 12588 -3380
rect 6720 -3470 11294 -3434
rect 12222 -3470 13744 -3414
rect 6720 -3658 13744 -3470
rect 16120 -3442 16212 -3004
rect 15034 -3516 16212 -3442
rect 22662 -3490 23754 -1138
rect 6720 -3948 13814 -3658
rect 6720 -5446 8452 -3948
rect 12318 -4018 13814 -3948
rect 22968 -3976 23752 -3490
rect 24460 -3984 25194 -898
rect 13740 -4020 13814 -4018
rect 6720 -7614 7418 -5446
rect 6720 -9330 8426 -7614
rect 1910 -10544 8428 -9330
rect 8900 -4548 25134 -4316
rect 8900 -4734 11694 -4548
rect 8900 -4970 10462 -4734
rect 12058 -4750 16094 -4548
rect 16958 -4556 17330 -4548
rect 8900 -5346 11224 -4970
rect 8900 -5476 10462 -5346
rect 11452 -5354 11992 -4958
rect 12122 -5346 12488 -4970
rect 12604 -5358 12826 -4958
rect 12924 -5346 13168 -4970
rect 13276 -5346 13642 -4970
rect 13768 -5354 14308 -4958
rect 15282 -4970 16094 -4750
rect 14538 -5346 16094 -4970
rect 15282 -5530 16094 -5346
rect 16666 -4794 16878 -4744
rect 16228 -5484 16878 -4794
rect 16666 -5530 16878 -5484
rect 17044 -5526 17246 -4750
rect 17514 -5526 18064 -4750
rect 15260 -5640 15938 -5636
rect 8878 -5758 15938 -5640
rect 18192 -5218 25134 -4548
rect 18192 -5352 21246 -5218
rect 18192 -5548 18848 -5352
rect 18192 -5674 18862 -5548
rect 8878 -5776 16602 -5758
rect 8878 -6000 10492 -5776
rect 15260 -5888 16602 -5776
rect 16776 -5888 17510 -5762
rect 17700 -5864 18728 -5762
rect 18808 -5790 18862 -5674
rect 20732 -5486 21246 -5352
rect 20732 -5776 21214 -5486
rect 17700 -5886 20504 -5864
rect 8878 -6378 11242 -6000
rect 8878 -6528 10492 -6378
rect 11602 -6378 11878 -6000
rect 12176 -6378 12452 -6000
rect 12924 -6392 13252 -5982
rect 13316 -6378 13592 -6000
rect 13886 -6378 14162 -6000
rect 15260 -6000 15938 -5888
rect 14526 -6378 15938 -6000
rect 8878 -6906 11242 -6528
rect 8878 -7114 10492 -6906
rect 11602 -6906 11878 -6528
rect 12238 -6530 12388 -6528
rect 12174 -6908 12450 -6530
rect 12742 -6906 13018 -6528
rect 13316 -6906 13592 -6528
rect 13888 -6906 14164 -6528
rect 15260 -6528 15938 -6378
rect 14526 -6906 15938 -6528
rect 15260 -7114 15938 -6906
rect 16162 -6050 16608 -5960
rect 16770 -6050 17066 -5956
rect 17228 -6050 17524 -5956
rect 17686 -6050 18132 -5960
rect 16224 -6886 16758 -6108
rect 17014 -6890 17280 -6106
rect 17532 -6886 18066 -6108
rect 16162 -7034 17078 -6944
rect 17216 -7034 18132 -6944
rect 18330 -6354 20504 -5886
rect 18330 -6844 18834 -6354
rect 20736 -6580 21184 -5870
rect 22086 -5298 25134 -5218
rect 22086 -5406 23274 -5298
rect 22086 -5758 22816 -5406
rect 22086 -5852 22638 -5758
rect 23778 -5834 25134 -5298
rect 22398 -6224 22620 -5948
rect 20736 -6844 21202 -6580
rect 18330 -6930 21202 -6844
rect 22118 -6694 22620 -6224
rect 24312 -6246 25178 -5946
rect 22118 -6802 22930 -6694
rect 24114 -6802 25178 -6246
rect 22118 -6930 25180 -6802
rect 18330 -7114 25180 -6930
rect 8878 -7248 25180 -7114
rect 8878 -7250 21202 -7248
rect 8878 -7366 10008 -7250
rect 8940 -9442 9046 -7608
rect 9208 -9240 9304 -7774
rect 9788 -9050 9904 -7570
rect 10162 -9408 10362 -9088
rect 9466 -9442 10362 -9408
rect 8940 -9960 10362 -9442
rect 24788 -9960 25116 -7404
rect 8940 -10142 25116 -9960
rect 1910 -11092 15780 -10544
rect 1910 -11096 8428 -11092
rect 1674 -11595 1772 -11588
rect 1674 -11629 1743 -11595
rect 1743 -11629 1772 -11595
rect 1674 -11655 1772 -11629
rect 1674 -23587 1683 -11655
rect 1683 -23587 1717 -11655
rect 1717 -23554 1772 -11655
rect 1996 -12862 7070 -11824
rect 7814 -12034 21870 -11798
rect 13436 -12194 21870 -12034
rect 8348 -12382 9840 -12322
rect 13436 -12680 20150 -12510
rect 20656 -12646 21870 -12194
rect 7778 -12752 20150 -12680
rect 1996 -13538 2982 -12862
rect 7778 -12898 19808 -12752
rect 19070 -13098 19808 -12898
rect 20008 -13352 20788 -13244
rect 20918 -13350 21698 -13242
rect 1996 -13814 19328 -13538
rect 19998 -13600 20798 -13452
rect 20908 -13600 21708 -13452
rect 20010 -13870 20786 -13702
rect 20920 -13800 21696 -13700
rect 22152 -12538 25456 -11668
rect 20204 -14336 20622 -13870
rect 20920 -13952 21696 -13856
rect 21828 -13874 21944 -13758
rect 20916 -14308 21698 -14052
rect 20010 -14500 20786 -14336
rect 20920 -14504 21696 -14404
rect 19998 -14750 20798 -14602
rect 20908 -14748 21708 -14600
rect 20008 -14962 20788 -14854
rect 20920 -14962 21700 -14854
rect 19534 -15878 21862 -15548
rect 19534 -16020 20220 -15878
rect 19534 -17992 20222 -16020
rect 20474 -16268 21252 -16008
rect 21532 -16254 21862 -15878
rect 20476 -16424 21252 -16332
rect 20476 -16582 21252 -16490
rect 20476 -16740 21252 -16648
rect 20476 -16898 21252 -16806
rect 20476 -17056 21252 -16964
rect 20476 -17214 21252 -17122
rect 20476 -17372 21252 -17280
rect 20476 -17530 21252 -17438
rect 20476 -17688 21252 -17596
rect 19534 -18128 20220 -17992
rect 20472 -17996 21252 -17756
rect 20474 -18010 21252 -17996
rect 22608 -13138 23388 -13092
rect 22608 -13344 23390 -13138
rect 22608 -13392 23388 -13344
rect 23538 -13390 24318 -13090
rect 22610 -13968 23390 -13668
rect 23536 -13716 24316 -13666
rect 23536 -13922 24318 -13716
rect 23536 -13966 24316 -13922
rect 22608 -14298 23388 -14242
rect 22608 -14504 23390 -14298
rect 22608 -14542 23388 -14504
rect 23538 -14538 24318 -14238
rect 22610 -14976 23390 -14814
rect 22612 -15642 23390 -15598
rect 23570 -15622 24284 -14908
rect 22610 -15914 23392 -15642
rect 22610 -16288 23390 -15988
rect 23538 -16288 24318 -15988
rect 22610 -16852 23390 -16552
rect 23536 -16606 24316 -16552
rect 23536 -16812 24318 -16606
rect 23536 -16852 24316 -16812
rect 22610 -17438 23390 -17138
rect 23538 -17436 24318 -17136
rect 24616 -17924 25456 -12538
rect 1996 -18408 18346 -18128
rect 18856 -18408 20220 -18128
rect 19534 -18466 20220 -18408
rect 1890 -23440 20268 -22710
rect 21482 -23096 21544 -22828
rect 21226 -23158 21544 -23096
rect 1717 -23587 20600 -23554
rect 1674 -23613 20600 -23587
rect 21764 -23598 22366 -23090
rect 22604 -23098 22666 -22830
rect 25228 -22730 25456 -17924
rect 22604 -23160 22922 -23098
rect 24070 -23230 25456 -22730
rect 23578 -23613 25456 -23230
rect 1674 -23647 1743 -23613
rect 1743 -23647 20600 -23613
rect 23578 -23630 25453 -23613
rect 25453 -23630 25456 -23613
rect 1674 -23656 20600 -23647
<< metal1 >>
rect 1626 -826 2026 -812
rect 1626 -1200 1638 -826
rect 2012 -1200 2026 -826
rect 1626 -1212 2026 -1200
rect 2178 -826 2578 -812
rect 2178 -1200 2190 -826
rect 2564 -1200 2578 -826
rect 3592 -826 3992 -812
rect 2178 -1212 2578 -1200
rect 2676 -864 2820 -850
rect 2676 -1182 2748 -864
rect 2806 -1110 2820 -864
rect 3592 -946 3606 -826
rect 2882 -956 3606 -946
rect 2882 -1046 3156 -956
rect 2806 -1128 3046 -1110
rect 3018 -1182 3046 -1128
rect 2676 -1236 3046 -1182
rect 3146 -1180 3156 -1046
rect 3236 -1046 3606 -956
rect 3236 -1180 3246 -1046
rect 3146 -1194 3246 -1180
rect 3592 -1200 3606 -1046
rect 3980 -1200 3992 -826
rect 3592 -1212 3992 -1200
rect 4338 -824 4738 -812
rect 4338 -1198 4350 -824
rect 4724 -948 4738 -824
rect 8076 -822 8476 -812
rect 5516 -852 6032 -850
rect 5516 -854 6112 -852
rect 7030 -854 7966 -852
rect 5516 -884 7966 -854
rect 4724 -958 5454 -948
rect 4724 -1048 5096 -958
rect 4724 -1198 4738 -1048
rect 5086 -1180 5096 -1048
rect 5176 -1048 5454 -958
rect 5176 -1180 5186 -1048
rect 5516 -1110 5530 -884
rect 5086 -1192 5186 -1180
rect 5290 -1126 5530 -1110
rect 5586 -890 7966 -884
rect 5290 -1180 5316 -1126
rect 5586 -1180 6110 -890
rect 7000 -896 7966 -890
rect 4338 -1212 4738 -1198
rect 5290 -1236 6110 -1180
rect 2676 -1354 2946 -1236
rect 1752 -1378 2946 -1354
rect 1752 -3222 1782 -1378
rect 2162 -1600 2946 -1378
rect 2162 -1856 2756 -1600
rect 3038 -1690 3426 -1680
rect 3038 -1772 3046 -1690
rect 3414 -1772 3426 -1690
rect 3038 -1780 3426 -1772
rect 3038 -1842 3278 -1780
rect 2162 -2476 2428 -1856
rect 3518 -1864 4838 -1286
rect 5414 -1600 6110 -1236
rect 7934 -1272 7966 -896
rect 8076 -1200 8088 -822
rect 8464 -1200 8476 -822
rect 9976 -818 10376 -812
rect 9976 -846 9982 -818
rect 8076 -1212 8476 -1200
rect 8592 -882 9982 -846
rect 10370 -846 10376 -818
rect 11192 -822 11592 -812
rect 10370 -882 11094 -846
rect 4904 -1682 5292 -1672
rect 4904 -1764 4912 -1682
rect 5280 -1764 5292 -1682
rect 4904 -1772 5292 -1764
rect 5058 -1842 5292 -1772
rect 5578 -1846 6110 -1600
rect 3894 -1866 4838 -1864
rect 4060 -1886 4294 -1866
rect 4110 -2044 4228 -1886
rect 2162 -2854 3056 -2476
rect 3632 -2726 3788 -2488
rect 5702 -2482 6110 -1846
rect 4544 -2726 4692 -2488
rect 3632 -2770 4692 -2726
rect 5276 -2854 6110 -2482
rect 2162 -2870 6110 -2854
rect 2162 -2952 3880 -2870
rect 4452 -2952 6110 -2870
rect 7000 -1294 7966 -1272
rect 8592 -1262 8606 -882
rect 11080 -1262 11094 -882
rect 11192 -1204 11200 -822
rect 11580 -1204 11592 -822
rect 23912 -820 24312 -812
rect 22388 -842 23810 -840
rect 14212 -846 23810 -842
rect 11192 -1212 11592 -1204
rect 11644 -914 23810 -846
rect 8592 -1276 11094 -1262
rect 11644 -1262 11672 -914
rect 23756 -1138 23810 -914
rect 13494 -1242 22662 -1138
rect 11644 -1286 12602 -1262
rect 1752 -3248 3880 -3222
rect 2084 -3308 3880 -3248
rect 4452 -3308 6720 -3222
rect 2084 -3330 6720 -3308
rect 2300 -3594 6034 -3578
rect 1626 -3600 6034 -3594
rect 1626 -5026 1636 -3600
rect 1920 -3858 6034 -3600
rect 1920 -5026 2452 -3858
rect 1626 -5036 2452 -5026
rect 4108 -5044 4226 -3858
rect 1936 -5122 2328 -5102
rect 4098 -5116 4232 -5102
rect 1936 -5154 2048 -5122
rect 1936 -6772 1990 -5154
rect 2476 -6772 3952 -6542
rect 1936 -6798 2048 -6772
rect 2454 -6798 3952 -6772
rect 1936 -6808 3952 -6798
rect 5958 -5156 6416 -5104
rect 4374 -6774 5838 -6542
rect 6324 -6774 6416 -5156
rect 4374 -6808 6416 -6774
rect 1936 -6822 6416 -6808
rect 3364 -7116 3370 -6962
rect 2496 -7126 3370 -7116
rect 2496 -7214 2510 -7126
rect 3230 -7214 3370 -7126
rect 2496 -7222 3370 -7214
rect 3478 -7222 3484 -6962
rect 3614 -7214 3620 -6954
rect 3728 -7110 3734 -6954
rect 3728 -7120 4600 -7110
rect 3728 -7208 3888 -7120
rect 4588 -7208 4600 -7120
rect 3728 -7214 4600 -7208
rect 2406 -8054 2412 -7254
rect 2520 -8054 2526 -7254
rect 2564 -8054 2570 -7254
rect 2678 -8054 2684 -7254
rect 2722 -8054 2728 -7254
rect 2836 -8054 2842 -7254
rect 2880 -8054 2886 -7254
rect 2994 -8054 3000 -7254
rect 3036 -8054 3042 -7254
rect 3150 -8054 3156 -7254
rect 3196 -8054 3202 -7254
rect 3310 -8054 3316 -7254
rect 3364 -8078 3370 -7906
rect 3478 -8078 3484 -7906
rect 3364 -8086 3484 -8078
rect 2496 -8092 3484 -8086
rect 2496 -8172 2512 -8092
rect 3212 -8172 3484 -8092
rect 2496 -8184 3484 -8172
rect 3614 -8078 3620 -7916
rect 3728 -8078 3734 -7916
rect 3782 -8054 3790 -7254
rect 3894 -8054 3902 -7254
rect 3940 -8054 3946 -7254
rect 4054 -8054 4060 -7254
rect 4098 -8054 4104 -7254
rect 4212 -8054 4218 -7254
rect 4256 -8054 4262 -7254
rect 4370 -8054 4376 -7254
rect 4414 -8054 4420 -7254
rect 4528 -8054 4534 -7254
rect 4572 -8054 4578 -7254
rect 4686 -8054 4692 -7254
rect 3614 -8096 3734 -8078
rect 3614 -8102 4608 -8096
rect 3614 -8188 3888 -8102
rect 4594 -8188 4608 -8102
rect 3614 -8196 4608 -8188
rect 6654 -9258 6720 -3330
rect 7000 -3410 7048 -1294
rect 7372 -1344 7472 -1338
rect 7234 -1444 7372 -1344
rect 7472 -1444 12358 -1344
rect 12458 -1444 12464 -1344
rect 7235 -2028 7334 -1444
rect 7372 -1450 7472 -1444
rect 7378 -1500 7478 -1494
rect 7478 -1600 12184 -1500
rect 12284 -1600 12290 -1500
rect 12558 -1582 12602 -1286
rect 13494 -1484 13950 -1242
rect 14430 -1260 22662 -1242
rect 14434 -1282 22662 -1260
rect 13494 -1490 13562 -1484
rect 13370 -1582 13562 -1490
rect 7378 -1606 7478 -1600
rect 7378 -1684 7478 -1678
rect 7478 -1784 12006 -1684
rect 12106 -1784 12112 -1684
rect 12424 -1740 13562 -1582
rect 7378 -1790 7478 -1784
rect 7234 -2082 9044 -2028
rect 7234 -2128 7514 -2082
rect 9032 -2128 9044 -2082
rect 7234 -2136 9044 -2128
rect 9222 -2048 9322 -1784
rect 9222 -2092 10966 -2048
rect 7235 -2612 7334 -2136
rect 9222 -2140 9438 -2092
rect 10952 -2140 10966 -2092
rect 9222 -2148 10966 -2140
rect 7432 -2194 7552 -2188
rect 7235 -2685 7336 -2612
rect 7236 -3038 7336 -2685
rect 7432 -2982 7434 -2194
rect 7550 -2982 7552 -2194
rect 7432 -2988 7552 -2982
rect 7592 -2194 7712 -2188
rect 7592 -2982 7594 -2194
rect 7710 -2982 7712 -2194
rect 7592 -2988 7712 -2982
rect 7750 -2194 7870 -2188
rect 7750 -2982 7752 -2194
rect 7868 -2982 7870 -2194
rect 7750 -2988 7870 -2982
rect 7908 -2194 8028 -2188
rect 7908 -2982 7910 -2194
rect 8026 -2982 8028 -2194
rect 7908 -2988 8028 -2982
rect 8066 -2194 8186 -2188
rect 8066 -2982 8068 -2194
rect 8184 -2982 8186 -2194
rect 8066 -2988 8186 -2982
rect 8222 -2192 8342 -2186
rect 8222 -2980 8224 -2192
rect 8340 -2980 8342 -2192
rect 8222 -2986 8342 -2980
rect 8380 -2194 8500 -2188
rect 8380 -2982 8382 -2194
rect 8498 -2982 8500 -2194
rect 8380 -2988 8500 -2982
rect 8540 -2192 8660 -2186
rect 8540 -2980 8542 -2192
rect 8658 -2980 8660 -2192
rect 8540 -2986 8660 -2980
rect 8696 -2194 8816 -2188
rect 8696 -2982 8698 -2194
rect 8814 -2982 8816 -2194
rect 8696 -2988 8816 -2982
rect 8854 -2194 8974 -2188
rect 8854 -2982 8856 -2194
rect 8972 -2982 8974 -2194
rect 8854 -2988 8974 -2982
rect 9012 -2194 9132 -2188
rect 9012 -2982 9014 -2194
rect 9130 -2982 9132 -2194
rect 9012 -2988 9132 -2982
rect 9222 -3036 9322 -2148
rect 11300 -2176 11474 -2164
rect 9358 -2198 9478 -2192
rect 9358 -2986 9360 -2198
rect 9476 -2986 9478 -2198
rect 9358 -2992 9478 -2986
rect 9516 -2198 9636 -2192
rect 9516 -2986 9518 -2198
rect 9634 -2986 9636 -2198
rect 9516 -2992 9636 -2986
rect 9676 -2198 9796 -2192
rect 9676 -2986 9678 -2198
rect 9794 -2986 9796 -2198
rect 9676 -2992 9796 -2986
rect 9834 -2198 9954 -2192
rect 9834 -2986 9836 -2198
rect 9952 -2986 9954 -2198
rect 9834 -2992 9954 -2986
rect 9990 -2198 10110 -2192
rect 9990 -2986 9992 -2198
rect 10108 -2986 10110 -2198
rect 9990 -2992 10110 -2986
rect 10150 -2198 10270 -2192
rect 10150 -2986 10152 -2198
rect 10268 -2986 10270 -2198
rect 10150 -2992 10270 -2986
rect 10306 -2198 10426 -2192
rect 10306 -2986 10308 -2198
rect 10424 -2986 10426 -2198
rect 10306 -2992 10426 -2986
rect 10464 -2198 10584 -2192
rect 10464 -2986 10466 -2198
rect 10582 -2986 10584 -2198
rect 10464 -2992 10584 -2986
rect 10624 -2198 10744 -2192
rect 10624 -2986 10626 -2198
rect 10742 -2986 10744 -2198
rect 10624 -2992 10744 -2986
rect 10780 -2198 10900 -2192
rect 10780 -2986 10782 -2198
rect 10898 -2986 10900 -2198
rect 10780 -2992 10900 -2986
rect 10938 -2198 11058 -2192
rect 10938 -2986 10940 -2198
rect 11056 -2986 11058 -2198
rect 11300 -2964 11310 -2176
rect 11462 -2180 11474 -2176
rect 11468 -2958 11474 -2180
rect 11462 -2964 11474 -2958
rect 11300 -2974 11474 -2964
rect 10938 -2992 11058 -2986
rect 11504 -3012 11550 -2082
rect 12204 -2154 13562 -1740
rect 12204 -2156 13048 -2154
rect 11592 -2182 11980 -2170
rect 11592 -2956 11606 -2182
rect 11666 -2956 11980 -2182
rect 11592 -2968 11980 -2956
rect 11772 -2980 11980 -2968
rect 7236 -3046 9046 -3038
rect 7236 -3092 7512 -3046
rect 9034 -3092 9046 -3046
rect 7236 -3138 9046 -3092
rect 9222 -3044 10966 -3036
rect 9222 -3092 9436 -3044
rect 10952 -3092 10966 -3044
rect 9222 -3136 10966 -3092
rect 11480 -3198 11580 -3012
rect 11772 -3164 11780 -2980
rect 11972 -3164 11980 -2980
rect 11772 -3172 11980 -3164
rect 12204 -2224 12634 -2156
rect 12770 -2224 12878 -2156
rect 13014 -2224 13048 -2156
rect 11416 -3208 11616 -3198
rect 11416 -3386 11426 -3208
rect 11604 -3386 11616 -3208
rect 11416 -3398 11616 -3386
rect 12204 -3216 12616 -2224
rect 13700 -2300 13800 -1724
rect 14866 -1750 22662 -1282
rect 12702 -2400 13800 -2300
rect 13028 -2468 13960 -2446
rect 13028 -3026 13052 -2468
rect 13648 -3026 13960 -2468
rect 22388 -2834 22662 -1750
rect 13028 -3044 13960 -3026
rect 16104 -3004 22662 -2834
rect 12204 -3380 12462 -3216
rect 7000 -3412 7506 -3410
rect 7000 -3434 11330 -3412
rect 11294 -3444 11330 -3434
rect 12204 -3444 12222 -3380
rect 12588 -3390 12616 -3216
rect 12772 -3176 12874 -3062
rect 12772 -3294 13942 -3176
rect 12588 -3414 13840 -3390
rect 11294 -3470 12222 -3444
rect 13744 -3658 13840 -3414
rect 16104 -3422 16120 -3004
rect 16212 -3136 22662 -3004
rect 15008 -3442 16120 -3422
rect 15008 -3516 15034 -3442
rect 17524 -3490 22662 -3136
rect 23754 -3490 23810 -1138
rect 23912 -1200 23924 -820
rect 24302 -1200 24312 -820
rect 23912 -1212 24312 -1200
rect 24418 -898 25270 -834
rect 17524 -3514 22968 -3490
rect 16212 -3516 22968 -3514
rect 15008 -3534 22968 -3516
rect 8452 -3978 12318 -3948
rect 8452 -5446 8542 -3978
rect 12260 -4018 12318 -3978
rect 12260 -4020 13740 -4018
rect 13814 -4020 13840 -3658
rect 9140 -4152 9146 -4052
rect 9246 -4152 11462 -4052
rect 11562 -4152 11568 -4052
rect 12260 -4066 13840 -4020
rect 22916 -3976 22968 -3534
rect 23752 -3976 23810 -3490
rect 22916 -4026 23810 -3976
rect 24418 -3984 24460 -898
rect 25194 -3984 25270 -898
rect 24418 -4022 25270 -3984
rect 7418 -5528 8542 -5446
rect 8880 -4310 25158 -4298
rect 8880 -4316 12112 -4310
rect 15250 -4316 25158 -4310
rect 8880 -5476 8900 -4316
rect 11694 -4574 12058 -4548
rect 11694 -4734 11724 -4574
rect 10476 -4768 11724 -4734
rect 11772 -4626 11980 -4616
rect 10476 -4958 10494 -4768
rect 11772 -4810 11780 -4626
rect 11972 -4810 11980 -4626
rect 12034 -4750 12058 -4574
rect 16094 -4556 16958 -4548
rect 17330 -4556 18192 -4548
rect 16094 -4574 18192 -4556
rect 12034 -4760 12112 -4750
rect 15250 -4760 15282 -4750
rect 12034 -4768 15282 -4760
rect 11772 -4816 11980 -4810
rect 10662 -4896 15100 -4816
rect 11436 -4958 12014 -4896
rect 12592 -4958 12844 -4896
rect 13748 -4958 14326 -4896
rect 15264 -4958 15282 -4768
rect 10476 -4970 11230 -4958
rect 11224 -5346 11230 -4970
rect 10462 -5358 11230 -5346
rect 11436 -5354 11452 -4958
rect 11992 -5354 12014 -4958
rect 10462 -5476 10494 -5358
rect 11436 -5420 12014 -5354
rect 12104 -4970 12504 -4958
rect 12104 -5346 12122 -4970
rect 12488 -5346 12504 -4970
rect 12104 -5358 12504 -5346
rect 12592 -5358 12604 -4958
rect 12826 -5358 12844 -4958
rect 12918 -4970 13178 -4958
rect 12918 -5346 12924 -4970
rect 13168 -5346 13178 -4970
rect 12918 -5358 13178 -5346
rect 13260 -4970 13660 -4958
rect 13260 -5346 13276 -4970
rect 13642 -5346 13660 -4970
rect 13260 -5358 13660 -5346
rect 13748 -5354 13768 -4958
rect 14308 -5354 14326 -4958
rect 12592 -5420 12844 -5358
rect 13748 -5420 14326 -5354
rect 14532 -4970 15282 -4958
rect 14532 -5346 14538 -4970
rect 14532 -5358 15282 -5346
rect 8880 -5494 10494 -5476
rect 10662 -5500 15100 -5420
rect 7418 -7534 7506 -5528
rect 15264 -5530 15282 -5358
rect 16094 -5530 16118 -4574
rect 16260 -4700 17076 -4640
rect 16648 -4744 16924 -4700
rect 17106 -4734 17186 -4574
rect 17218 -4700 18034 -4640
rect 17266 -4706 17486 -4700
rect 16648 -4776 16666 -4744
rect 16210 -4794 16666 -4776
rect 16210 -5484 16228 -4794
rect 16210 -5502 16666 -5484
rect 15264 -5548 16118 -5530
rect 16648 -5530 16666 -5502
rect 16878 -5530 16924 -4744
rect 16648 -5576 16924 -5530
rect 17026 -4750 17266 -4734
rect 17026 -5526 17044 -4750
rect 17246 -5526 17266 -4750
rect 17026 -5542 17266 -5526
rect 17328 -5570 17424 -4706
rect 17498 -4742 18082 -4734
rect 17498 -5530 17508 -4742
rect 17702 -4750 18082 -4742
rect 18064 -5526 18082 -4750
rect 18002 -5530 18082 -5526
rect 17498 -5542 18082 -5530
rect 17266 -5576 17486 -5570
rect 7588 -7438 7604 -5608
rect 8962 -5636 16060 -5608
rect 8962 -5640 15260 -5636
rect 15938 -5752 16060 -5636
rect 16648 -5636 17534 -5576
rect 15938 -5758 16614 -5752
rect 10492 -5814 15260 -5776
rect 10492 -5988 10580 -5814
rect 10682 -5948 15086 -5888
rect 10492 -6000 11248 -5988
rect 11242 -6378 11248 -6000
rect 10492 -6388 11248 -6378
rect 10492 -6390 10680 -6388
rect 10492 -6516 10580 -6390
rect 10492 -6518 10680 -6516
rect 11088 -6518 11248 -6388
rect 10492 -6528 11248 -6518
rect 11242 -6906 11248 -6528
rect 10492 -6918 11248 -6906
rect 10492 -7086 10580 -6918
rect 11088 -7056 11248 -6918
rect 11362 -6958 11542 -5948
rect 11588 -5990 11892 -5984
rect 11588 -6000 11666 -5990
rect 11814 -6000 11892 -5990
rect 11588 -6378 11602 -6000
rect 11878 -6378 11892 -6000
rect 11588 -6388 11666 -6378
rect 11814 -6388 11892 -6378
rect 11588 -6394 11892 -6388
rect 11660 -6512 11820 -6394
rect 11586 -6518 11890 -6512
rect 11586 -6528 11666 -6518
rect 11814 -6528 11890 -6518
rect 11586 -6906 11602 -6528
rect 11878 -6906 11890 -6528
rect 11586 -6916 11666 -6906
rect 11814 -6916 11890 -6906
rect 11586 -6922 11890 -6916
rect 11936 -6958 12116 -5948
rect 12912 -5982 13260 -5948
rect 12164 -5988 12468 -5984
rect 12164 -6000 12850 -5988
rect 12164 -6378 12176 -6000
rect 12452 -6378 12850 -6000
rect 12164 -6394 12850 -6378
rect 12234 -6512 12394 -6394
rect 12912 -6430 12924 -5982
rect 13252 -6392 13260 -5982
rect 12440 -6468 12924 -6430
rect 13250 -6468 13260 -6392
rect 13300 -6000 13604 -5984
rect 13300 -6378 13316 -6000
rect 13592 -6378 13604 -6000
rect 13300 -6394 13604 -6378
rect 12440 -6476 13260 -6468
rect 12160 -6528 12464 -6512
rect 12160 -6530 12238 -6528
rect 12388 -6530 12464 -6528
rect 12160 -6908 12174 -6530
rect 12450 -6908 12464 -6530
rect 12160 -6922 12464 -6908
rect 11294 -7018 12184 -6958
rect 12234 -7056 12394 -6922
rect 12508 -6958 12688 -6476
rect 12730 -6518 13034 -6512
rect 12730 -6528 12810 -6518
rect 12958 -6528 13034 -6518
rect 12730 -6906 12742 -6528
rect 13018 -6906 13034 -6528
rect 12730 -6916 12810 -6906
rect 12958 -6916 13034 -6906
rect 12730 -6922 13034 -6916
rect 13080 -6958 13260 -6476
rect 13376 -6512 13536 -6394
rect 13304 -6528 13608 -6512
rect 13304 -6906 13316 -6528
rect 13592 -6906 13608 -6528
rect 13304 -6922 13608 -6906
rect 12440 -7018 13330 -6958
rect 13376 -7056 13536 -6922
rect 13650 -6958 13830 -5948
rect 13874 -5990 14178 -5984
rect 13874 -6000 13954 -5990
rect 14102 -6000 14178 -5990
rect 13874 -6378 13886 -6000
rect 14162 -6378 14178 -6000
rect 13874 -6388 13954 -6378
rect 14102 -6388 14178 -6378
rect 13874 -6394 14178 -6388
rect 13948 -6512 14108 -6394
rect 13876 -6518 14180 -6512
rect 13876 -6528 13954 -6518
rect 14102 -6528 14180 -6518
rect 13876 -6906 13888 -6528
rect 14164 -6906 14180 -6528
rect 13876 -6916 13954 -6906
rect 14102 -6916 14180 -6906
rect 13876 -6922 14180 -6916
rect 14222 -6958 14402 -5948
rect 15228 -5988 15260 -5814
rect 16602 -5888 16614 -5758
rect 14520 -6000 15260 -5988
rect 15938 -5894 16614 -5888
rect 14520 -6378 14526 -6000
rect 14520 -6388 15260 -6378
rect 14520 -6518 14680 -6388
rect 15228 -6518 15260 -6388
rect 14520 -6528 15260 -6518
rect 14520 -6906 14526 -6528
rect 14520 -6918 15260 -6906
rect 13584 -7018 14474 -6958
rect 14520 -7056 14680 -6918
rect 11088 -7086 14680 -7056
rect 15228 -7086 15260 -6918
rect 10492 -7114 15260 -7086
rect 15938 -7086 15964 -5894
rect 16036 -5960 16620 -5950
rect 16036 -6050 16162 -5960
rect 16608 -6050 16620 -5960
rect 16036 -6056 16620 -6050
rect 16036 -6554 16156 -6056
rect 16648 -6092 16728 -5636
rect 16762 -5762 17524 -5752
rect 16762 -5888 16776 -5762
rect 17510 -5888 17524 -5762
rect 16762 -5894 17524 -5888
rect 16758 -5956 17078 -5950
rect 16758 -6050 16770 -5956
rect 17066 -6050 17078 -5956
rect 16758 -6056 17078 -6050
rect 17216 -5956 17536 -5950
rect 17216 -6050 17228 -5956
rect 17524 -6050 17536 -5956
rect 17216 -6056 17536 -6050
rect 16036 -7036 16044 -6554
rect 16148 -6938 16156 -6554
rect 16208 -6108 16770 -6092
rect 16208 -6886 16224 -6108
rect 16758 -6886 16770 -6108
rect 16208 -6902 16770 -6886
rect 16830 -6938 16954 -6056
rect 16998 -6106 17298 -6092
rect 16998 -6890 17014 -6106
rect 17280 -6890 17298 -6106
rect 16998 -6902 17298 -6890
rect 17340 -6938 17464 -6056
rect 17564 -6092 17644 -5542
rect 18174 -5674 18192 -4574
rect 21246 -5244 22086 -5218
rect 21246 -5274 21272 -5244
rect 18848 -5382 20732 -5352
rect 18848 -5530 18878 -5382
rect 18848 -5548 18900 -5530
rect 18174 -5694 18808 -5674
rect 17684 -5762 18742 -5752
rect 17684 -5886 17700 -5762
rect 18728 -5850 18742 -5762
rect 18788 -5790 18808 -5694
rect 18862 -5790 18900 -5548
rect 19036 -5696 19090 -5478
rect 19230 -5696 20470 -5478
rect 18788 -5808 18900 -5790
rect 18728 -5864 20528 -5850
rect 17684 -5894 18330 -5886
rect 17674 -5960 18258 -5950
rect 17674 -6050 17686 -5960
rect 18132 -6050 18258 -5960
rect 17674 -6056 18258 -6050
rect 17520 -6100 18082 -6092
rect 17520 -6894 17528 -6100
rect 17782 -6108 18082 -6100
rect 18066 -6886 18082 -6108
rect 17782 -6894 18082 -6886
rect 17520 -6902 18082 -6894
rect 18138 -6554 18258 -6056
rect 18138 -6938 18146 -6554
rect 16148 -6944 17118 -6938
rect 16148 -7034 16162 -6944
rect 17078 -7034 17118 -6944
rect 16148 -7036 17118 -7034
rect 16036 -7044 17118 -7036
rect 16160 -7046 17118 -7044
rect 17176 -6944 18146 -6938
rect 17176 -7034 17216 -6944
rect 18132 -7034 18146 -6944
rect 17176 -7036 18146 -7034
rect 18250 -7036 18258 -6554
rect 17176 -7046 18258 -7036
rect 18304 -7086 18330 -5894
rect 20504 -6354 20528 -5864
rect 18834 -6382 20528 -6354
rect 20574 -6016 20674 -5530
rect 20714 -5776 20732 -5382
rect 21246 -5402 21270 -5274
rect 21462 -5334 21562 -5328
rect 21246 -5486 21400 -5402
rect 21214 -5508 21400 -5486
rect 21214 -5776 21232 -5508
rect 20714 -5790 21232 -5776
rect 20574 -6104 20580 -6016
rect 20668 -6104 20674 -6016
rect 18834 -6816 18898 -6382
rect 19036 -6702 19092 -6484
rect 19232 -6702 20460 -6484
rect 20574 -6654 20674 -6104
rect 20712 -5870 21212 -5850
rect 20712 -6816 20736 -5870
rect 21184 -6560 21212 -5870
rect 21290 -6010 21390 -5610
rect 21462 -5788 21468 -5334
rect 21556 -5788 21562 -5334
rect 21620 -5716 21662 -5244
rect 21462 -5794 21562 -5788
rect 21718 -6010 21818 -5328
rect 21290 -6110 21818 -6010
rect 21290 -6516 21390 -6110
rect 21464 -6330 21564 -6324
rect 21184 -6580 21272 -6560
rect 18834 -6844 20736 -6816
rect 21202 -6636 21272 -6580
rect 21202 -6742 21400 -6636
rect 21202 -6878 21272 -6742
rect 21464 -6820 21470 -6330
rect 21560 -6820 21564 -6330
rect 21464 -6826 21564 -6820
rect 21202 -6902 21274 -6878
rect 21620 -6902 21662 -6412
rect 21718 -6828 21818 -6110
rect 21900 -5990 22000 -5406
rect 22066 -5852 22086 -5244
rect 23274 -5322 23778 -5298
rect 23274 -5406 23294 -5322
rect 23376 -5404 23642 -5322
rect 23724 -5404 23778 -5322
rect 22816 -5422 23294 -5406
rect 22816 -5758 22836 -5422
rect 22638 -5776 22836 -5758
rect 22914 -5594 23666 -5494
rect 22638 -5852 22654 -5776
rect 22914 -5842 23014 -5594
rect 22066 -5872 22654 -5852
rect 22714 -5852 23014 -5842
rect 22374 -5948 22652 -5924
rect 21900 -5996 22308 -5990
rect 21900 -6124 22006 -5996
rect 22302 -6124 22308 -5996
rect 21900 -6130 22308 -6124
rect 21900 -6738 22000 -6130
rect 22374 -6188 22398 -5948
rect 22070 -6224 22398 -6188
rect 22070 -6902 22118 -6224
rect 22620 -6674 22652 -5948
rect 22714 -6132 22726 -5852
rect 23002 -6132 23014 -5852
rect 22714 -6142 23014 -6132
rect 23434 -5930 23584 -5654
rect 23756 -5834 23778 -5404
rect 25134 -5834 25158 -4316
rect 23756 -5858 25158 -5834
rect 24010 -5930 24210 -5924
rect 23434 -6130 24010 -5930
rect 22714 -6496 22814 -6142
rect 23434 -6438 23584 -6130
rect 24010 -6136 24210 -6130
rect 24286 -5946 25202 -5924
rect 24286 -6220 24312 -5946
rect 24082 -6246 24312 -6220
rect 22714 -6596 24016 -6496
rect 24082 -6674 24114 -6246
rect 22620 -6694 22982 -6674
rect 22930 -6776 22982 -6694
rect 23332 -6774 23730 -6674
rect 24080 -6774 24114 -6674
rect 23332 -6776 24114 -6774
rect 22930 -6802 24114 -6776
rect 25178 -6674 25202 -5946
rect 25178 -6802 25204 -6674
rect 21202 -6930 22118 -6902
rect 15938 -7114 18330 -7086
rect 25180 -7248 25204 -6802
rect 21202 -7250 25204 -7248
rect 10008 -7290 25204 -7250
rect 10008 -7366 10100 -7290
rect 8962 -7410 10100 -7366
rect 8962 -7438 9648 -7410
rect 7588 -7454 9648 -7438
rect 9792 -7454 9902 -7410
rect 10046 -7454 10100 -7410
rect 24218 -7402 24654 -7390
rect 9792 -7474 9798 -7454
rect 9896 -7474 9902 -7454
rect 7418 -7614 8512 -7534
rect 9736 -7570 9952 -7548
rect 1858 -9330 6720 -9258
rect 8426 -9258 8512 -7614
rect 8920 -7608 9068 -7586
rect 8426 -9330 8516 -9258
rect 1858 -11096 1910 -9330
rect 8428 -10482 8516 -9330
rect 8920 -10142 8940 -7608
rect 9046 -9422 9068 -7608
rect 9148 -7774 9364 -7684
rect 9148 -9240 9208 -7774
rect 9304 -8908 9364 -7774
rect 9736 -8908 9788 -7570
rect 9304 -9002 9788 -8908
rect 9304 -9240 9364 -9002
rect 9736 -9050 9788 -9002
rect 9904 -8908 9952 -7570
rect 10618 -7674 11048 -7438
rect 24218 -7540 24230 -7402
rect 24644 -7540 24654 -7402
rect 24218 -7550 24654 -7540
rect 24760 -7404 25152 -7368
rect 10620 -8006 11050 -7770
rect 24220 -7840 24650 -7604
rect 10620 -8338 11050 -8102
rect 24220 -8172 24650 -7936
rect 10620 -8670 11050 -8434
rect 24220 -8502 24650 -8266
rect 9904 -9002 10547 -8908
rect 10620 -9002 11050 -8766
rect 24220 -8834 24650 -8598
rect 9904 -9050 9952 -9002
rect 9736 -9132 9952 -9050
rect 10146 -9088 10384 -9066
rect 9148 -9268 9364 -9240
rect 10146 -9386 10162 -9088
rect 9208 -9422 9308 -9386
rect 9448 -9406 10162 -9386
rect 9448 -9408 9636 -9406
rect 10048 -9408 10162 -9406
rect 9448 -9422 9466 -9408
rect 9046 -9442 9466 -9422
rect 10362 -9940 10384 -9088
rect 10453 -9751 10547 -9002
rect 10620 -9334 11050 -9098
rect 24220 -9166 24650 -8930
rect 10620 -9664 11050 -9428
rect 24220 -9500 24650 -9264
rect 10453 -9845 11069 -9751
rect 24220 -9832 24650 -9596
rect 24760 -9940 24788 -7404
rect 10362 -9960 24788 -9940
rect 25116 -10142 25152 -7404
rect 8920 -10144 24792 -10142
rect 25112 -10144 25152 -10142
rect 8920 -10176 25152 -10144
rect 15968 -10464 25450 -10450
rect 8428 -10544 15856 -10482
rect 15780 -11092 15856 -10544
rect 8428 -11096 15856 -11092
rect 1858 -11146 15856 -11096
rect 15968 -11130 15988 -10464
rect 16648 -10898 17142 -10464
rect 18052 -10898 25450 -10464
rect 16648 -11130 25450 -10898
rect 1858 -11148 8516 -11146
rect 15968 -11150 25450 -11130
rect 1844 -11310 21916 -11292
rect 1844 -11314 17714 -11310
rect 1662 -11588 1786 -11576
rect 1662 -23656 1674 -11588
rect 1772 -23544 1786 -11588
rect 1844 -11824 2030 -11314
rect 3298 -11484 17714 -11314
rect 3298 -11798 15036 -11484
rect 15812 -11798 17714 -11484
rect 18284 -11798 21916 -11310
rect 3298 -11824 7814 -11798
rect 1844 -13814 1996 -11824
rect 7070 -12022 7814 -11824
rect 7070 -12862 7118 -12022
rect 7752 -12034 7814 -12022
rect 7752 -12082 13436 -12034
rect 13404 -12194 13436 -12082
rect 7370 -12501 7478 -12200
rect 13404 -12226 20656 -12194
rect 7534 -12270 7714 -12260
rect 7534 -12430 7542 -12270
rect 7704 -12430 7714 -12270
rect 7534 -12440 7714 -12430
rect 8336 -12264 9798 -12262
rect 8336 -12322 9886 -12264
rect 8336 -12382 8348 -12322
rect 9840 -12382 9886 -12322
rect 8336 -12442 9886 -12382
rect 9978 -12268 11464 -12252
rect 9978 -12434 9998 -12268
rect 11440 -12434 11464 -12268
rect 9978 -12452 11464 -12434
rect 11640 -12268 13126 -12252
rect 11640 -12434 11662 -12268
rect 13104 -12434 13126 -12268
rect 20278 -12298 20478 -12284
rect 20278 -12302 20292 -12298
rect 13236 -12306 20292 -12302
rect 13190 -12398 20292 -12306
rect 13236 -12402 20292 -12398
rect 11640 -12452 13126 -12434
rect 20278 -12468 20292 -12402
rect 20464 -12468 20478 -12298
rect 2982 -12958 7118 -12862
rect 7339 -12620 7514 -12501
rect 13404 -12510 20194 -12474
rect 20278 -12484 20478 -12468
rect 13404 -12618 13436 -12510
rect 7339 -12910 7346 -12620
rect 7506 -12910 7514 -12620
rect 7339 -12916 7514 -12910
rect 7744 -12680 13436 -12618
rect 20150 -12618 20194 -12510
rect 20610 -12618 20656 -12226
rect 20150 -12646 20656 -12618
rect 21870 -12646 21916 -11798
rect 22120 -11596 25450 -11150
rect 22120 -11668 25512 -11596
rect 22120 -12538 22152 -11668
rect 22120 -12574 24616 -12538
rect 7744 -12898 7778 -12680
rect 20150 -12752 21916 -12646
rect 7744 -12954 19070 -12898
rect 2982 -13448 3002 -12958
rect 3134 -13314 3566 -13098
rect 4022 -13448 4422 -12958
rect 6016 -13448 6416 -12958
rect 8000 -13448 8400 -12954
rect 10006 -13448 10406 -12954
rect 12016 -13448 12416 -12954
rect 14008 -13448 14408 -12954
rect 16002 -13448 16402 -12954
rect 18008 -13098 19070 -12954
rect 19808 -13098 21916 -12752
rect 18008 -13112 21916 -13098
rect 22452 -12834 22556 -12794
rect 23444 -12834 23486 -12794
rect 22452 -12836 23486 -12834
rect 24374 -12796 24416 -12794
rect 24374 -12836 24376 -12796
rect 22452 -13028 24376 -12836
rect 18008 -13448 18408 -13112
rect 18532 -13242 21712 -13228
rect 18532 -13244 20918 -13242
rect 18532 -13322 20008 -13244
rect 18532 -13350 19822 -13322
rect 19460 -13368 19822 -13350
rect 19994 -13352 20008 -13322
rect 20788 -13330 20918 -13244
rect 20788 -13352 20802 -13330
rect 19994 -13368 20802 -13352
rect 20904 -13350 20918 -13330
rect 21698 -13350 21712 -13242
rect 20904 -13368 21712 -13350
rect 2982 -13538 19350 -13448
rect 19328 -13814 19350 -13538
rect 1844 -13888 19350 -13814
rect 1844 -13892 4972 -13888
rect 5450 -13890 19350 -13888
rect 5450 -13892 8958 -13890
rect 9436 -13892 19350 -13890
rect 1844 -18044 1970 -13892
rect 2132 -14254 2564 -14038
rect 2134 -14584 2566 -14368
rect 2132 -14916 2564 -14700
rect 2132 -15248 2564 -15032
rect 2130 -15578 2562 -15362
rect 2132 -15912 2564 -15696
rect 2132 -16242 2564 -16026
rect 2132 -16576 2564 -16360
rect 2130 -16908 2562 -16692
rect 2130 -17240 2562 -17024
rect 2132 -17570 2564 -17354
rect 2132 -17904 2564 -17688
rect 5008 -18044 5408 -18040
rect 7024 -18044 7424 -13892
rect 9006 -18044 9406 -18042
rect 11014 -18044 11414 -13892
rect 14994 -18044 15394 -13892
rect 16042 -13978 16556 -13972
rect 16042 -13980 19366 -13978
rect 16042 -14472 16050 -13980
rect 16548 -13994 19366 -13980
rect 16548 -14456 18384 -13994
rect 19346 -14132 19366 -13994
rect 18848 -14146 19366 -14132
rect 18848 -14456 18870 -14146
rect 18932 -14418 19364 -14202
rect 16548 -14466 18870 -14456
rect 16548 -14472 16556 -14466
rect 16042 -14480 16556 -14472
rect 18932 -14750 19364 -14534
rect 19460 -14838 19640 -13368
rect 19698 -13440 21780 -13426
rect 19698 -14762 19712 -13440
rect 19844 -13452 21780 -13440
rect 19844 -13600 19998 -13452
rect 20798 -13600 20908 -13452
rect 21708 -13600 21780 -13452
rect 19844 -13626 21780 -13600
rect 22452 -13450 22554 -13028
rect 23442 -13070 23488 -13028
rect 22596 -13092 23404 -13078
rect 22596 -13392 22608 -13092
rect 23388 -13138 23404 -13092
rect 23390 -13160 23404 -13138
rect 23524 -13090 24332 -13078
rect 23524 -13160 23538 -13090
rect 23390 -13326 23538 -13160
rect 23390 -13344 23404 -13326
rect 23388 -13392 23404 -13344
rect 22596 -13402 23404 -13392
rect 23524 -13390 23538 -13326
rect 24318 -13160 24332 -13090
rect 24548 -13160 24616 -12574
rect 24318 -13326 24616 -13160
rect 24318 -13390 24332 -13326
rect 23524 -13402 24332 -13390
rect 24376 -13450 24478 -13374
rect 22452 -13618 24478 -13450
rect 19844 -14576 19858 -13626
rect 19994 -13702 20802 -13680
rect 19994 -13870 20010 -13702
rect 19994 -13896 20204 -13870
rect 20174 -14308 20204 -13896
rect 19994 -14336 20204 -14308
rect 19994 -14500 20010 -14336
rect 20786 -13718 20802 -13702
rect 20904 -13700 21712 -13680
rect 20904 -13718 20920 -13700
rect 20786 -13800 20920 -13718
rect 21696 -13800 21712 -13700
rect 21816 -13758 21956 -13746
rect 20786 -13820 21712 -13800
rect 20786 -13870 20802 -13820
rect 21748 -13848 21828 -13758
rect 20622 -13896 20802 -13870
rect 20908 -13856 21828 -13848
rect 20622 -14308 20654 -13896
rect 20908 -13952 20920 -13856
rect 21696 -13874 21828 -13856
rect 21944 -13874 21956 -13758
rect 21696 -13908 21956 -13874
rect 21696 -13952 21708 -13908
rect 20908 -13964 21708 -13952
rect 20854 -14030 21764 -14008
rect 20854 -14306 20882 -14030
rect 21736 -14170 21764 -14030
rect 22452 -14022 22554 -13618
rect 22594 -13668 23402 -13656
rect 22594 -13968 22610 -13668
rect 23390 -13702 23402 -13668
rect 23520 -13666 24328 -13656
rect 23390 -13738 23404 -13702
rect 23520 -13738 23536 -13666
rect 24316 -13702 24328 -13666
rect 24316 -13714 24330 -13702
rect 23390 -13904 23536 -13738
rect 23390 -13942 23404 -13904
rect 23390 -13968 23402 -13942
rect 22594 -13980 23402 -13968
rect 23520 -13966 23536 -13904
rect 24318 -13922 24330 -13714
rect 24316 -13942 24330 -13922
rect 24316 -13966 24328 -13942
rect 23520 -13980 24328 -13966
rect 24376 -14022 24478 -13618
rect 21736 -14306 22400 -14170
rect 20854 -14308 20916 -14306
rect 21698 -14308 22400 -14306
rect 20622 -14336 20802 -14308
rect 20854 -14330 22400 -14308
rect 20786 -14384 20802 -14336
rect 20786 -14404 22156 -14384
rect 20786 -14486 20920 -14404
rect 20786 -14500 20802 -14486
rect 19994 -14524 20802 -14500
rect 20904 -14504 20920 -14486
rect 21696 -14482 22156 -14404
rect 21696 -14504 21712 -14482
rect 20904 -14524 21712 -14504
rect 19844 -14600 21782 -14576
rect 19844 -14602 20908 -14600
rect 19844 -14750 19998 -14602
rect 20798 -14748 20908 -14602
rect 21708 -14748 21782 -14600
rect 20798 -14750 21782 -14748
rect 19844 -14762 21782 -14750
rect 19698 -14776 21782 -14762
rect 18932 -15082 19364 -14866
rect 19460 -14884 19822 -14838
rect 19994 -14854 20802 -14838
rect 19994 -14884 20008 -14854
rect 19460 -14962 20008 -14884
rect 20788 -14876 20802 -14854
rect 20904 -14854 21712 -14838
rect 20904 -14876 20920 -14854
rect 20788 -14962 20920 -14876
rect 21700 -14962 21712 -14854
rect 19460 -14978 21712 -14962
rect 18402 -15164 18802 -15148
rect 18402 -15530 18420 -15164
rect 18784 -15530 18802 -15164
rect 18932 -15414 19364 -15198
rect 18402 -15548 18802 -15530
rect 18426 -17798 18776 -15548
rect 18932 -15746 19364 -15530
rect 19502 -15548 21878 -15122
rect 18932 -16078 19364 -15862
rect 18932 -16410 19364 -16194
rect 18932 -16742 19364 -16526
rect 18932 -17074 19364 -16858
rect 18932 -17406 19364 -17190
rect 18932 -17738 19364 -17522
rect 18426 -17958 19376 -17798
rect 1844 -18128 18352 -18044
rect 1844 -18408 1996 -18128
rect 18346 -18408 18352 -18128
rect 1844 -18484 18352 -18408
rect 1844 -18486 4962 -18484
rect 5456 -18486 18352 -18484
rect 1844 -22670 1970 -18486
rect 2130 -18850 2564 -18616
rect 2130 -19184 2564 -18950
rect 2130 -19514 2564 -19280
rect 2130 -19846 2564 -19612
rect 2130 -20180 2564 -19946
rect 2130 -20510 2564 -20276
rect 2130 -20842 2564 -20608
rect 2128 -21174 2562 -20940
rect 2130 -21506 2564 -21272
rect 2130 -21838 2564 -21604
rect 2128 -22170 2562 -21936
rect 2136 -22232 2670 -22222
rect 2136 -22372 2148 -22232
rect 2654 -22372 2670 -22232
rect 2136 -22382 2670 -22372
rect 5008 -22670 5408 -22668
rect 9006 -22670 9406 -18486
rect 13040 -22670 13440 -18486
rect 16960 -22670 17360 -18486
rect 18426 -18578 18776 -17958
rect 19502 -18044 19534 -15548
rect 20220 -15918 21532 -15878
rect 20220 -15994 20252 -15918
rect 20220 -16020 20254 -15994
rect 20222 -17992 20254 -16020
rect 20464 -16008 21264 -15994
rect 18850 -18128 19534 -18044
rect 20220 -18022 20254 -17992
rect 18850 -18408 18856 -18128
rect 18850 -18466 19534 -18408
rect 20220 -18466 20252 -18022
rect 20332 -18116 20432 -16094
rect 20464 -16268 20474 -16008
rect 21252 -16268 21264 -16008
rect 20464 -16284 21264 -16268
rect 20464 -16324 21264 -16312
rect 20464 -16430 20474 -16324
rect 21252 -16430 21264 -16324
rect 20464 -16442 21264 -16430
rect 20464 -16482 21264 -16470
rect 20464 -16588 20474 -16482
rect 21252 -16588 21264 -16482
rect 20464 -16600 21264 -16588
rect 20464 -16640 21264 -16628
rect 20464 -16746 20474 -16640
rect 21252 -16746 21264 -16640
rect 20464 -16758 21264 -16746
rect 20464 -16798 21264 -16786
rect 20464 -16904 20474 -16798
rect 21252 -16904 21264 -16798
rect 20464 -16916 21264 -16904
rect 20464 -16956 21264 -16944
rect 20464 -17062 20474 -16956
rect 21252 -17062 21264 -16956
rect 20464 -17074 21264 -17062
rect 20464 -17114 21264 -17102
rect 20464 -17220 20476 -17114
rect 21254 -17220 21264 -17114
rect 20464 -17232 21264 -17220
rect 20464 -17272 21264 -17260
rect 20464 -17378 20474 -17272
rect 21252 -17378 21264 -17272
rect 20464 -17390 21264 -17378
rect 20464 -17430 21264 -17418
rect 20464 -17536 20474 -17430
rect 21252 -17536 21264 -17430
rect 20464 -17548 21264 -17536
rect 20464 -17588 21264 -17576
rect 20464 -17694 20474 -17588
rect 21252 -17694 21264 -17588
rect 20464 -17706 21264 -17694
rect 20464 -17750 21264 -17734
rect 20464 -17756 20476 -17750
rect 21250 -17756 21264 -17750
rect 20464 -17996 20472 -17756
rect 20464 -18010 20474 -17996
rect 21252 -18010 21264 -17756
rect 20464 -18022 21264 -18010
rect 21296 -18116 21396 -16094
rect 21520 -16254 21532 -15918
rect 21862 -16254 21878 -15548
rect 21956 -15590 22156 -14482
rect 22240 -14884 22400 -14330
rect 22452 -14190 24478 -14022
rect 22452 -14598 22554 -14190
rect 22596 -14242 23404 -14230
rect 22596 -14542 22608 -14242
rect 23388 -14298 23404 -14242
rect 23390 -14316 23404 -14298
rect 23524 -14238 24332 -14230
rect 23524 -14316 23538 -14238
rect 23390 -14482 23538 -14316
rect 23390 -14504 23404 -14482
rect 23388 -14542 23404 -14504
rect 22596 -14554 23404 -14542
rect 23524 -14538 23538 -14482
rect 24318 -14316 24332 -14238
rect 24376 -14268 24478 -14190
rect 24548 -14316 24616 -13326
rect 24318 -14482 24616 -14316
rect 24318 -14538 24332 -14482
rect 23524 -14554 24332 -14538
rect 24376 -14598 24478 -14532
rect 22452 -14766 24478 -14598
rect 22452 -14834 22554 -14766
rect 22596 -14814 23404 -14802
rect 22596 -14884 22610 -14814
rect 22240 -14976 22610 -14884
rect 23390 -14976 23404 -14814
rect 22240 -14982 23404 -14976
rect 23552 -14908 24300 -14894
rect 22452 -15184 22554 -15040
rect 22452 -15352 23448 -15184
rect 22452 -15560 22554 -15352
rect 22452 -15590 23486 -15560
rect 21956 -15598 23486 -15590
rect 21956 -15642 22612 -15598
rect 23390 -15642 23486 -15598
rect 23552 -15622 23570 -14908
rect 24284 -15622 24300 -14908
rect 23552 -15638 24300 -15622
rect 21956 -15750 22610 -15642
rect 21520 -16266 21878 -16254
rect 22452 -15914 22610 -15750
rect 23392 -15752 23486 -15642
rect 24376 -15752 24478 -14766
rect 23392 -15914 24478 -15752
rect 22452 -15920 24478 -15914
rect 22452 -15946 23486 -15920
rect 22452 -16332 22554 -15946
rect 22596 -15988 23404 -15978
rect 22596 -16288 22610 -15988
rect 23390 -16050 23404 -15988
rect 23522 -15988 24330 -15978
rect 23522 -16050 23538 -15988
rect 23390 -16216 23538 -16050
rect 23390 -16288 23404 -16216
rect 22596 -16302 23404 -16288
rect 23522 -16288 23538 -16216
rect 24318 -16050 24330 -15988
rect 24376 -16000 24478 -15920
rect 24548 -16050 24616 -14482
rect 24318 -16216 24616 -16050
rect 24318 -16288 24330 -16216
rect 23522 -16302 24330 -16288
rect 24376 -16332 24478 -16264
rect 22452 -16500 24478 -16332
rect 21704 -16590 22104 -16576
rect 21704 -17098 21718 -16590
rect 22090 -17098 22104 -16590
rect 21704 -17112 22104 -17098
rect 22452 -16906 22554 -16500
rect 22596 -16552 23404 -16540
rect 22596 -16852 22610 -16552
rect 23390 -16628 23404 -16552
rect 23524 -16552 24332 -16540
rect 23524 -16628 23536 -16552
rect 24316 -16604 24332 -16552
rect 23390 -16794 23536 -16628
rect 23390 -16852 23404 -16794
rect 22596 -16864 23404 -16852
rect 23524 -16852 23536 -16794
rect 24318 -16812 24332 -16604
rect 24316 -16852 24332 -16812
rect 23524 -16864 24332 -16852
rect 24376 -16906 24478 -16500
rect 22452 -17074 24478 -16906
rect 20332 -18216 21396 -18116
rect 18850 -18486 20252 -18466
rect 17754 -18590 19608 -18578
rect 17754 -19030 17768 -18590
rect 19592 -19030 19608 -18590
rect 17754 -19040 19608 -19030
rect 19848 -22670 20248 -18486
rect 20776 -20592 20936 -18216
rect 21830 -18388 21990 -17112
rect 22452 -17502 22554 -17074
rect 22596 -17138 23404 -17126
rect 22596 -17438 22610 -17138
rect 23390 -17206 23404 -17138
rect 23524 -17136 24332 -17126
rect 23524 -17206 23538 -17136
rect 23390 -17372 23538 -17206
rect 23390 -17438 23404 -17372
rect 22596 -17450 23404 -17438
rect 23524 -17436 23538 -17372
rect 24318 -17206 24332 -17136
rect 24376 -17158 24478 -17074
rect 24548 -17206 24616 -16216
rect 24318 -17372 24616 -17206
rect 24318 -17436 24332 -17372
rect 23524 -17450 24332 -17436
rect 23442 -17502 23486 -17460
rect 24374 -17502 24376 -17460
rect 22452 -17694 24376 -17502
rect 22452 -17696 23484 -17694
rect 22452 -17736 22560 -17696
rect 23448 -17736 23484 -17696
rect 24372 -17736 24376 -17694
rect 24548 -17820 24616 -17372
rect 22120 -17924 24616 -17820
rect 22120 -17984 25228 -17924
rect 24548 -17986 25228 -17984
rect 21830 -18548 23334 -18388
rect 23174 -18572 23334 -18548
rect 23174 -18732 24982 -18572
rect 23174 -19970 23334 -18732
rect 24530 -19016 24964 -18782
rect 24530 -19348 24964 -19114
rect 24530 -19680 24964 -19446
rect 23102 -19984 23402 -19970
rect 23102 -20260 23114 -19984
rect 23386 -20260 23402 -19984
rect 24530 -20012 24964 -19778
rect 23102 -20270 23402 -20260
rect 20704 -20606 21004 -20592
rect 20704 -20882 20718 -20606
rect 20990 -20882 21004 -20606
rect 20704 -20892 21004 -20882
rect 20776 -22154 20936 -20892
rect 20706 -22168 21006 -22154
rect 20706 -22440 20720 -22168
rect 20992 -22440 21006 -22168
rect 20706 -22454 21006 -22440
rect 1844 -22710 20318 -22670
rect 1844 -23440 1890 -22710
rect 20268 -23440 20318 -22710
rect 20776 -22932 20936 -22454
rect 21474 -22828 22674 -22792
rect 20458 -23032 21408 -22932
rect 20776 -23304 20936 -23032
rect 21474 -23088 21482 -22828
rect 21214 -23096 21482 -23088
rect 21544 -22830 22674 -22828
rect 21544 -23090 22604 -22830
rect 21214 -23158 21226 -23096
rect 21544 -23158 21764 -23090
rect 21214 -23186 21764 -23158
rect 1844 -23486 20318 -23440
rect 20656 -23312 21056 -23304
rect 1772 -23554 20612 -23544
rect 20600 -23656 20612 -23554
rect 1662 -23668 20612 -23656
rect 20656 -23696 20664 -23312
rect 21048 -23696 21056 -23312
rect 21288 -23598 21764 -23186
rect 22366 -23160 22604 -23090
rect 22666 -23090 22674 -22830
rect 23174 -22932 23334 -20270
rect 24530 -20344 24964 -20110
rect 24530 -20676 24964 -20442
rect 24530 -21008 24964 -20774
rect 24528 -21342 24962 -21108
rect 24530 -21672 24964 -21438
rect 24528 -22004 24962 -21770
rect 24528 -22338 24962 -22104
rect 25198 -22706 25228 -17986
rect 24040 -22730 25228 -22706
rect 22740 -23032 23658 -22932
rect 22666 -23098 22934 -23090
rect 22922 -23160 22934 -23098
rect 22366 -23348 22934 -23160
rect 23174 -23304 23334 -23032
rect 24040 -23206 24070 -22730
rect 23544 -23230 24070 -23206
rect 23054 -23316 23454 -23304
rect 22366 -23598 22968 -23348
rect 21288 -23646 22968 -23598
rect 20656 -23704 21056 -23696
rect 23054 -23690 23070 -23316
rect 23440 -23690 23454 -23316
rect 23544 -23630 23578 -23230
rect 25456 -23630 25512 -11668
rect 23544 -23646 25512 -23630
rect 23054 -23704 23454 -23690
<< via1 >>
rect 1638 -1200 2012 -826
rect 2190 -1200 2564 -826
rect 3606 -1200 3980 -826
rect 4350 -1198 4724 -824
rect 3046 -1694 3414 -1690
rect 3046 -1768 3050 -1694
rect 3050 -1768 3412 -1694
rect 3412 -1768 3414 -1694
rect 3046 -1772 3414 -1768
rect 8088 -1200 8464 -822
rect 9982 -882 10370 -818
rect 4912 -1686 5280 -1682
rect 4912 -1760 4916 -1686
rect 4916 -1760 5278 -1686
rect 5278 -1760 5280 -1686
rect 4912 -1764 5280 -1760
rect 3788 -2726 4544 -2044
rect 3880 -2952 4452 -2870
rect 9982 -1206 10370 -882
rect 11200 -1204 11580 -822
rect 12730 -1138 13494 -960
rect 12730 -1262 13372 -1138
rect 13372 -1262 13494 -1138
rect 3880 -3222 4452 -2952
rect 3880 -3308 4452 -3222
rect 1636 -5026 1920 -3600
rect 2048 -5154 2454 -5122
rect 2048 -6772 2454 -5154
rect 2048 -6798 2454 -6772
rect 3952 -6808 4374 -5116
rect 3370 -7222 3478 -6962
rect 3620 -7214 3728 -6954
rect 2412 -7266 2520 -7254
rect 2412 -8042 2420 -7266
rect 2420 -8042 2512 -7266
rect 2512 -8042 2520 -7266
rect 2412 -8054 2520 -8042
rect 2570 -7266 2678 -7254
rect 2570 -8042 2578 -7266
rect 2578 -8042 2670 -7266
rect 2670 -8042 2678 -7266
rect 2570 -8054 2678 -8042
rect 2728 -7266 2836 -7254
rect 2728 -8042 2736 -7266
rect 2736 -8042 2828 -7266
rect 2828 -8042 2836 -7266
rect 2728 -8054 2836 -8042
rect 2886 -7266 2994 -7254
rect 2886 -8042 2894 -7266
rect 2894 -8042 2986 -7266
rect 2986 -8042 2994 -7266
rect 2886 -8054 2994 -8042
rect 3042 -7266 3150 -7254
rect 3042 -8042 3050 -7266
rect 3050 -8042 3142 -7266
rect 3142 -8042 3150 -7266
rect 3042 -8054 3150 -8042
rect 3202 -7266 3310 -7254
rect 3202 -8042 3210 -7266
rect 3210 -8042 3302 -7266
rect 3302 -8042 3310 -7266
rect 3202 -8054 3310 -8042
rect 3370 -8078 3478 -7906
rect 3620 -8078 3728 -7916
rect 3790 -7266 3894 -7254
rect 3790 -8044 3796 -7266
rect 3796 -8044 3888 -7266
rect 3888 -8044 3894 -7266
rect 3790 -8054 3894 -8044
rect 3946 -7266 4054 -7254
rect 3946 -8044 3954 -7266
rect 3954 -8044 4046 -7266
rect 4046 -8044 4054 -7266
rect 3946 -8054 4054 -8044
rect 4104 -7266 4212 -7254
rect 4104 -8044 4112 -7266
rect 4112 -8044 4204 -7266
rect 4204 -8044 4212 -7266
rect 4104 -8054 4212 -8044
rect 4262 -7266 4370 -7254
rect 4262 -8044 4270 -7266
rect 4270 -8044 4362 -7266
rect 4362 -8044 4370 -7266
rect 4262 -8054 4370 -8044
rect 4420 -7266 4528 -7254
rect 4420 -8044 4428 -7266
rect 4428 -8044 4520 -7266
rect 4520 -8044 4528 -7266
rect 4420 -8054 4528 -8044
rect 4578 -7266 4686 -7254
rect 4578 -8044 4586 -7266
rect 4586 -8044 4678 -7266
rect 4678 -8044 4686 -7266
rect 4578 -8054 4686 -8044
rect 7372 -1444 7472 -1344
rect 12358 -1444 12458 -1344
rect 7378 -1600 7478 -1500
rect 12184 -1600 12284 -1500
rect 12730 -1490 13370 -1262
rect 13370 -1490 13494 -1262
rect 7378 -1784 7478 -1684
rect 12006 -1784 12106 -1684
rect 7434 -2198 7550 -2194
rect 7434 -2976 7444 -2198
rect 7444 -2976 7540 -2198
rect 7540 -2976 7550 -2198
rect 7434 -2982 7550 -2976
rect 7594 -2198 7710 -2194
rect 7594 -2976 7604 -2198
rect 7604 -2976 7700 -2198
rect 7700 -2976 7710 -2198
rect 7594 -2982 7710 -2976
rect 7752 -2198 7868 -2194
rect 7752 -2976 7762 -2198
rect 7762 -2976 7858 -2198
rect 7858 -2976 7868 -2198
rect 7752 -2982 7868 -2976
rect 7910 -2198 8026 -2194
rect 7910 -2976 7920 -2198
rect 7920 -2976 8016 -2198
rect 8016 -2976 8026 -2198
rect 7910 -2982 8026 -2976
rect 8068 -2198 8184 -2194
rect 8068 -2976 8078 -2198
rect 8078 -2976 8174 -2198
rect 8174 -2976 8184 -2198
rect 8068 -2982 8184 -2976
rect 8224 -2198 8340 -2192
rect 8224 -2976 8234 -2198
rect 8234 -2976 8330 -2198
rect 8330 -2976 8340 -2198
rect 8224 -2980 8340 -2976
rect 8382 -2198 8498 -2194
rect 8382 -2976 8392 -2198
rect 8392 -2976 8488 -2198
rect 8488 -2976 8498 -2198
rect 8382 -2982 8498 -2976
rect 8542 -2198 8658 -2192
rect 8542 -2976 8552 -2198
rect 8552 -2976 8648 -2198
rect 8648 -2976 8658 -2198
rect 8542 -2980 8658 -2976
rect 8698 -2198 8814 -2194
rect 8698 -2976 8708 -2198
rect 8708 -2976 8804 -2198
rect 8804 -2976 8814 -2198
rect 8698 -2982 8814 -2976
rect 8856 -2198 8972 -2194
rect 8856 -2976 8866 -2198
rect 8866 -2976 8962 -2198
rect 8962 -2976 8972 -2198
rect 8856 -2982 8972 -2976
rect 9014 -2198 9130 -2194
rect 9014 -2976 9024 -2198
rect 9024 -2976 9120 -2198
rect 9120 -2976 9130 -2198
rect 9014 -2982 9130 -2976
rect 9360 -2202 9476 -2198
rect 9360 -2980 9370 -2202
rect 9370 -2980 9466 -2202
rect 9466 -2980 9476 -2202
rect 9360 -2986 9476 -2980
rect 9518 -2202 9634 -2198
rect 9518 -2980 9528 -2202
rect 9528 -2980 9624 -2202
rect 9624 -2980 9634 -2202
rect 9518 -2986 9634 -2980
rect 9678 -2202 9794 -2198
rect 9678 -2980 9688 -2202
rect 9688 -2980 9784 -2202
rect 9784 -2980 9794 -2202
rect 9678 -2986 9794 -2980
rect 9836 -2202 9952 -2198
rect 9836 -2980 9846 -2202
rect 9846 -2980 9942 -2202
rect 9942 -2980 9952 -2202
rect 9836 -2986 9952 -2980
rect 9992 -2202 10108 -2198
rect 9992 -2980 10002 -2202
rect 10002 -2980 10098 -2202
rect 10098 -2980 10108 -2202
rect 9992 -2986 10108 -2980
rect 10152 -2202 10268 -2198
rect 10152 -2980 10162 -2202
rect 10162 -2980 10258 -2202
rect 10258 -2980 10268 -2202
rect 10152 -2986 10268 -2980
rect 10308 -2202 10424 -2198
rect 10308 -2980 10318 -2202
rect 10318 -2980 10414 -2202
rect 10414 -2980 10424 -2202
rect 10308 -2986 10424 -2980
rect 10466 -2202 10582 -2198
rect 10466 -2980 10476 -2202
rect 10476 -2980 10572 -2202
rect 10572 -2980 10582 -2202
rect 10466 -2986 10582 -2980
rect 10626 -2202 10742 -2198
rect 10626 -2980 10636 -2202
rect 10636 -2980 10732 -2202
rect 10732 -2980 10742 -2202
rect 10626 -2986 10742 -2980
rect 10782 -2202 10898 -2198
rect 10782 -2980 10792 -2202
rect 10792 -2980 10888 -2202
rect 10888 -2980 10898 -2202
rect 10782 -2986 10898 -2980
rect 10940 -2202 11056 -2198
rect 10940 -2980 10950 -2202
rect 10950 -2980 11046 -2202
rect 11046 -2980 11056 -2202
rect 10940 -2986 11056 -2980
rect 11310 -2180 11462 -2176
rect 11310 -2958 11462 -2180
rect 11310 -2964 11462 -2958
rect 11780 -3164 11972 -2980
rect 11426 -3386 11604 -3208
rect 13942 -3470 14128 -3124
rect 14344 -3464 14520 -3152
rect 16124 -3514 16212 -3136
rect 16212 -3514 17524 -3136
rect 23924 -1200 24302 -820
rect 9146 -4152 9246 -4052
rect 11462 -4152 11562 -4052
rect 12112 -4316 15250 -4310
rect 9534 -4734 10888 -4324
rect 9534 -4970 10462 -4734
rect 10462 -4970 10476 -4734
rect 11780 -4810 11972 -4626
rect 12112 -4750 15250 -4316
rect 12112 -4760 15250 -4750
rect 9534 -5346 11224 -4970
rect 12122 -5346 12488 -4970
rect 12924 -5346 13168 -4970
rect 13276 -5346 13642 -4970
rect 14538 -5346 15284 -4970
rect 17508 -4750 17702 -4742
rect 17508 -5526 17514 -4750
rect 17514 -5004 17702 -4750
rect 17514 -5526 18002 -5004
rect 17508 -5530 18002 -5526
rect 7604 -5640 8962 -5608
rect 7604 -7366 8878 -5640
rect 8878 -7366 8962 -5640
rect 11666 -6000 11814 -5990
rect 11666 -6378 11814 -6000
rect 11666 -6388 11814 -6378
rect 11666 -6528 11814 -6518
rect 11666 -6906 11814 -6528
rect 11666 -6916 11814 -6906
rect 12924 -6392 13250 -5982
rect 12924 -6468 13250 -6392
rect 12810 -6528 12958 -6518
rect 12810 -6906 12958 -6528
rect 12810 -6916 12958 -6906
rect 13954 -6000 14102 -5990
rect 13954 -6378 14102 -6000
rect 13954 -6388 14102 -6378
rect 13954 -6528 14102 -6518
rect 13954 -6906 14102 -6528
rect 13954 -6916 14102 -6906
rect 16044 -7036 16148 -6554
rect 17014 -6890 17280 -6106
rect 19090 -5706 19230 -5466
rect 17528 -6108 17782 -6100
rect 17528 -6886 17532 -6108
rect 17532 -6886 17782 -6108
rect 17528 -6894 17782 -6886
rect 18146 -7036 18250 -6554
rect 20580 -6104 20668 -6016
rect 19092 -6714 19232 -6474
rect 21468 -5788 21556 -5334
rect 21470 -6820 21560 -6330
rect 23006 -5246 23868 -4406
rect 22006 -6124 22302 -5996
rect 22726 -6132 23002 -5852
rect 24796 -5830 25120 -4334
rect 24010 -6130 24210 -5930
rect 22262 -7202 24596 -6846
rect 7604 -7438 8962 -7366
rect 24230 -7540 24644 -7402
rect 9636 -9408 10048 -9406
rect 9636 -9922 10048 -9408
rect 24792 -10142 25112 -7416
rect 24792 -10144 25112 -10142
rect 15988 -11130 16648 -10464
rect 17142 -10898 18052 -10464
rect 2030 -11824 3298 -11314
rect 15036 -11798 15812 -11484
rect 17714 -11798 18284 -11310
rect 2030 -11974 3298 -11824
rect 2032 -12806 3288 -11974
rect 2032 -13766 2930 -12806
rect 15036 -12058 15812 -11798
rect 17714 -12066 18284 -11798
rect 7542 -12430 7704 -12270
rect 9998 -12434 11440 -12268
rect 11662 -12434 13104 -12268
rect 20292 -12468 20464 -12298
rect 7346 -12910 7506 -12620
rect 16050 -14472 16548 -13980
rect 18384 -14132 19346 -13994
rect 18384 -14456 18848 -14132
rect 19712 -14762 19844 -13440
rect 20214 -14482 20590 -13716
rect 20882 -14052 21736 -14030
rect 20882 -14306 20916 -14052
rect 20916 -14306 21698 -14052
rect 21698 -14306 21736 -14052
rect 22612 -13924 23390 -13716
rect 23540 -13716 24316 -13714
rect 24316 -13716 24318 -13714
rect 23540 -13922 24318 -13716
rect 18420 -15530 18784 -15164
rect 2148 -22372 2654 -22232
rect 19884 -17992 20222 -16020
rect 20476 -16268 21250 -16010
rect 20474 -16332 21252 -16324
rect 20474 -16424 20476 -16332
rect 20476 -16424 21252 -16332
rect 20474 -16430 21252 -16424
rect 20474 -16490 21252 -16482
rect 20474 -16582 20476 -16490
rect 20476 -16582 21252 -16490
rect 20474 -16588 21252 -16582
rect 20474 -16648 21252 -16640
rect 20474 -16740 20476 -16648
rect 20476 -16740 21252 -16648
rect 20474 -16746 21252 -16740
rect 20474 -16806 21252 -16798
rect 20474 -16898 20476 -16806
rect 20476 -16898 21252 -16806
rect 20474 -16904 21252 -16898
rect 20474 -16964 21252 -16956
rect 20474 -17056 20476 -16964
rect 20476 -17056 21252 -16964
rect 20474 -17062 21252 -17056
rect 20476 -17122 21254 -17114
rect 20476 -17214 21252 -17122
rect 21252 -17214 21254 -17122
rect 20476 -17220 21254 -17214
rect 20474 -17280 21252 -17272
rect 20474 -17372 20476 -17280
rect 20476 -17372 21252 -17280
rect 20474 -17378 21252 -17372
rect 20474 -17438 21252 -17430
rect 20474 -17530 20476 -17438
rect 20476 -17530 21252 -17438
rect 20474 -17536 21252 -17530
rect 20474 -17596 21252 -17588
rect 20474 -17688 20476 -17596
rect 20476 -17688 21252 -17596
rect 20474 -17694 21252 -17688
rect 20476 -17756 21250 -17750
rect 20476 -18008 21250 -17756
rect 23628 -15592 24228 -14938
rect 21718 -17098 22090 -16590
rect 22610 -16812 23388 -16604
rect 23540 -16606 24316 -16604
rect 24316 -16606 24318 -16604
rect 23540 -16812 24318 -16606
rect 17768 -19030 19592 -18590
rect 23114 -20260 23386 -19984
rect 20718 -20882 20990 -20606
rect 20720 -22440 20992 -22168
rect 20664 -23696 21048 -23312
rect 23070 -23690 23440 -23316
<< metal2 >>
rect 1626 -826 2026 -812
rect 1626 -1200 1638 -826
rect 2012 -1200 2026 -826
rect 1626 -1212 2026 -1200
rect 2178 -826 2578 -812
rect 2178 -1200 2190 -826
rect 2564 -1200 2578 -826
rect 2178 -1212 2578 -1200
rect 3592 -826 3992 -812
rect 3592 -1200 3606 -826
rect 3980 -1200 3992 -826
rect 3592 -1212 3992 -1200
rect 4338 -824 4738 -812
rect 4338 -1198 4350 -824
rect 4724 -1198 4738 -824
rect 4338 -1212 4738 -1198
rect 8076 -822 8476 -812
rect 8076 -1200 8088 -822
rect 8464 -1200 8476 -822
rect 8076 -1210 8476 -1200
rect 9976 -818 10376 -812
rect 9976 -1206 9982 -818
rect 10370 -1206 10376 -818
rect 9976 -1210 10376 -1206
rect 11192 -822 11592 -812
rect 11192 -1204 11200 -822
rect 11580 -1204 11592 -822
rect 23912 -820 24312 -812
rect 14082 -936 23806 -852
rect 1626 -3600 1926 -1212
rect 2226 -1362 2526 -1212
rect 7542 -1220 9136 -1210
rect 1626 -7264 1636 -3600
rect 1920 -5026 1926 -3600
rect 1830 -6974 1926 -5026
rect 2026 -1662 2526 -1362
rect 6632 -1444 7372 -1344
rect 7472 -1444 7478 -1344
rect 2026 -5102 2326 -1662
rect 6632 -1672 6732 -1444
rect 3038 -1690 4632 -1680
rect 3038 -1772 3046 -1690
rect 3414 -1772 4632 -1690
rect 4904 -1682 6732 -1672
rect 4904 -1764 4912 -1682
rect 5280 -1764 6732 -1682
rect 4904 -1772 6732 -1764
rect 6812 -1600 7378 -1500
rect 7478 -1600 7484 -1500
rect 7542 -1562 7548 -1220
rect 9128 -1562 9136 -1220
rect 3038 -1780 4632 -1772
rect 4532 -1864 4632 -1780
rect 6812 -1864 6912 -1600
rect 4532 -1964 6912 -1864
rect 6974 -1784 7378 -1684
rect 7478 -1784 7484 -1684
rect 6974 -2026 7074 -1784
rect 7542 -1854 9136 -1562
rect 3772 -2044 4562 -2026
rect 3772 -2272 3788 -2044
rect 3770 -2726 3788 -2272
rect 4544 -2726 4562 -2044
rect 3770 -2742 4562 -2726
rect 6042 -2126 7074 -2026
rect 7428 -2084 9136 -1854
rect 3864 -2870 4470 -2854
rect 3864 -3308 3880 -2870
rect 4452 -3308 4470 -2870
rect 6042 -3082 6142 -2126
rect 7428 -2194 7556 -2084
rect 7428 -2982 7434 -2194
rect 7550 -2982 7556 -2194
rect 7428 -2992 7556 -2982
rect 7588 -2194 7716 -2184
rect 7588 -2982 7594 -2194
rect 7710 -2982 7716 -2194
rect 5274 -3182 6142 -3082
rect 7588 -3092 7716 -2982
rect 7746 -2194 7874 -2084
rect 7746 -2982 7752 -2194
rect 7868 -2982 7874 -2194
rect 7746 -2992 7874 -2982
rect 7904 -2194 8032 -2184
rect 7904 -2982 7910 -2194
rect 8026 -2982 8032 -2194
rect 7904 -3092 8032 -2982
rect 8062 -2194 8190 -2084
rect 8062 -2982 8068 -2194
rect 8184 -2982 8190 -2194
rect 8062 -2992 8190 -2982
rect 8218 -2192 8346 -2184
rect 8218 -2980 8224 -2192
rect 8340 -2980 8346 -2192
rect 8218 -3092 8346 -2980
rect 8376 -2194 8504 -2084
rect 8376 -2982 8382 -2194
rect 8498 -2982 8504 -2194
rect 8376 -2992 8504 -2982
rect 8536 -2192 8664 -2184
rect 8536 -2980 8542 -2192
rect 8658 -2980 8664 -2192
rect 8536 -3092 8664 -2980
rect 8692 -2194 8820 -2084
rect 8692 -2982 8698 -2194
rect 8814 -2982 8820 -2194
rect 8692 -2992 8820 -2982
rect 8850 -2194 8978 -2184
rect 8850 -2982 8856 -2194
rect 8972 -2982 8978 -2194
rect 8850 -3092 8978 -2982
rect 9008 -2194 9136 -2084
rect 9008 -2982 9014 -2194
rect 9130 -2982 9136 -2194
rect 9008 -2992 9136 -2982
rect 9354 -1238 11062 -1210
rect 11192 -1212 11592 -1204
rect 12712 -960 13510 -946
rect 9354 -1640 9390 -1238
rect 11028 -1640 11062 -1238
rect 9354 -2088 11062 -1640
rect 9354 -2198 9482 -2088
rect 9354 -2986 9360 -2198
rect 9476 -2986 9482 -2198
rect 9354 -2996 9482 -2986
rect 9512 -2198 9640 -2188
rect 9512 -2986 9518 -2198
rect 9634 -2986 9640 -2198
rect 3864 -3324 4470 -3308
rect 2026 -5122 2480 -5102
rect 2026 -6798 2048 -5122
rect 2454 -6798 2480 -5122
rect 3940 -5116 4386 -5102
rect 2026 -6822 2480 -6798
rect 2610 -6860 3484 -6740
rect 3364 -6962 3484 -6860
rect 1830 -7174 3158 -6974
rect 1830 -7254 2526 -7174
rect 2722 -7254 2842 -7174
rect 3036 -7254 3158 -7174
rect 3364 -7222 3370 -6962
rect 3478 -7222 3484 -6962
rect 1830 -7264 2412 -7254
rect 1626 -7274 2412 -7264
rect 2406 -8054 2412 -7274
rect 2520 -8054 2526 -7254
rect 2564 -8054 2570 -7254
rect 2678 -8054 2684 -7254
rect 2722 -8054 2728 -7254
rect 2836 -8054 2842 -7254
rect 2880 -8054 2886 -7254
rect 2994 -8054 3000 -7254
rect 3036 -8054 3042 -7254
rect 3150 -7554 3158 -7254
rect 3150 -8054 3156 -7554
rect 3196 -8054 3202 -7254
rect 3310 -8054 3316 -7254
rect 2564 -8134 2684 -8054
rect 2880 -8134 3000 -8054
rect 3196 -8134 3316 -8054
rect 3364 -7906 3484 -7222
rect 3364 -8078 3370 -7906
rect 3478 -8078 3484 -7906
rect 3614 -6954 3734 -6750
rect 3614 -7214 3620 -6954
rect 3728 -7214 3734 -6954
rect 3614 -7916 3734 -7214
rect 3940 -6808 3952 -5116
rect 4374 -6808 4386 -5116
rect 7588 -5608 8978 -3092
rect 9512 -3096 9640 -2986
rect 9672 -2198 9800 -2088
rect 9672 -2986 9678 -2198
rect 9794 -2986 9800 -2198
rect 9672 -2996 9800 -2986
rect 9830 -2198 9958 -2188
rect 9830 -2986 9836 -2198
rect 9952 -2986 9958 -2198
rect 9830 -3096 9958 -2986
rect 9986 -2198 10114 -2088
rect 9986 -2986 9992 -2198
rect 10108 -2986 10114 -2198
rect 9986 -2996 10114 -2986
rect 10146 -2198 10274 -2188
rect 10146 -2986 10152 -2198
rect 10268 -2986 10274 -2198
rect 10146 -3096 10274 -2986
rect 10302 -2198 10430 -2088
rect 10302 -2986 10308 -2198
rect 10424 -2986 10430 -2198
rect 10302 -2996 10430 -2986
rect 10460 -2198 10588 -2188
rect 10460 -2986 10466 -2198
rect 10582 -2986 10588 -2198
rect 10460 -3096 10588 -2986
rect 10620 -2198 10748 -2088
rect 10620 -2986 10626 -2198
rect 10742 -2986 10748 -2198
rect 10620 -2996 10748 -2986
rect 10776 -2198 10904 -2188
rect 10776 -2986 10782 -2198
rect 10898 -2986 10904 -2198
rect 10776 -3096 10904 -2986
rect 10934 -2198 11062 -2088
rect 10934 -2986 10940 -2198
rect 11056 -2986 11062 -2198
rect 11300 -2176 11474 -1212
rect 12358 -1344 12458 -1338
rect 12184 -1500 12284 -1494
rect 12006 -1684 12106 -1678
rect 12006 -1874 12106 -1784
rect 12184 -1736 12284 -1600
rect 12358 -1586 12458 -1444
rect 12712 -1490 12730 -960
rect 13494 -1490 13510 -960
rect 12712 -1504 13510 -1490
rect 14082 -1508 15334 -936
rect 15922 -1508 23806 -936
rect 23912 -1200 23924 -820
rect 24302 -1200 24312 -820
rect 23912 -1212 24312 -1200
rect 14082 -1530 23806 -1508
rect 14434 -1532 23806 -1530
rect 12358 -1686 13790 -1586
rect 12184 -1836 13542 -1736
rect 12006 -1974 13372 -1874
rect 11300 -2964 11310 -2176
rect 11462 -2964 11474 -2176
rect 13272 -2204 13372 -1974
rect 13442 -1926 13542 -1836
rect 15402 -1838 23806 -1532
rect 13442 -2026 13808 -1926
rect 15402 -2058 21844 -1838
rect 13272 -2304 13800 -2204
rect 11300 -2974 11474 -2964
rect 16192 -2550 21842 -2532
rect 10934 -2996 11062 -2986
rect 11772 -2980 11980 -2972
rect 5526 -6710 5726 -6660
rect 3940 -7014 4000 -6808
rect 4308 -6974 4386 -6808
rect 5592 -6810 5692 -6710
rect 5526 -6860 5726 -6810
rect 4308 -7014 4692 -6974
rect 3940 -7174 4692 -7014
rect 3940 -7254 4060 -7174
rect 4256 -7254 4376 -7174
rect 4572 -7254 4692 -7174
rect 3614 -8078 3620 -7916
rect 3728 -8078 3734 -7916
rect 3782 -8054 3790 -7254
rect 3894 -8054 3902 -7254
rect 3940 -8054 3946 -7254
rect 4054 -8054 4060 -7254
rect 4098 -8054 4104 -7254
rect 4212 -8054 4218 -7254
rect 4256 -8054 4262 -7254
rect 4370 -8054 4376 -7254
rect 4414 -8054 4420 -7254
rect 4528 -8054 4534 -7254
rect 4572 -8054 4578 -7254
rect 4686 -8054 4692 -7254
rect 5592 -7536 5692 -6860
rect 7588 -7438 7604 -5608
rect 8962 -7438 8978 -5608
rect 7588 -7454 8978 -7438
rect 9146 -4052 9246 -4046
rect 9146 -7536 9246 -4152
rect 9512 -4324 10904 -3096
rect 11772 -3164 11780 -2980
rect 11972 -3164 11980 -2980
rect 16192 -3006 16208 -2550
rect 17532 -2752 21842 -2550
rect 22136 -2752 23806 -1838
rect 17532 -3006 23812 -2752
rect 16192 -3022 23812 -3006
rect 11772 -3172 11980 -3164
rect 13934 -3124 14136 -3116
rect 11416 -3208 11616 -3198
rect 11416 -3386 11426 -3208
rect 11604 -3386 11616 -3208
rect 11416 -3398 11616 -3386
rect 11462 -4052 11568 -3398
rect 11562 -4152 11568 -4052
rect 11462 -4156 11568 -4152
rect 11462 -4158 11562 -4156
rect 9512 -5346 9534 -4324
rect 10888 -4734 10904 -4324
rect 11826 -4616 11926 -3172
rect 13934 -3470 13942 -3124
rect 14128 -3470 14136 -3124
rect 16104 -3136 17546 -3120
rect 13934 -3476 14136 -3470
rect 14332 -3152 14532 -3140
rect 14332 -3464 14344 -3152
rect 14520 -3464 14532 -3152
rect 14332 -3476 14532 -3464
rect 13962 -3882 14102 -3476
rect 14360 -3640 14500 -3476
rect 16104 -3514 16124 -3136
rect 17524 -3514 17546 -3136
rect 16104 -3534 17546 -3514
rect 17668 -3530 23812 -3022
rect 14360 -3780 22856 -3640
rect 13962 -4022 22308 -3882
rect 12104 -4310 15264 -4298
rect 10476 -4958 10904 -4734
rect 11772 -4626 11980 -4616
rect 11772 -4810 11780 -4626
rect 11972 -4810 11980 -4626
rect 11772 -4816 11980 -4810
rect 12104 -4760 12112 -4310
rect 15250 -4760 15264 -4310
rect 12104 -4768 15264 -4760
rect 17500 -4742 17712 -4734
rect 12104 -4958 12504 -4768
rect 13260 -4958 13660 -4768
rect 10476 -4970 12504 -4958
rect 11224 -5346 12122 -4970
rect 12488 -5346 12504 -4970
rect 9512 -5358 12504 -5346
rect 12918 -4970 13178 -4958
rect 12918 -5346 12924 -4970
rect 13168 -5346 13178 -4970
rect 12918 -5358 13178 -5346
rect 13260 -4970 15296 -4958
rect 13260 -5346 13276 -4970
rect 13642 -5346 14538 -4970
rect 15284 -5346 15296 -4970
rect 17500 -4994 17508 -4742
rect 13260 -5358 15296 -5346
rect 17212 -5014 17508 -4994
rect 17702 -4994 17712 -4742
rect 17702 -5004 18012 -4994
rect 5592 -7636 9246 -7536
rect 2564 -8280 3316 -8134
rect 3782 -8134 3902 -8054
rect 4098 -8134 4218 -8054
rect 4414 -8134 4534 -8054
rect 2018 -10686 3318 -8280
rect 3782 -8282 4534 -8134
rect 2016 -11314 3318 -10686
rect 3780 -10450 5080 -8282
rect 9616 -9406 10068 -5358
rect 12998 -5896 13098 -5358
rect 17212 -5772 17232 -5014
rect 18002 -5530 18012 -5004
rect 21462 -5334 21562 -5328
rect 17990 -5772 18012 -5530
rect 17212 -5794 18012 -5772
rect 19082 -5466 19242 -5462
rect 19082 -5706 19090 -5466
rect 19230 -5706 19242 -5466
rect 12912 -5982 13260 -5896
rect 11660 -5990 11820 -5984
rect 11660 -6388 11666 -5990
rect 11814 -6388 11820 -5990
rect 11660 -6512 11820 -6388
rect 12912 -6468 12924 -5982
rect 13250 -6468 13260 -5982
rect 12912 -6482 13260 -6468
rect 13948 -5990 14108 -5984
rect 13948 -6388 13954 -5990
rect 14102 -6388 14108 -5990
rect 17500 -6092 17712 -5794
rect 19082 -6036 19242 -5706
rect 21462 -5788 21468 -5334
rect 21556 -5788 21562 -5334
rect 21462 -5794 21562 -5788
rect 21466 -6010 21562 -5794
rect 22168 -5990 22308 -4022
rect 22716 -5842 22856 -3780
rect 22972 -4394 23904 -4378
rect 22972 -4406 23036 -4394
rect 23488 -4406 23904 -4394
rect 22972 -5246 23006 -4406
rect 23868 -5246 23904 -4406
rect 22972 -5266 23036 -5246
rect 23488 -5266 23904 -5246
rect 22972 -5276 23904 -5266
rect 13948 -6402 14108 -6388
rect 16998 -6106 17298 -6092
rect 16998 -6402 17014 -6106
rect 13948 -6502 17014 -6402
rect 13948 -6512 14108 -6502
rect 11660 -6518 14108 -6512
rect 11660 -6916 11666 -6518
rect 11814 -6916 12810 -6518
rect 12958 -6916 13954 -6518
rect 14102 -6916 14108 -6518
rect 11660 -6922 14108 -6916
rect 16036 -6554 16156 -6544
rect 16036 -7036 16044 -6554
rect 16148 -7036 16156 -6554
rect 16998 -6890 17014 -6502
rect 17280 -6890 17298 -6106
rect 16998 -6902 17298 -6890
rect 17500 -6100 17790 -6092
rect 17500 -6894 17528 -6100
rect 17782 -6894 17790 -6100
rect 17500 -6902 17790 -6894
rect 17854 -6196 19242 -6036
rect 20574 -6016 21562 -6010
rect 20574 -6104 20580 -6016
rect 20668 -6104 21562 -6016
rect 20574 -6110 21562 -6104
rect 16036 -7424 16156 -7036
rect 16036 -7544 16904 -7424
rect 9616 -9922 9636 -9406
rect 10048 -9922 10068 -9406
rect 9616 -9948 10068 -9922
rect 3780 -10464 16668 -10450
rect 3780 -10468 15988 -10464
rect 3780 -11132 5904 -10468
rect 7226 -11124 12774 -10468
rect 13664 -11124 15988 -10468
rect 7226 -11130 15988 -11124
rect 16648 -11130 16668 -10464
rect 7226 -11132 16668 -11130
rect 3780 -11150 16668 -11132
rect 2016 -11974 2030 -11314
rect 3298 -11974 3318 -11314
rect 15028 -11482 15826 -11470
rect 15028 -11484 15304 -11482
rect 15554 -11484 15826 -11482
rect 2016 -13536 2032 -11974
rect 3288 -11990 3318 -11974
rect 5808 -11778 7106 -11760
rect 5808 -11790 7984 -11778
rect 3288 -12806 3304 -11990
rect 5808 -12116 5830 -11790
rect 7082 -11968 7984 -11790
rect 7082 -12116 7106 -11968
rect 5808 -12148 7106 -12116
rect 7534 -12270 7714 -12260
rect 7534 -12430 7542 -12270
rect 7704 -12272 7714 -12270
rect 7816 -12272 7984 -11968
rect 15028 -12058 15036 -11484
rect 15812 -12058 15826 -11484
rect 9978 -12268 13126 -12252
rect 9978 -12272 9998 -12268
rect 7704 -12428 9998 -12272
rect 7704 -12430 7714 -12428
rect 7534 -12440 7714 -12430
rect 9978 -12434 9998 -12428
rect 11440 -12434 11662 -12268
rect 13104 -12434 13126 -12268
rect 15028 -12262 15304 -12058
rect 15554 -12262 15826 -12058
rect 15028 -12272 15826 -12262
rect 9978 -12452 13126 -12434
rect 1900 -13570 2032 -13536
rect 2930 -13536 3304 -12806
rect 7334 -12620 7520 -12612
rect 7334 -12910 7346 -12620
rect 7506 -12910 7520 -12620
rect 2930 -13570 3682 -13536
rect 1900 -14770 1946 -13570
rect 3638 -14770 3682 -13570
rect 7334 -13976 7520 -12910
rect 7334 -13978 9618 -13976
rect 16042 -13978 16556 -13972
rect 7334 -13980 16556 -13978
rect 7334 -14146 16050 -13980
rect 7334 -14148 9618 -14146
rect 7334 -14154 7520 -14148
rect 16042 -14472 16050 -14146
rect 16548 -14472 16556 -13980
rect 16042 -14480 16556 -14472
rect 1900 -14810 3682 -14770
rect 16784 -20684 16904 -7544
rect 17854 -7546 18014 -6196
rect 19082 -6474 19242 -6196
rect 21466 -6324 21562 -6110
rect 22000 -5996 22308 -5990
rect 22000 -6124 22006 -5996
rect 22302 -6124 22308 -5996
rect 22000 -6130 22308 -6124
rect 22714 -5852 23014 -5842
rect 22714 -6132 22726 -5852
rect 23002 -6132 23014 -5852
rect 24010 -5930 24210 -1212
rect 24762 -4334 25158 -4298
rect 24762 -5830 24796 -4334
rect 25120 -5830 25158 -4334
rect 24004 -6130 24010 -5930
rect 24210 -6130 24216 -5930
rect 22714 -6142 23014 -6132
rect 17214 -7568 18014 -7546
rect 17214 -8326 17236 -7568
rect 17994 -8326 18014 -7568
rect 17214 -8346 18014 -8326
rect 18138 -6554 18258 -6546
rect 18138 -7036 18146 -6554
rect 18250 -7036 18258 -6554
rect 17112 -10446 18066 -10434
rect 17112 -10904 17124 -10446
rect 17812 -10464 18066 -10446
rect 18052 -10898 18066 -10464
rect 17812 -10904 18066 -10898
rect 17112 -10906 18066 -10904
rect 18138 -10970 18258 -7036
rect 19082 -6714 19092 -6474
rect 19232 -6714 19242 -6474
rect 19082 -7390 19242 -6714
rect 21464 -6330 21564 -6324
rect 21464 -6820 21470 -6330
rect 21560 -6820 21564 -6330
rect 21464 -6826 21564 -6820
rect 22244 -6836 24622 -6828
rect 22244 -6846 22880 -6836
rect 23376 -6846 24622 -6836
rect 22244 -7202 22262 -6846
rect 24596 -7202 24622 -6846
rect 22244 -7224 24622 -7202
rect 19082 -7402 24654 -7390
rect 19082 -7540 24230 -7402
rect 24644 -7540 24654 -7402
rect 19082 -7550 24654 -7540
rect 24762 -7416 25158 -5830
rect 24762 -10144 24792 -7416
rect 25112 -10144 25158 -7416
rect 24762 -10176 25158 -10144
rect 17400 -11090 18258 -10970
rect 17400 -20062 17520 -11090
rect 17700 -11310 18300 -11292
rect 17700 -12066 17714 -11310
rect 18284 -12066 18300 -11310
rect 17700 -15994 18300 -12066
rect 20278 -12298 20478 -12284
rect 20278 -12468 20292 -12298
rect 20464 -12468 20478 -12298
rect 20278 -12484 20478 -12468
rect 19698 -13440 19858 -13426
rect 19698 -13978 19712 -13440
rect 18372 -13994 19712 -13978
rect 18372 -14456 18384 -13994
rect 19346 -14132 19712 -13994
rect 18848 -14146 19712 -14132
rect 18848 -14456 18870 -14146
rect 18372 -14466 18870 -14456
rect 19698 -14762 19712 -14146
rect 19844 -14762 19858 -13440
rect 20328 -13702 20478 -12484
rect 20200 -13716 20600 -13702
rect 20200 -14482 20214 -13716
rect 20590 -14482 20600 -13716
rect 22596 -13714 24330 -13688
rect 22596 -13716 23540 -13714
rect 22596 -13924 22612 -13716
rect 23390 -13922 23540 -13716
rect 24318 -13922 24330 -13714
rect 23390 -13924 24330 -13922
rect 22596 -13956 24330 -13924
rect 20200 -14496 20600 -14482
rect 20856 -14030 21760 -14010
rect 20856 -14306 20882 -14030
rect 21736 -14306 21760 -14030
rect 20856 -14328 21760 -14306
rect 19698 -14776 19858 -14762
rect 20856 -15148 21256 -14328
rect 18402 -15164 21256 -15148
rect 18402 -15530 18420 -15164
rect 18784 -15530 21256 -15164
rect 18402 -15546 21256 -15530
rect 23584 -14938 24274 -13956
rect 18402 -15548 21222 -15546
rect 23584 -15592 23628 -14938
rect 24228 -15592 24274 -14938
rect 17700 -16010 21264 -15994
rect 17700 -16020 20476 -16010
rect 17700 -16410 19884 -16020
rect 17700 -16810 18944 -16410
rect 19854 -16810 19884 -16410
rect 17700 -17210 19884 -16810
rect 17700 -17610 18944 -17210
rect 19854 -17610 19884 -17210
rect 17700 -17992 19884 -17610
rect 20222 -16268 20476 -16020
rect 21250 -16268 21264 -16010
rect 20222 -16284 21264 -16268
rect 20222 -16470 20432 -16284
rect 20464 -16324 21704 -16312
rect 20464 -16430 20474 -16324
rect 21252 -16430 21704 -16324
rect 20464 -16442 21704 -16430
rect 20222 -16482 21264 -16470
rect 20222 -16588 20474 -16482
rect 21252 -16588 21264 -16482
rect 20222 -16600 21264 -16588
rect 21296 -16576 21704 -16442
rect 23584 -16576 24274 -15592
rect 21296 -16590 24330 -16576
rect 20222 -16786 20432 -16600
rect 21296 -16628 21718 -16590
rect 20464 -16640 21718 -16628
rect 20464 -16746 20474 -16640
rect 21252 -16746 21718 -16640
rect 20464 -16758 21718 -16746
rect 20222 -16798 21264 -16786
rect 20222 -16904 20474 -16798
rect 21252 -16904 21264 -16798
rect 20222 -16916 21264 -16904
rect 20222 -17102 20432 -16916
rect 21296 -16944 21718 -16758
rect 20464 -16956 21718 -16944
rect 20464 -17062 20474 -16956
rect 21252 -17062 21718 -16956
rect 20464 -17074 21718 -17062
rect 21296 -17098 21718 -17074
rect 22090 -16604 24330 -16590
rect 22090 -16812 22610 -16604
rect 23388 -16812 23540 -16604
rect 24318 -16812 24330 -16604
rect 22090 -16844 24330 -16812
rect 22090 -17098 22104 -16844
rect 20222 -17114 21264 -17102
rect 20222 -17220 20476 -17114
rect 21254 -17220 21264 -17114
rect 20222 -17232 21264 -17220
rect 21296 -17112 22104 -17098
rect 20222 -17418 20432 -17232
rect 21296 -17260 21704 -17112
rect 20464 -17272 21704 -17260
rect 20464 -17378 20474 -17272
rect 21252 -17378 21704 -17272
rect 20464 -17390 21704 -17378
rect 20222 -17430 21264 -17418
rect 20222 -17536 20474 -17430
rect 21252 -17536 21264 -17430
rect 20222 -17548 21264 -17536
rect 20222 -17734 20432 -17548
rect 21296 -17576 21704 -17390
rect 20464 -17588 21704 -17576
rect 20464 -17694 20474 -17588
rect 21252 -17694 21704 -17588
rect 20464 -17706 21704 -17694
rect 20222 -17750 21264 -17734
rect 20222 -17992 20476 -17750
rect 17700 -18008 20476 -17992
rect 21250 -18008 21264 -17750
rect 17700 -18010 21264 -18008
rect 17700 -18012 18300 -18010
rect 19854 -18022 21264 -18010
rect 17556 -18474 19806 -18462
rect 17556 -18744 17574 -18474
rect 19792 -18744 19806 -18474
rect 17556 -18758 17768 -18744
rect 17680 -19030 17768 -18758
rect 19592 -18758 19806 -18744
rect 19592 -19030 19684 -18758
rect 17680 -19098 19684 -19030
rect 23102 -19984 23402 -19970
rect 23102 -20062 23114 -19984
rect 17400 -20182 23114 -20062
rect 23102 -20260 23114 -20182
rect 23386 -20260 23402 -19984
rect 23102 -20270 23402 -20260
rect 20704 -20606 21004 -20592
rect 20704 -20684 20718 -20606
rect 16784 -20804 20718 -20684
rect 20704 -20882 20718 -20804
rect 20990 -20882 21004 -20606
rect 20704 -20892 21004 -20882
rect 6298 -21038 6540 -21026
rect 6298 -22222 6310 -21038
rect 2136 -22232 6310 -22222
rect 2136 -22372 2148 -22232
rect 2654 -22372 6310 -22232
rect 2136 -22382 6310 -22372
rect 6298 -23318 6310 -22382
rect 6530 -22222 6540 -21038
rect 11016 -21038 11258 -21024
rect 11016 -22222 11030 -21038
rect 6530 -22382 11030 -22222
rect 6530 -23318 6540 -22382
rect 6298 -23330 6540 -23318
rect 11016 -23318 11030 -22382
rect 11250 -22222 11258 -21038
rect 15738 -21036 15980 -21026
rect 15738 -22222 15744 -21036
rect 11250 -22382 15744 -22222
rect 11250 -23318 11258 -22382
rect 11016 -23328 11258 -23318
rect 15738 -23316 15744 -22382
rect 15970 -22222 15980 -21036
rect 20706 -22168 21006 -22154
rect 20706 -22222 20720 -22168
rect 15970 -22382 20720 -22222
rect 15970 -23316 15980 -22382
rect 20706 -22440 20720 -22382
rect 20992 -22440 21006 -22168
rect 20706 -22454 21006 -22440
rect 15738 -23330 15980 -23316
rect 20656 -23312 21056 -23304
rect 20656 -23696 20664 -23312
rect 21048 -23696 21056 -23312
rect 20656 -23704 21056 -23696
rect 23054 -23316 23454 -23304
rect 23054 -23690 23070 -23316
rect 23440 -23690 23454 -23316
rect 23054 -23704 23454 -23690
<< via2 >>
rect 1636 -5026 1830 -3912
rect 1636 -7264 1830 -5026
rect 7548 -1562 9128 -1220
rect 3788 -2726 4544 -2044
rect 3880 -3308 4452 -2870
rect 9390 -1640 11028 -1238
rect 4000 -5886 4308 -5136
rect 3956 -6210 4358 -5886
rect 4000 -6808 4308 -6210
rect 12730 -1490 13494 -960
rect 15334 -1508 15922 -936
rect 4000 -7014 4308 -6808
rect 16208 -3006 17532 -2550
rect 16124 -3514 17524 -3136
rect 17232 -5530 17508 -5014
rect 17508 -5530 17990 -5014
rect 17232 -5772 17990 -5530
rect 23036 -4406 23488 -4394
rect 23036 -5246 23488 -4406
rect 23036 -5266 23488 -5246
rect 5904 -11132 7226 -10468
rect 12774 -11124 13664 -10468
rect 15304 -11484 15554 -11482
rect 5830 -12116 7082 -11790
rect 15304 -11764 15554 -11484
rect 15038 -12026 15810 -11764
rect 15304 -12058 15554 -12026
rect 15304 -12262 15554 -12058
rect 1946 -13766 2032 -13570
rect 2032 -13766 2930 -13570
rect 2930 -13766 3638 -13570
rect 1946 -14770 3638 -13766
rect 16050 -14470 16546 -13980
rect 17236 -8326 17994 -7568
rect 17124 -10464 17812 -10446
rect 17124 -10898 17142 -10464
rect 17142 -10898 17812 -10464
rect 17124 -10904 17812 -10898
rect 22880 -6846 23376 -6836
rect 22880 -7182 23376 -6846
rect 17574 -18590 19792 -18474
rect 17574 -18744 17768 -18590
rect 17768 -18744 19592 -18590
rect 19592 -18744 19792 -18590
rect 6310 -23318 6530 -21038
rect 11030 -23318 11250 -21038
rect 15744 -23316 15970 -21036
<< metal3 >>
rect 15322 -936 15936 -922
rect 12712 -960 13510 -946
rect 7540 -1216 9136 -1210
rect 7540 -1562 7548 -1216
rect 9128 -1562 9136 -1216
rect 7540 -1570 9136 -1562
rect 9356 -1238 11066 -1212
rect 9356 -1640 9390 -1238
rect 11028 -1640 11066 -1238
rect 9356 -1758 11066 -1640
rect 12712 -1490 12730 -960
rect 13494 -1490 13510 -960
rect 12712 -1798 13510 -1490
rect 15322 -1508 15334 -936
rect 15922 -1508 15936 -936
rect 15322 -1520 15936 -1508
rect 3772 -2044 4562 -2026
rect 3772 -2272 3788 -2044
rect 3770 -2726 3788 -2272
rect 4544 -2726 4562 -2044
rect 3770 -2742 4562 -2726
rect 16192 -2550 17548 -2532
rect 3864 -2870 7396 -2854
rect 3864 -3308 3880 -2870
rect 4452 -3308 7396 -2870
rect 16192 -3006 16208 -2550
rect 17532 -3006 17548 -2550
rect 16192 -3022 17548 -3006
rect 3864 -3324 7396 -3308
rect 15918 -3136 17546 -3120
rect 15918 -3514 16124 -3136
rect 17524 -3514 17546 -3136
rect 15918 -3534 17546 -3514
rect 1626 -3906 1842 -3900
rect 1626 -7268 1632 -3906
rect 1836 -7268 1842 -3906
rect 23024 -4394 23524 -4378
rect 17212 -5014 18012 -4994
rect 3886 -5136 4460 -5120
rect 3886 -5886 4000 -5136
rect 4308 -5886 4460 -5136
rect 17212 -5238 17232 -5014
rect 16654 -5538 17232 -5238
rect 17212 -5772 17232 -5538
rect 17990 -5772 18012 -5014
rect 23024 -5266 23036 -4394
rect 23488 -5266 23524 -4394
rect 23024 -5276 23524 -5266
rect 17212 -5794 18012 -5772
rect 3886 -6210 3956 -5886
rect 4358 -6210 4460 -5886
rect 3886 -7014 4000 -6210
rect 4308 -7014 4460 -6210
rect 3886 -7028 4460 -7014
rect 22870 -6836 23384 -6830
rect 22870 -7182 22880 -6836
rect 23376 -7182 23384 -6836
rect 22870 -7190 23384 -7182
rect 1626 -7274 1842 -7268
rect 17214 -7568 18014 -7546
rect 17214 -8326 17236 -7568
rect 17994 -8326 18014 -7568
rect 17214 -8346 18014 -8326
rect 5864 -10412 7262 -10390
rect 5864 -11184 5884 -10412
rect 7244 -11184 7262 -10412
rect 5864 -11204 7262 -11184
rect 12752 -10430 13730 -10410
rect 12752 -11172 12774 -10430
rect 13704 -11172 13730 -10430
rect 17112 -10446 17824 -10432
rect 17112 -10904 17124 -10446
rect 17812 -10904 17824 -10446
rect 17112 -11156 17128 -10904
rect 17808 -11156 17824 -10904
rect 17112 -11168 17824 -11156
rect 12752 -11190 13730 -11172
rect 15026 -11482 15830 -11470
rect 5700 -11790 7106 -11760
rect 5700 -12116 5830 -11790
rect 7082 -12116 7106 -11790
rect 5700 -12148 7106 -12116
rect 15026 -11764 15304 -11482
rect 15554 -11764 15830 -11482
rect 15026 -12026 15038 -11764
rect 15810 -12026 15830 -11764
rect 15026 -12262 15304 -12026
rect 15554 -12262 15830 -12026
rect 15026 -12272 15830 -12262
rect 1898 -13570 3682 -13536
rect 1898 -13572 1946 -13570
rect 3638 -13572 3682 -13570
rect 1898 -14772 1932 -13572
rect 3642 -14772 3682 -13572
rect 1898 -14810 3682 -14772
rect 16042 -13980 16556 -13972
rect 16042 -14470 16050 -13980
rect 16546 -14470 16556 -13980
rect 16042 -15062 16556 -14470
rect 5242 -17098 14268 -16466
rect 17544 -18462 19818 -18448
rect 17544 -18758 17556 -18462
rect 19806 -18758 19818 -18462
rect 17544 -18770 19818 -18758
rect 2044 -21036 24966 -21016
rect 2044 -21038 15744 -21036
rect 2044 -23112 6310 -21038
rect 6298 -23318 6310 -23112
rect 6530 -23112 11030 -21038
rect 6530 -23318 6540 -23112
rect 6298 -23330 6540 -23318
rect 11018 -23318 11030 -23112
rect 11250 -23112 15744 -21038
rect 11250 -23318 11260 -23112
rect 11018 -23326 11260 -23318
rect 15738 -23316 15744 -23112
rect 15970 -21412 24966 -21036
rect 15970 -23112 17354 -21412
rect 15970 -23316 15980 -23112
rect 15738 -23328 15980 -23316
<< via3 >>
rect 7548 -1220 9128 -1216
rect 7548 -1562 9128 -1220
rect 15334 -1508 15922 -936
rect 3788 -2726 4544 -2044
rect 16208 -3006 17532 -2550
rect 1632 -3912 1836 -3906
rect 1632 -7264 1636 -3912
rect 1636 -7264 1830 -3912
rect 1830 -7264 1836 -3912
rect 1632 -7268 1836 -7264
rect 22880 -7182 23376 -6836
rect 17236 -8326 17994 -7568
rect 5884 -10468 7244 -10412
rect 5884 -11132 5904 -10468
rect 5904 -11132 7226 -10468
rect 7226 -11132 7244 -10468
rect 5884 -11184 7244 -11132
rect 12774 -10468 13704 -10430
rect 12774 -11124 13664 -10468
rect 13664 -11124 13704 -10468
rect 12774 -11172 13704 -11124
rect 17128 -10904 17808 -10448
rect 17128 -11156 17808 -10904
rect 1932 -14770 1946 -13572
rect 1946 -14770 3638 -13572
rect 3638 -14770 3642 -13572
rect 1932 -14772 3642 -14770
rect 17556 -18474 19806 -18462
rect 17556 -18744 17574 -18474
rect 17574 -18744 19792 -18474
rect 19792 -18744 19806 -18474
rect 17556 -18758 19806 -18744
<< metal4 >>
rect 15322 -936 15936 -922
rect 7540 -1216 9136 -1210
rect 7540 -1562 7548 -1216
rect 9128 -1562 9136 -1216
rect 7540 -1758 9136 -1562
rect 15322 -1508 15334 -936
rect 15922 -1508 15936 -936
rect 15322 -1792 15936 -1508
rect 3772 -2044 4562 -2026
rect 3772 -2726 3788 -2044
rect 4544 -2272 4562 -2044
rect 4544 -2726 7328 -2272
rect 3772 -2742 7328 -2726
rect 15884 -2550 17548 -2532
rect 15884 -3006 16208 -2550
rect 17532 -3006 17548 -2550
rect 15884 -3022 17548 -3006
rect 1626 -3906 2088 -3900
rect 1626 -7268 1632 -3906
rect 1836 -7268 2088 -3906
rect 1626 -7274 2088 -7268
rect 22664 -6836 23608 -6828
rect 22664 -7182 22880 -6836
rect 23376 -7182 23608 -6836
rect 22664 -7284 23608 -7182
rect 17214 -7568 18014 -7546
rect 17214 -7802 17236 -7568
rect 16472 -8102 17236 -7802
rect 17214 -8326 17236 -8102
rect 17994 -8326 18014 -7568
rect 17214 -8346 18014 -8326
rect 5658 -10412 7262 -10390
rect 5658 -11184 5884 -10412
rect 7244 -11184 7262 -10412
rect 5658 -11204 7262 -11184
rect 12752 -10430 13950 -10410
rect 12752 -11172 12774 -10430
rect 13704 -11172 13950 -10430
rect 15104 -10608 15704 -10396
rect 16932 -10448 17824 -10434
rect 16932 -11156 17128 -10448
rect 17808 -11156 17824 -10448
rect 16932 -11168 17824 -11156
rect 12752 -11190 13950 -11172
rect 14052 -12138 14260 -11586
rect 16656 -12160 16864 -11608
rect 15136 -13354 15736 -13142
rect 1900 -13572 3680 -13538
rect 1900 -14772 1932 -13572
rect 3642 -14772 3680 -13572
rect 1900 -15092 3680 -14772
rect 5242 -17098 14268 -16466
rect 17542 -18462 19822 -18442
rect 17542 -18758 17556 -18462
rect 19806 -18758 19822 -18462
rect 17542 -19024 19822 -18758
rect 5950 -21440 21402 -20766
use sky130_fd_pr__cap_mim_m3_1_67RTNB  amp_XC1
timestamp 1713225924
transform 0 1 12312 -1 0 -8182
box -3798 -4532 6070 4534
use sky130_fd_pr__nfet_g5v0d10v5_Z6W9J4  amp_XM1_2
timestamp 1713225924
transform 1 0 12881 0 1 -5158
box -2451 -458 2451 458
use sky130_fd_pr__pfet_g5v0d10v5_8CDM6Z  amp_XM3_5
timestamp 1713225924
transform 1 0 17147 0 1 -6497
box -1145 -697 1145 697
use sky130_fd_pr__nfet_01v8_LHQHT5  amp_XM4_18
timestamp 1713225924
transform 1 0 17147 0 1 -5138
box -1083 -610 1083 610
use sky130_fd_pr__pfet_01v8_EDYT7U  amp_XM6
timestamp 1713225924
transform -1 0 19728 0 -1 -6597
box -996 -269 996 269
use sky130_fd_pr__nfet_01v8_UY343Z  amp_XM7
timestamp 1713225924
transform -1 0 19748 0 -1 -5584
box -996 -260 996 260
use sky130_fd_pr__pfet_01v8_EDYT7U  amp_XM8
timestamp 1713225924
transform 0 1 9847 -1 0 -8280
box -996 -269 996 269
use sky130_fd_pr__nfet_01v8_UY343Z  amp_XM9
timestamp 1713225924
transform 0 1 9258 -1 0 -8546
box -996 -260 996 260
use sky130_fd_pr__pfet_01v8_M6QFHF  amp_XM10_12
timestamp 1713225924
transform 1 0 21641 0 1 -6575
box -425 -383 425 383
use sky130_fd_pr__nfet_01v8_6G4XAN  amp_XM11_13
timestamp 1713225924
transform 1 0 21641 0 1 -5561
box -425 -365 425 365
use sky130_fd_pr__pfet_01v8_LL48TN  amp_XM16_17
timestamp 1713225924
transform 1 0 12884 0 1 -6453
box -2398 -683 2398 683
use sky130_fd_pr__res_xhigh_po_0p35_WHP78W  amp_XR1
timestamp 1713225924
transform 0 1 17636 -1 0 -8635
box -1363 -7182 1363 7182
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  ant_diode_ena
timestamp 1713225924
transform 1 0 2933 0 1 -997
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  ant_diode_standby
timestamp 1713225924
transform 1 0 5403 0 1 -997
box -183 -183 183 183
use sky130_fd_pr__cap_mim_m3_1_VMUSDZ  bias_XC1
timestamp 1713225924
transform 0 1 13498 -1 0 -21238
box -2386 -11680 2092 11684
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  bias_XC2
timestamp 1713362484
transform -1 0 3588 0 -1 -11370
box -2186 -2040 1882 2040
use sky130_fd_pr__cap_mim_m3_1_F5PPB9  bias_XC3
timestamp 1713225924
transform 0 -1 9528 1 0 -16620
box -1986 -7722 1700 7724
use sky130_fd_pr__nfet_g5v0d10v5_BKL7UB  bias_XM1_2
timestamp 1713225924
transform 0 1 20853 -1 0 -14102
box -1584 -1113 1584 1113
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  bias_XM5
timestamp 1713225924
transform 1 0 7426 0 1 -12350
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_H6M2KM  bias_XM6_7_8
timestamp 1713225924
transform -1 0 10726 0 -1 -12352
box -2686 -300 2686 300
use sky130_fd_pr__res_xhigh_po_0p35_M35ED8  bias_XR2
timestamp 1713225924
transform 0 1 10748 -1 0 -15970
box -2276 -8782 2276 8782
use sky130_fd_pr__res_xhigh_po_0p35_VTNT3C  bias_XR3
timestamp 1713225924
transform 0 1 11050 -1 0 -13206
box -450 -8082 450 8082
use sky130_fd_sc_hd__tapvpwrvgnd_1  ena_buf_tap $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712500979
transform 0 1 2950 -1 0 -1232
box -38 -48 130 592
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  esd_n_xin
timestamp 1713225924
transform 1 0 20505 0 1 -22985
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  esd_n_xout
timestamp 1713225924
transform 1 0 23613 0 1 -22987
box -183 -183 183 183
use sky130_fd_pr__diode_pd2nw_05v5_K4SERG  esd_p_xin
timestamp 1713225924
transform 1 0 21361 0 1 -22975
box -321 -321 321 321
use sky130_fd_pr__diode_pd2nw_05v5_K4SERG  esd_p_xout
timestamp 1713225924
transform 1 0 22787 0 1 -22977
box -321 -321 321 321
use sky130_fd_sc_hd__tapvpwrvgnd_1  standby_buf_tap
timestamp 1712500979
transform 0 -1 5380 1 0 -1324
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712500979
transform 0 1 2950 -1 0 -1324
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x2
timestamp 1712500979
transform 0 -1 5380 -1 0 -1324
box -38 -48 314 592
use level_shift  x3
timestamp 1713225924
transform 0 1 4250 -1 0 -1190
box 652 -1950 5670 -128
use level_shift  x4
timestamp 1713225924
transform 0 -1 4086 -1 0 -1190
box 652 -1950 5670 -128
use ripl_dly_clk_buf  x7
timestamp 1713360460
transform 1 0 13446 0 1 -1060
box 216 -2416 9016 -120
use sky130_fd_pr__cap_mim_m3_1_UYSCL3  XC1
timestamp 1713225924
transform 0 1 15424 -1 0 -12168
box -1892 -1614 1336 1624
use sky130_fd_pr__cap_mim_m3_1_43FTN9  XC2
timestamp 1713225924
transform 1 0 21888 0 1 -9798
box -3546 -8008 3672 8020
use sky130_fd_pr__cap_mim_m3_1_3DMTNZ  XC3
timestamp 1713225924
transform 1 0 4424 0 1 -6020
box -2492 -2268 1950 2222
use sky130_fd_pr__cap_mim_m3_1_4HHTN9  XC4
timestamp 1713225924
transform 0 -1 11504 1 0 -2544
box -1186 -4640 890 4640
use sky130_fd_pr__nfet_g5v0d10v5_YG6WAD  XM1
timestamp 1713225924
transform 0 1 20864 -1 0 -17009
box -1147 -658 1147 658
use sky130_fd_pr__pfet_g5v0d10v5_E4RF2H  XM2_bias_XM3_4
timestamp 1713225924
transform 0 1 23465 -1 0 -15266
box -2770 -1161 2770 1161
use sky130_fd_pr__nfet_01v8_AHZR5K  XM3
timestamp 1713225924
transform 0 1 12824 -1 0 -2652
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_HZ6WG7  XM4
timestamp 1713225924
transform 0 1 23509 -1 0 -5548
box -296 -285 296 285
use sky130_fd_pr__nfet_g5v0d10v5_GZN5JV  XM5
timestamp 1713225924
transform -1 0 2863 0 1 -7653
box -594 -658 594 658
use sky130_fd_pr__pfet_g5v0d10v5_74GBJT  XM6
timestamp 1713225924
transform 1 0 4238 0 -1 -7655
box -624 -697 624 697
use sky130_fd_pr__pfet_01v8_3H68VM  XM7
timestamp 1713225924
transform 0 -1 23531 1 0 -6550
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_MTZJAC  XM8
timestamp 1713225924
transform 1 0 8283 0 1 -2587
box -957 -619 957 619
use sky130_fd_pr__pfet_g5v0d10v5_6RLJVT  XM9
timestamp 1713225924
transform -1 0 11530 0 -1 -2569
box -308 -697 308 697
use sky130_fd_pr__nfet_01v8_Y7GPAW  XM11
timestamp 1713225924
transform 1 0 10209 0 1 -2592
box -957 -610 957 610
use sky130_fd_pr__res_xhigh_po_0p35_68VL2P  XR2
timestamp 1713225924
transform 0 1 13546 -1 0 -20477
box -2193 -11582 2193 11582
<< labels >>
flabel metal2 2178 -1212 2578 -812 0 FreeSans 1200 0 0 0 avdd
port 1 nsew
flabel metal2 1626 -1212 2026 -812 0 FreeSans 1200 0 0 0 avss
port 2 nsew
flabel metal2 8076 -1212 8476 -812 0 FreeSans 1200 0 0 0 dvdd
port 3 nsew
flabel metal2 9976 -1212 10376 -812 0 FreeSans 1200 0 0 0 dvss
port 4 nsew
flabel metal2 11192 -1212 11592 -812 0 FreeSans 1200 0 0 0 ibias
port 5 nsew
flabel metal2 3592 -1212 3992 -812 0 FreeSans 1200 0 0 0 ena
port 6 nsew
flabel metal2 4338 -1212 4738 -812 0 FreeSans 1200 0 0 0 standby
port 7 nsew
flabel metal2 23912 -1212 24312 -812 0 FreeSans 1200 0 0 0 dout
port 8 nsew
flabel metal1 23054 -23704 23454 -23304 0 FreeSans 1200 0 0 0 xout
port 9 nsew
flabel metal1 20656 -23704 21056 -23304 0 FreeSans 1200 0 0 0 xin
port 10 nsew
flabel metal1 19460 -14978 19640 -13228 0 FreeSans 400 0 0 0 vrb
flabel metal1 22240 -14982 22400 -14170 0 FreeSans 400 0 0 0 vg1
flabel metal1 22120 -11668 25450 -10450 0 FreeSans 3200 0 0 0 avdd_ip
flabel metal1 18284 -11798 21916 -11292 0 FreeSans 3200 0 0 0 avss_ip
flabel metal2 18932 -14146 19712 -13978 0 FreeSans 400 0 0 0 vg2
flabel metal1 21956 -15750 22156 -14384 0 FreeSans 400 0 0 0 vbreg
flabel metal2 7082 -11968 7984 -11778 0 FreeSans 800 0 0 0 icnode
flabel metal2 5592 -7636 9246 -7536 0 FreeSans 800 0 0 0 standby_33
flabel metal2 6632 -1444 7372 -1344 0 FreeSans 800 0 0 0 standby_ip
flabel metal2 6812 -1600 7378 -1500 0 FreeSans 800 0 0 0 ena_ip
flabel metal2 6974 -1784 7378 -1684 0 FreeSans 800 0 0 0 standby_b
flabel viali 8878 -7250 10492 -5640 0 FreeSans 3200 0 0 0 dvdd_ip
flabel viali 8900 -5476 10462 -4316 0 FreeSans 3200 0 0 0 dvss_ip
flabel metal2 13962 -4022 22308 -3882 0 FreeSans 800 0 0 0 dout_ip
flabel metal2 14360 -3780 22856 -3640 0 FreeSans 800 0 0 0 dout_filt
flabel metal2 11826 -4626 11926 -3164 0 FreeSans 800 0 0 0 ibias_ip
flabel metal2 12998 -5906 13098 -5346 0 FreeSans 800 0 0 0 vbp
flabel metal2 13948 -6502 17014 -6402 0 FreeSans 800 0 0 0 tail
flabel metal1 16648 -6108 16728 -5530 0 FreeSans 800 0 0 0 vn
flabel metal2 17500 -6100 17712 -5772 0 FreeSans 800 0 0 0 xin_buf
flabel metal2 19082 -6474 19242 -5706 0 FreeSans 800 0 0 0 inv_in
flabel metal2 20668 -6110 21562 -6010 0 FreeSans 800 0 0 0 inv_m1
flabel metal1 21718 -6828 21818 -5328 0 FreeSans 800 0 0 0 inv_m2
<< end >>
