magic
tech sky130A
magscale 1 2
timestamp 1712954147
<< pwell >>
rect -2276 -8782 2276 8782
<< psubdiff >>
rect -2240 8712 -2144 8746
rect 2144 8712 2240 8746
rect -2240 8650 -2206 8712
rect 2206 8650 2240 8712
rect -2240 -8712 -2206 -8650
rect 2206 -8712 2240 -8650
rect -2240 -8746 -2144 -8712
rect 2144 -8746 2240 -8712
<< psubdiffcont >>
rect -2144 8712 2144 8746
rect -2240 -8650 -2206 8650
rect 2206 -8650 2240 8650
rect -2144 -8746 2144 -8712
<< xpolycontact >>
rect -2110 8184 -2040 8616
rect -2110 -8616 -2040 -8184
rect -1944 8184 -1874 8616
rect -1944 -8616 -1874 -8184
rect -1778 8184 -1708 8616
rect -1778 -8616 -1708 -8184
rect -1612 8184 -1542 8616
rect -1612 -8616 -1542 -8184
rect -1446 8184 -1376 8616
rect -1446 -8616 -1376 -8184
rect -1280 8184 -1210 8616
rect -1280 -8616 -1210 -8184
rect -1114 8184 -1044 8616
rect -1114 -8616 -1044 -8184
rect -948 8184 -878 8616
rect -948 -8616 -878 -8184
rect -782 8184 -712 8616
rect -782 -8616 -712 -8184
rect -616 8184 -546 8616
rect -616 -8616 -546 -8184
rect -450 8184 -380 8616
rect -450 -8616 -380 -8184
rect -284 8184 -214 8616
rect -284 -8616 -214 -8184
rect -118 8184 -48 8616
rect -118 -8616 -48 -8184
rect 48 8184 118 8616
rect 48 -8616 118 -8184
rect 214 8184 284 8616
rect 214 -8616 284 -8184
rect 380 8184 450 8616
rect 380 -8616 450 -8184
rect 546 8184 616 8616
rect 546 -8616 616 -8184
rect 712 8184 782 8616
rect 712 -8616 782 -8184
rect 878 8184 948 8616
rect 878 -8616 948 -8184
rect 1044 8184 1114 8616
rect 1044 -8616 1114 -8184
rect 1210 8184 1280 8616
rect 1210 -8616 1280 -8184
rect 1376 8184 1446 8616
rect 1376 -8616 1446 -8184
rect 1542 8184 1612 8616
rect 1542 -8616 1612 -8184
rect 1708 8184 1778 8616
rect 1708 -8616 1778 -8184
rect 1874 8184 1944 8616
rect 1874 -8616 1944 -8184
rect 2040 8184 2110 8616
rect 2040 -8616 2110 -8184
<< xpolyres >>
rect -2110 -8184 -2040 8184
rect -1944 -8184 -1874 8184
rect -1778 -8184 -1708 8184
rect -1612 -8184 -1542 8184
rect -1446 -8184 -1376 8184
rect -1280 -8184 -1210 8184
rect -1114 -8184 -1044 8184
rect -948 -8184 -878 8184
rect -782 -8184 -712 8184
rect -616 -8184 -546 8184
rect -450 -8184 -380 8184
rect -284 -8184 -214 8184
rect -118 -8184 -48 8184
rect 48 -8184 118 8184
rect 214 -8184 284 8184
rect 380 -8184 450 8184
rect 546 -8184 616 8184
rect 712 -8184 782 8184
rect 878 -8184 948 8184
rect 1044 -8184 1114 8184
rect 1210 -8184 1280 8184
rect 1376 -8184 1446 8184
rect 1542 -8184 1612 8184
rect 1708 -8184 1778 8184
rect 1874 -8184 1944 8184
rect 2040 -8184 2110 8184
<< locali >>
rect -2240 8712 -2144 8746
rect 2144 8712 2240 8746
rect -2240 8650 -2206 8712
rect 2206 8650 2240 8712
rect -2240 -8712 -2206 -8650
rect 2206 -8712 2240 -8650
rect -2240 -8746 -2144 -8712
rect 2144 -8746 2240 -8712
<< viali >>
rect -2094 8201 -2056 8598
rect -1928 8201 -1890 8598
rect -1762 8201 -1724 8598
rect -1596 8201 -1558 8598
rect -1430 8201 -1392 8598
rect -1264 8201 -1226 8598
rect -1098 8201 -1060 8598
rect -932 8201 -894 8598
rect -766 8201 -728 8598
rect -600 8201 -562 8598
rect -434 8201 -396 8598
rect -268 8201 -230 8598
rect -102 8201 -64 8598
rect 64 8201 102 8598
rect 230 8201 268 8598
rect 396 8201 434 8598
rect 562 8201 600 8598
rect 728 8201 766 8598
rect 894 8201 932 8598
rect 1060 8201 1098 8598
rect 1226 8201 1264 8598
rect 1392 8201 1430 8598
rect 1558 8201 1596 8598
rect 1724 8201 1762 8598
rect 1890 8201 1928 8598
rect 2056 8201 2094 8598
rect -2094 -8598 -2056 -8201
rect -1928 -8598 -1890 -8201
rect -1762 -8598 -1724 -8201
rect -1596 -8598 -1558 -8201
rect -1430 -8598 -1392 -8201
rect -1264 -8598 -1226 -8201
rect -1098 -8598 -1060 -8201
rect -932 -8598 -894 -8201
rect -766 -8598 -728 -8201
rect -600 -8598 -562 -8201
rect -434 -8598 -396 -8201
rect -268 -8598 -230 -8201
rect -102 -8598 -64 -8201
rect 64 -8598 102 -8201
rect 230 -8598 268 -8201
rect 396 -8598 434 -8201
rect 562 -8598 600 -8201
rect 728 -8598 766 -8201
rect 894 -8598 932 -8201
rect 1060 -8598 1098 -8201
rect 1226 -8598 1264 -8201
rect 1392 -8598 1430 -8201
rect 1558 -8598 1596 -8201
rect 1724 -8598 1762 -8201
rect 1890 -8598 1928 -8201
rect 2056 -8598 2094 -8201
<< metal1 >>
rect -2100 8598 -2050 8610
rect -2100 8201 -2094 8598
rect -2056 8201 -2050 8598
rect -2100 8189 -2050 8201
rect -1934 8598 -1884 8610
rect -1934 8201 -1928 8598
rect -1890 8201 -1884 8598
rect -1934 8189 -1884 8201
rect -1768 8598 -1718 8610
rect -1768 8201 -1762 8598
rect -1724 8201 -1718 8598
rect -1768 8189 -1718 8201
rect -1602 8598 -1552 8610
rect -1602 8201 -1596 8598
rect -1558 8201 -1552 8598
rect -1602 8189 -1552 8201
rect -1436 8598 -1386 8610
rect -1436 8201 -1430 8598
rect -1392 8201 -1386 8598
rect -1436 8189 -1386 8201
rect -1270 8598 -1220 8610
rect -1270 8201 -1264 8598
rect -1226 8201 -1220 8598
rect -1270 8189 -1220 8201
rect -1104 8598 -1054 8610
rect -1104 8201 -1098 8598
rect -1060 8201 -1054 8598
rect -1104 8189 -1054 8201
rect -938 8598 -888 8610
rect -938 8201 -932 8598
rect -894 8201 -888 8598
rect -938 8189 -888 8201
rect -772 8598 -722 8610
rect -772 8201 -766 8598
rect -728 8201 -722 8598
rect -772 8189 -722 8201
rect -606 8598 -556 8610
rect -606 8201 -600 8598
rect -562 8201 -556 8598
rect -606 8189 -556 8201
rect -440 8598 -390 8610
rect -440 8201 -434 8598
rect -396 8201 -390 8598
rect -440 8189 -390 8201
rect -274 8598 -224 8610
rect -274 8201 -268 8598
rect -230 8201 -224 8598
rect -274 8189 -224 8201
rect -108 8598 -58 8610
rect -108 8201 -102 8598
rect -64 8201 -58 8598
rect -108 8189 -58 8201
rect 58 8598 108 8610
rect 58 8201 64 8598
rect 102 8201 108 8598
rect 58 8189 108 8201
rect 224 8598 274 8610
rect 224 8201 230 8598
rect 268 8201 274 8598
rect 224 8189 274 8201
rect 390 8598 440 8610
rect 390 8201 396 8598
rect 434 8201 440 8598
rect 390 8189 440 8201
rect 556 8598 606 8610
rect 556 8201 562 8598
rect 600 8201 606 8598
rect 556 8189 606 8201
rect 722 8598 772 8610
rect 722 8201 728 8598
rect 766 8201 772 8598
rect 722 8189 772 8201
rect 888 8598 938 8610
rect 888 8201 894 8598
rect 932 8201 938 8598
rect 888 8189 938 8201
rect 1054 8598 1104 8610
rect 1054 8201 1060 8598
rect 1098 8201 1104 8598
rect 1054 8189 1104 8201
rect 1220 8598 1270 8610
rect 1220 8201 1226 8598
rect 1264 8201 1270 8598
rect 1220 8189 1270 8201
rect 1386 8598 1436 8610
rect 1386 8201 1392 8598
rect 1430 8201 1436 8598
rect 1386 8189 1436 8201
rect 1552 8598 1602 8610
rect 1552 8201 1558 8598
rect 1596 8201 1602 8598
rect 1552 8189 1602 8201
rect 1718 8598 1768 8610
rect 1718 8201 1724 8598
rect 1762 8201 1768 8598
rect 1718 8189 1768 8201
rect 1884 8598 1934 8610
rect 1884 8201 1890 8598
rect 1928 8201 1934 8598
rect 1884 8189 1934 8201
rect 2050 8598 2100 8610
rect 2050 8201 2056 8598
rect 2094 8201 2100 8598
rect 2050 8189 2100 8201
rect -2100 -8201 -2050 -8189
rect -2100 -8598 -2094 -8201
rect -2056 -8598 -2050 -8201
rect -2100 -8610 -2050 -8598
rect -1934 -8201 -1884 -8189
rect -1934 -8598 -1928 -8201
rect -1890 -8598 -1884 -8201
rect -1934 -8610 -1884 -8598
rect -1768 -8201 -1718 -8189
rect -1768 -8598 -1762 -8201
rect -1724 -8598 -1718 -8201
rect -1768 -8610 -1718 -8598
rect -1602 -8201 -1552 -8189
rect -1602 -8598 -1596 -8201
rect -1558 -8598 -1552 -8201
rect -1602 -8610 -1552 -8598
rect -1436 -8201 -1386 -8189
rect -1436 -8598 -1430 -8201
rect -1392 -8598 -1386 -8201
rect -1436 -8610 -1386 -8598
rect -1270 -8201 -1220 -8189
rect -1270 -8598 -1264 -8201
rect -1226 -8598 -1220 -8201
rect -1270 -8610 -1220 -8598
rect -1104 -8201 -1054 -8189
rect -1104 -8598 -1098 -8201
rect -1060 -8598 -1054 -8201
rect -1104 -8610 -1054 -8598
rect -938 -8201 -888 -8189
rect -938 -8598 -932 -8201
rect -894 -8598 -888 -8201
rect -938 -8610 -888 -8598
rect -772 -8201 -722 -8189
rect -772 -8598 -766 -8201
rect -728 -8598 -722 -8201
rect -772 -8610 -722 -8598
rect -606 -8201 -556 -8189
rect -606 -8598 -600 -8201
rect -562 -8598 -556 -8201
rect -606 -8610 -556 -8598
rect -440 -8201 -390 -8189
rect -440 -8598 -434 -8201
rect -396 -8598 -390 -8201
rect -440 -8610 -390 -8598
rect -274 -8201 -224 -8189
rect -274 -8598 -268 -8201
rect -230 -8598 -224 -8201
rect -274 -8610 -224 -8598
rect -108 -8201 -58 -8189
rect -108 -8598 -102 -8201
rect -64 -8598 -58 -8201
rect -108 -8610 -58 -8598
rect 58 -8201 108 -8189
rect 58 -8598 64 -8201
rect 102 -8598 108 -8201
rect 58 -8610 108 -8598
rect 224 -8201 274 -8189
rect 224 -8598 230 -8201
rect 268 -8598 274 -8201
rect 224 -8610 274 -8598
rect 390 -8201 440 -8189
rect 390 -8598 396 -8201
rect 434 -8598 440 -8201
rect 390 -8610 440 -8598
rect 556 -8201 606 -8189
rect 556 -8598 562 -8201
rect 600 -8598 606 -8201
rect 556 -8610 606 -8598
rect 722 -8201 772 -8189
rect 722 -8598 728 -8201
rect 766 -8598 772 -8201
rect 722 -8610 772 -8598
rect 888 -8201 938 -8189
rect 888 -8598 894 -8201
rect 932 -8598 938 -8201
rect 888 -8610 938 -8598
rect 1054 -8201 1104 -8189
rect 1054 -8598 1060 -8201
rect 1098 -8598 1104 -8201
rect 1054 -8610 1104 -8598
rect 1220 -8201 1270 -8189
rect 1220 -8598 1226 -8201
rect 1264 -8598 1270 -8201
rect 1220 -8610 1270 -8598
rect 1386 -8201 1436 -8189
rect 1386 -8598 1392 -8201
rect 1430 -8598 1436 -8201
rect 1386 -8610 1436 -8598
rect 1552 -8201 1602 -8189
rect 1552 -8598 1558 -8201
rect 1596 -8598 1602 -8201
rect 1552 -8610 1602 -8598
rect 1718 -8201 1768 -8189
rect 1718 -8598 1724 -8201
rect 1762 -8598 1768 -8201
rect 1718 -8610 1768 -8598
rect 1884 -8201 1934 -8189
rect 1884 -8598 1890 -8201
rect 1928 -8598 1934 -8201
rect 1884 -8610 1934 -8598
rect 2050 -8201 2100 -8189
rect 2050 -8598 2056 -8201
rect 2094 -8598 2100 -8201
rect 2050 -8610 2100 -8598
<< properties >>
string FIXED_BBOX -2223 -8729 2223 8729
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 82 m 1 nx 26 wmin 0.350 lmin 0.50 rho 2000 val 469.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
