magic
tech sky130A
timestamp 1712087189
<< metal1 >>
rect 372 -278 472 -178
rect 122 -490 222 -390
rect 3653 -521 3753 -421
rect 369 -727 469 -627
rect 2053 -727 2153 -627
rect 3465 -727 3565 -627
use sky130_fd_sc_hd__and2_0  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 173 0 1 -589
box -19 -24 249 296
use sky130_fd_sc_hd__dfrbp_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 441 0 1 -589
box -19 -24 1077 296
use sky130_fd_sc_hd__dfrbp_1  x3
timestamp 1707688321
transform 1 0 1537 0 1 -589
box -19 -24 1077 296
use sky130_fd_sc_hd__dfrbp_1  x4
timestamp 1707688321
transform 1 0 2633 0 1 -589
box -19 -24 1077 296
<< labels >>
flabel metal1 3465 -727 3565 -627 0 FreeSans 64 0 0 0 done
port 3 nsew
flabel metal1 2053 -727 2153 -627 0 FreeSans 64 0 0 0 ena
port 5 nsew
flabel metal1 3653 -521 3753 -421 0 FreeSans 64 0 0 0 doneb
port 4 nsew
flabel metal1 122 -490 222 -390 0 FreeSans 64 0 0 0 clkin
port 2 nsew
flabel metal1 369 -727 469 -627 0 FreeSans 64 0 0 0 dvss
port 1 nsew
flabel metal1 372 -278 472 -178 0 FreeSans 64 0 0 0 dvdd
port 0 nsew
<< end >>
