* PEX produced on Sun Apr 14 23:49:44 EDT 2024 using /home/brady/sources/osic-multitool-src/iic-pex.sh with m=3 and s=1
* NGSPICE file created from sky130_be_ip__lsxo.ext - technology: sky130A

.subckt sky130_be_ip__lsxo dout ibias xin xout ena avss avdd standby dvss dvdd
X0 a_16620_n1869.t1 a_15705_n2241.t2 a_16273_n2273.t2 dvss.t210 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1 a_20376_n2791.t0 x7.x3.A2.t2 dvdd.t15 dvdd.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_21036_n1869.t0 a_19955_n2241.t2 a_20689_n2273.t0 dvdd.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3 a_10620_n8338.t0 a_24220_n8172.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X4 a_16795_n2817.t0 a_16620_n2791.t4 a_16974_n2791.t0 dvss.t289 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5 dvdd.t126 ena_ip.t2 x3.in_b.t0 dvdd.t125 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X6 dvdd.t159 a_21036_n1869.t4 a_21211_n1943.t0 dvdd.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_18828_n2791.t0 a_17913_n2791.t2 a_18481_n2549.t0 dvss.t118 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X8 a_2130_n19848.t0 a_24530_n20014.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X9 vbreg.t0 icnode.t2 a_11526_n12394.t1 dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X10 x7.x2.x2.CLK.t1 a_15000_n2791.t3 dvss.t57 dvss.t56 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X11 a_18168_n1881.t3 x7.x1.x4.CLK.t2 dvss.t274 dvss.t273 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X12 tail.t11 vbp.t3 dvdd_ip.t52 dvdd_ip.t42 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X13 a_16317_n2791.t1 a_16273_n2549.t4 a_16151_n2791.t1 dvss.t169 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X14 dvss.t250 x4.in_b.t0 dvss_ip dvss.t249 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X15 a_9120_n9346.t4 a_24220_n9832.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X16 a_16795_n1943.t1 a_16620_n1869.t4 a_16974_n1881.t0 dvss.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X17 x7.x3.B2.t0 a_21775_n2247.t2 dvdd.t17 dvdd.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X18 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X19 a_20121_n2241.t0 a_19955_n2241.t3 dvdd.t146 dvdd.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_2130_n21176.t1 a_24530_n21342.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X21 a_10658_n5446.t10 standby_33.t3 ibias.t1 ibias.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X22 xout.t20 vbreg.t9 avdd_ip.t28 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X23 inv_m1.t0 inv_in.t1 dvdd_ip.t7 dvdd_ip.t6 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X24 a_2132_n15590.t0 a_18932_n15756.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X25 dout_ip.t1 inv_m2.t2 dvdd_ip.t17 dvdd_ip.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X26 a_20733_n2791.t0 a_20689_n2549.t4 a_20567_n2791.t0 dvss.t5 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X27 inv_in.t2 a_17576_n6897.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X28 x7.x1.x2.CLK.t1 a_15000_n1881.t3 dvss.t108 dvss.t107 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X29 avdd_ip.t29 dvss sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X30 a_16317_n1881.t0 a_16273_n2273.t4 a_16151_n1869.t0 dvss.t65 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X31 x7.x3.A2.t0 a_21775_n2791.t2 dvss.t36 dvss.t35 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X32 a_14009_n2701.t1 x7.x5.TE_B.t2 dvss.t31 dvss.t30 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.07665 ps=0.785 w=0.42 l=0.15
X33 dvss.t29 standby_ip.t2 x4.in_b dvss.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X34 dvss.t63 a_2971_n1521.t2 ena_ip.t0 dvss.t62 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X35 dvss.t252 x4.in_b.t1 a_16317_n2791.t0 dvss.t251 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X36 avdd_ip.t30 dvss sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X37 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X38 dvss.t141 x7.x3.B2.t2 a_14035_n1997.t1 dvss.t98 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X39 x7.x3.A2.t1 a_21775_n2791.t3 dvdd.t117 dvdd.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X40 a_2132_n17582.t0 a_18932_n17416.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X41 inv_m1.t1 inv_in.t3 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X42 avss.t26 avdd.t11 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X43 a_10620_n9666.t0 a_24220_n9832.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X44 a_20733_n1881.t0 a_20689_n2273.t4 a_20567_n1869.t0 dvss.t41 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X45 dvdd.t29 x7.x2.x2.CLK.t2 a_15539_n2791.t0 dvdd.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X46 a_16782_n2425.t1 a_15705_n2791.t2 a_16620_n2791.t0 dvdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X47 dvdd_ip.t5 inv_m1.t2 inv_m2.t0 dvdd_ip.t4 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X48 a_4857_n1521.t0 standby.t0 dvdd.t33 dvdd.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X49 avdd_ip.t3 ena_b_33.t3 avdd.t14 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X50 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X51 a_20121_n2791.t1 a_19955_n2791.t2 dvss.t124 dvss.t123 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X52 dvss.t183 ena_ip.t3 a_16317_n1881.t1 dvss.t182 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X53 x7.x1.x4.CLK.t0 a_19567_n2247.t2 dvss.t219 dvss.t218 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X54 dvss.t93 ena.t0 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X55 dvdd.t88 a_19003_n2817.t3 a_19567_n2791.t0 dvdd.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X56 dvss vg1.t1 vg1.t2 dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X57 a_21145_n1869.t0 a_19955_n2241.t4 a_21036_n1869.t1 dvss.t170 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X58 avdd_ip.t21 vbreg.t10 avdd_ip.t20 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X59 a_21211_n2817.t2 x4.in_b.t2 dvdd.t31 dvdd.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X60 dvss xin.t6 dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=23.6118 ps=175.6 w=4 l=0.5
X61 a_19003_n2817.t1 a_18828_n2791.t4 a_19182_n2791.t0 dvss.t86 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X62 a_15000_n1881.t0 dout_ip.t5 dvdd.t53 dvdd.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
X63 a_2132_n17250.t0 a_18932_n17416.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X64 a_20121_n2241.t1 a_19955_n2241.t5 dvss.t172 dvss.t171 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X65 dvss_ip a_10658_n5446.t11 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=5.8 ps=45.8 w=2 l=2
X66 a_10620_n9666.t1 a_24220_n9500.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X67 a_18359_n1869.t0 a_17913_n2241.t2 a_18263_n1869.t2 dvss.t119 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X68 xout.t19 vbreg.t11 avdd_ip.t27 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X69 dvss dvss dvss sky130_fd_pr__res_xhigh_po_0p35 l=75
X70 vbreg.t2 vg2.t5 vrb.t4 dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X71 dvss ena_33.t3 avss.t7 avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X72 a_18525_n2791.t0 a_18481_n2549.t4 a_18359_n2791.t1 dvss.t148 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X73 a_2130_n20844.t1 a_24530_n21010.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X74 a_15083_n2791.t1 dout_ip.t6 a_15000_n2791.t1 dvss.t87 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X75 a_21036_n1869.t2 a_20121_n2241.t2 a_20689_n2273.t2 dvss.t227 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X76 dvss_ip x4.in_b.t3 dvss.t61 dvss.t60 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X77 a_2132_n15590.t1 a_18932_n15424.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X78 a_14285_n2079.t2 x7.x3.B2.t3 a_14285_n2281.t2 dvdd.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X79 a_19003_n1943.t1 a_18828_n1869.t4 a_19182_n1881.t0 dvss.t23 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X80 vn.t1 xin.t7 vn.t0 dvdd_ip.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X81 avss.t25 x4.in_b.t4 standby_33.t2 avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X82 a_10620_n7674.t1 a_24220_n7840.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X83 a_10658_n5446.t9 a_10658_n5446.t8 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X84 avdd.t3 ena_b_33.t4 avdd_ip.t0 avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X85 a_15960_n2791.t2 x7.x2.x3.CLK.t2 dvdd.t124 dvdd.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X86 a_2130_n19516.t1 a_24530_n19682.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X87 xin.t8 avdd_ip.t2 sky130_fd_pr__diode_pd2nw_05v5 perim=1.8e+06 area=2.025e+11
X88 a_20579_n2247.t2 ena_ip.t4 dvdd.t135 dvdd.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X89 dvdd.t42 a_2971_n1521.t3 ena_ip.t1 dvdd.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X90 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X91 a_15083_n1881.t0 dout_ip.t7 a_15000_n1881.t1 dvss.t88 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X92 a_18525_n1881.t0 a_18481_n2273.t4 a_18359_n1869.t1 dvss.t140 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X93 a_18168_n2791.t1 x7.x2.x4.CLK.t2 dvdd.t160 dvdd.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X94 dvss.t115 x4.in_b.t5 a_18525_n2791.t1 dvss.t114 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X95 a_17576_n6897.t4 xout.t23 tail.t0 dvdd_ip.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X96 a_16273_n2549.t2 a_16055_n2791.t4 dvdd.t122 dvdd.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X97 dvss.t135 x7.x3.A2.t3 a_15083_n2791.t0 dvss.t134 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X98 xout.t0 xin.t9 dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X99 x7.x1.x4.Q.t1 a_21211_n1943.t3 dvss.t224 dvss.t223 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X100 dvdd.t13 x7.x3.A2.t4 a_15000_n2791.t0 dvdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X101 a_14009_n2404.t0 standby_ip.t3 a_14285_n2079.t0 dvdd.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X102 dvss_ip x4.in_b.t6 dvss.t151 dvss.t150 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X103 avdd_ip.t23 vbreg.t12 xout.t18 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X104 tail.t10 vbp.t4 dvdd_ip.t51 dvdd_ip.t34 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X105 a_2130_n20844.t0 a_24530_n20678.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X106 a_16729_n1869.t1 a_15539_n2241.t2 a_16620_n1869.t3 dvss.t272 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X107 dvss vg2.t4 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X108 dvdd_ip.t50 vbp.t5 dvdd_ip.t49 dvdd_ip.t29 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X109 a_16273_n2273.t3 a_16055_n1869.t4 dvdd.t170 dvdd.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X110 a_2132_n15258.t1 a_18932_n15424.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X111 a_18990_n2425.t0 a_17913_n2791.t3 a_18828_n2791.t1 dvdd.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X112 a_14285_n2281.t0 x7.x3.A2.t5 dvdd.t11 dvdd.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X113 avdd_ip.t26 vbreg.t13 avdd_ip.t25 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X114 dvss.t191 ena_ip.t5 a_18525_n1881.t1 dvss.t190 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X115 dvdd.t151 a_21211_n1943.t4 a_21775_n2247.t0 dvdd.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X116 dvss.t246 x7.x3.B2.t4 a_15083_n1881.t1 dvss.t245 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X117 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X118 a_16795_n1943.t2 ena_ip.t6 dvdd.t90 dvdd.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X119 dvss.t0 standby.t1 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X120 dvss.t153 x4.in_b.t7 dvss_ip dvss.t152 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X121 a_2130_n19516.t0 a_24530_n19350.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X122 dvdd.t131 a_14009_n2404.t4 x7.x5.TE_B.t0 dvdd.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X123 dvss dvss dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X124 dvdd_ip.t54 standby_ip.t4 dvdd.t165 dvdd.t164 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X125 a_16163_n2247.t2 ena_ip.t7 dvdd.t92 dvdd.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X126 a_2132_n16918.t1 a_18932_n17084.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X127 dvdd.t120 x7.x2.x4.CLK.t3 a_19955_n2791.t1 dvdd.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X128 a_19003_n1943.t2 ena_ip.t8 dvdd.t150 dvdd.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X129 inv_in.t4 a_17576_n6897.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X130 a_10620_n9334.t1 a_24220_n9500.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X131 dvss.t69 a_21211_n2817.t3 a_21775_n2791.t0 dvss.t68 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X132 a_3134_n13324.t0 vrb.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=75
X133 dvdd_ip.t55 standby_ip.t5 dvdd.t167 dvdd.t166 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X134 a_16974_n2791.t1 x4.in_b.t8 dvss.t145 dvss.t144 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X135 x7.x1.x2.Q.t1 a_16795_n1943.t3 dvss.t49 dvss.t48 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X136 a_2132_n17582.t1 a_18932_n17748.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X137 dvdd.t127 x7.x1.x2.CLK.t2 a_15539_n2241.t0 dvdd.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X138 dvdd_ip.t48 vbp.t6 tail.t9 dvdd_ip.t27 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X139 a_19182_n2791.t1 x4.in_b.t9 dvss.t147 dvss.t146 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X140 dvss.t139 a_19003_n2817.t4 a_18937_n2791.t0 dvss.t138 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X141 dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X142 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X143 dout_ip.t3 inv_m2.t3 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X144 a_15705_n2791.t0 a_15539_n2791.t2 dvdd.t25 dvdd.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X145 avdd.t5 ena_b_33.t5 ena_33.t2 avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X146 dvdd.t59 a_16795_n2817.t3 a_16782_n2425.t0 dvdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X147 dvss.t229 a_21211_n1943.t5 a_21775_n2247.t1 dvss.t228 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X148 xout.t2 xin.t10 dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X149 dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X150 a_16974_n1881.t1 ena_ip.t9 dvss.t221 dvss.t220 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X151 dvdd.t27 a_16795_n1943.t4 a_17359_n2247.t0 dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X152 xin.t0 a_24530_n22338.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X153 dvss.t33 x7.x5.TE_B.t3 dout_filt.t2 dvss.t32 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X154 a_16055_n2791.t2 a_15539_n2791.t3 a_15960_n2791.t1 dvss.t163 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X155 dvdd.t23 standby_ip.t6 dvdd_ip.t8 dvdd.t22 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X156 standby_33.t0 x4.out_b.t3 avdd.t1 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X157 a_16055_n1869.t2 a_15705_n2241.t3 a_15960_n1881.t2 dvdd.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X158 dvdd_ip.t47 vbp.t7 tail.t8 dvdd_ip.t40 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X159 a_20471_n2791.t0 a_20121_n2791.t2 a_20376_n2791.t2 dvdd.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X160 dvss xout.t24 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X161 tail.t7 vbp.t8 dvdd_ip.t46 dvdd_ip.t38 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X162 dvdd.t87 a_19003_n2817.t5 a_18990_n2425.t1 dvdd.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X163 a_10620_n9334.t0 a_24220_n9168.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X164 a_19182_n1881.t1 ena_ip.t10 dvss.t216 dvss.t215 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X165 avdd_ip.t24 vbreg.t14 xout.t17 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X166 dvss xin.t11 xout.t10 dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X167 a_17576_n6897.t3 xout.t25 a_17576_n6897.t3 dvdd_ip.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0 ps=0 w=4 l=2
X168 a_3134_n13324.t1 dvss dvss sky130_fd_pr__res_xhigh_po_0p35 l=75
X169 a_21036_n2791.t2 a_19955_n2791.t3 a_20689_n2549.t3 dvdd.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X170 dvss.t178 a_19003_n1943.t3 a_18937_n1869.t0 dvss.t177 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X171 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X172 a_18937_n2791.t1 a_17747_n2791.t2 a_18828_n2791.t3 dvss.t255 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X173 dvss.t113 a_16795_n2817.t4 a_17359_n2791.t1 dvss.t112 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X174 a_16273_n2273.t0 a_16055_n1869.t5 dvss.t189 dvss.t188 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X175 dvdd.t9 a_16620_n1869.t5 a_16795_n1943.t0 dvdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X176 x7.x1.x2.Q.t0 a_16795_n1943.t5 dvdd.t102 dvdd.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X177 a_2130_n20512.t0 a_24530_n20678.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X178 dvss xin.t12 xout.t8 dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X179 dvdd.t51 a_21036_n2791.t4 a_21211_n2817.t1 dvdd.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X180 x4.out_b.t2 standby_ip.t7 avss.t13 avss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X181 a_18481_n2549.t2 a_18263_n2791.t4 dvdd.t80 dvdd.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X182 dvss_ip inv_m1.t3 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=7.9025 ps=61.46 w=0.5 l=1
X183 a_10658_n5446.t7 a_10658_n5446.t6 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X184 dvss.t59 x7.x2.x2.CLK.t3 a_15539_n2791.t1 dvss.t58 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X185 xout.t7 xin.t13 dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X186 a_2132_n14926.t1 a_18932_n15092.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X187 dvdd.t38 x7.x5.TE_B.t4 a_14357_n2743.t1 dvdd.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.005 as=0.0672 ps=0.85 w=0.64 l=0.15
X188 vn.t7 vn.t5 vn.t6 dvss_ip sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X189 a_20567_n2791.t1 a_20121_n2791.t3 a_20471_n2791.t1 dvss.t217 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X190 dvdd.t76 standby_ip.t8 dvdd_ip.t15 dvdd.t75 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X191 dvss_ip dout_filt.t3 dout.t1 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=1
X192 a_20471_n1869.t0 a_19955_n2241.t6 a_20376_n1881.t0 dvss.t149 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X193 a_18481_n2273.t1 a_18263_n1869.t4 dvdd.t107 dvdd.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X194 dvss.t143 a_16795_n1943.t6 a_17359_n2247.t1 dvss.t142 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X195 x7.x1.x3.CLK.t0 a_17359_n2247.t2 dvdd.t5 dvdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X196 dvdd_ip.t45 vbp.t9 tail.t6 dvdd_ip.t36 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X197 avss.t27 avdd.t10 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X198 x7.x2.x2.Q.t0 a_16795_n2817.t5 dvdd.t140 dvdd.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X199 a_14035_n2743.t0 dout_ip.t8 dout_filt.t1 dvss.t30 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X200 dvss.t185 x7.x1.x2.CLK.t3 a_15539_n2241.t1 dvss.t184 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X201 dout_ip.t2 inv_m2.t4 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X202 a_17576_n6897.t2 vn.t8 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X203 avdd_ip.t22 vbreg.t15 vg1.t3 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X204 a_2130_n19848.t1 a_24530_n19682.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X205 vrb.t3 vg2.t6 vbreg.t1 dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X206 a_18828_n1869.t1 a_17913_n2241.t3 a_18481_n2273.t0 dvss.t125 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X207 x7.x2.x3.CLK.t1 a_17359_n2791.t2 dvss.t83 dvss.t82 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X208 a_2130_n20512.t1 a_24530_n20346.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X209 dvdd.t174 a_20689_n2273.t5 a_20579_n2247.t0 dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X210 x7.x1.x2.CLK.t0 a_15000_n1881.t4 dvdd.t83 dvdd.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X211 dvdd_ip.t16 standby_ip.t9 dvdd.t78 dvdd.t77 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X212 a_2132_n14926.t0 a_18932_n14760.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X213 x7.x2.x3.CLK.t0 a_17359_n2791.t3 dvdd.t35 dvdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X214 x7.x1.x3.Q.t1 a_19003_n1943.t4 dvss.t103 dvss.t102 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X215 xout.t4 xin.t14 dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X216 avdd.t16 ena_b_33.t6 avdd_ip.t5 avdd.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X217 a_16273_n2549.t0 a_16055_n2791.t5 dvss.t67 dvss.t66 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X218 a_16151_n2791.t0 a_15705_n2791.t3 a_16055_n2791.t1 dvss.t45 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X219 vg1.t4 xin.t5 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X220 dvss xin.t15 xout.t6 dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X221 dvss_ip inv_m1.t4 inv_m2.t1 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X222 a_2130_n19184.t1 a_24530_n19018.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X223 dvdd_ip.t44 vbp.t10 dvdd_ip.t43 dvdd_ip.t42 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X224 inv_in.t5 a_17576_n6897.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X225 dvdd.t138 a_4857_n1521.t2 standby_ip.t1 dvdd.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X226 a_14035_n1997.t0 ena_ip.t11 a_14009_n2404.t2 dvss.t98 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X227 a_17913_n2791.t0 a_17747_n2791.t3 dvdd.t21 dvdd.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X228 a_4857_n1521.t1 standby.t2 dvss.t2 dvss.t1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X229 a_10620_n9002.t0 a_24220_n9168.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X230 a_18263_n2791.t2 a_17747_n2791.t4 a_18168_n2791.t3 dvss.t179 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X231 a_14009_n2404.t3 x4.in_b.t10 a_14035_n2281.t1 dvss.t98 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X232 a_16620_n1869.t0 a_15539_n2241.t3 a_16273_n2273.t1 dvdd.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X233 a_18263_n1869.t1 a_17913_n2241.t4 a_18168_n1881.t0 dvdd.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X234 a_10620_n9002.t1 a_24220_n8836.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X235 dvdd.t169 x7.x1.x4.CLK.t3 a_19955_n2241.t1 dvdd.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X236 a_2130_n20180.t1 a_24530_n20346.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X237 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X238 ena_b_33.t2 ena_33.t4 avdd.t19 avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X239 xout.t3 xin.t16 dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X240 avdd.t12 standby_33.t4 x4.out_b.t0 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X241 a_20579_n2247.t1 a_19955_n2241.t7 a_20471_n1869.t1 dvdd.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X242 dvdd.t44 a_16273_n2273.t5 a_16163_n2247.t1 dvdd.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X243 a_15000_n2791.t2 dout_ip.t9 dvdd.t118 dvdd.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
X244 dvdd.t156 a_18828_n1869.t5 a_19003_n1943.t0 dvdd.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X245 a_2130_n22172.t0 a_24530_n22006.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X246 dvss xin.t17 xout.t9 dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X247 avdd_ip.t31 dvss sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X248 a_15705_n2241.t0 a_15539_n2241.t4 dvdd.t155 dvdd.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X249 a_2130_n21840.t1 a_24530_n22006.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X250 avdd_ip.t19 vbreg.t16 xout.t16 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X251 dvdd.t47 x7.x2.x3.CLK.t3 a_17747_n2791.t0 dvdd.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X252 a_2132_n16586.t0 a_18932_n16420.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X253 dvss xin.t18 dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X254 a_10620_n8670.t1 a_24220_n8836.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X255 a_17576_n6897.t1 vn.t9 a_17576_n6897.t1 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0 ps=0 w=4 l=2
X256 x7.x1.x4.CLK.t1 a_19567_n2247.t3 dvdd.t149 dvdd.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X257 a_2132_n17250.t1 a_18932_n17084.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X258 a_14009_n2701.t0 x7.x5.TE_B.t5 dvdd.t40 dvdd.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.10855 ps=1.005 w=0.42 l=0.15
X259 dvss.t25 x7.x2.x4.CLK.t4 a_19955_n2791.t0 dvss.t24 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X260 dvss.t257 standby_ip.t10 dout_ip.t4 dvss.t256 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X261 dvss_ip a_10658_n5446.t12 vbp.t0 dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X262 inv_in.t6 a_17576_n6897.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X263 a_22601_n15524.t1 vbreg.t17 a_22601_n15524.t0 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X264 a_20579_n2425.t2 x4.in_b.t11 dvdd.t139 dvdd.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X265 a_16163_n2247.t0 a_15539_n2241.t5 a_16055_n1869.t0 dvdd.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X266 dvss xin.t19 xout.t5 dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X267 x7.x2.x4.CLK.t1 a_19567_n2791.t2 dvss.t55 dvss.t54 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X268 vbreg.t5 vg1.t5 vbreg.t4 dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X269 dvss ena_33.t5 avss.t21 avss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X270 vg1.t6 xin.t4 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X271 x3.in_b.t1 ena_ip.t12 dvss.t176 dvss.t175 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X272 x7.x2.x4.CLK.t0 a_19567_n2791.t3 dvdd.t109 dvdd.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X273 dvss.t92 x7.x1.x4.CLK.t4 a_19955_n2241.t0 dvss.t91 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X274 a_15705_n2791.t1 a_15539_n2791.t4 dvss.t165 dvss.t164 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X275 standby_33.t1 x4.in_b.t12 avss.t23 avss.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X276 vbreg.t8 vg2.t7 vrb.t2 dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X277 tail.t1 xin.t20 vn.t2 dvdd_ip.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X278 dout_ip.t0 inv_m2.t5 dvdd_ip.t3 dvdd_ip.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X279 dvdd.t175 dvss.t180 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X280 avss.t5 ena_33.t6 dvss avss.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X281 dvdd.t55 a_21211_n1943.t6 a_21198_n2247.t1 dvdd.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X282 a_2130_n20180.t0 a_24530_n20014.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X283 dvdd_ip.t33 vbp.t11 dvdd_ip.t32 dvdd_ip.t24 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X284 a_20376_n2791.t1 x7.x3.A2.t6 dvss.t167 dvss.t166 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X285 a_18828_n1869.t2 a_17747_n2241.t2 a_18481_n2273.t3 dvdd.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X286 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X287 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X288 a_16795_n2817.t2 x4.in_b.t13 dvdd.t66 dvdd.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X289 a_2132_n14594.t0 a_18932_n14428.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X290 a_15705_n2241.t1 a_15539_n2241.t6 dvss.t269 dvss.t268 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X291 ena_33.t1 x3.in_b.t2 avss.t3 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X292 a_16163_n2425.t2 x4.in_b.t14 dvdd.t93 dvdd.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X293 inv_in.t7 a_17576_n6897.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X294 a_2132_n15258.t0 a_18932_n15092.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X295 a_19003_n2817.t2 x4.in_b.t15 dvdd.t95 dvdd.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X296 dvdd.t168 a_18481_n2273.t5 a_18371_n2247.t0 dvdd.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X297 dvss dvss dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X298 a_20376_n1881.t3 x7.x3.B2.t5 dvss.t248 dvss.t247 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X299 dvdd_ip.t13 inv_m1.t5 dvdd_ip.t12 dvdd_ip.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=1
X300 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X301 dvss.t195 x4.in_b.t16 dvss_ip dvss.t194 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X302 vg1.t7 xin.t3 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X303 a_2130_n19184.t0 a_24530_n19350.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X304 a_10620_n8670.t0 a_24220_n8504.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X305 a_17913_n2241.t0 a_17747_n2241.t3 dvdd.t129 dvdd.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X306 x7.x2.x4.Q.t1 a_21211_n2817.t4 dvss.t226 dvss.t225 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X307 dvss_ip a_10658_n5446.t4 a_10658_n5446.t5 dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X308 a_21198_n2247.t0 a_20121_n2241.t3 a_21036_n1869.t3 dvdd.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X309 a_20689_n2273.t3 a_20471_n1869.t4 dvss.t263 dvss.t262 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X310 x7.x1.x4.Q.t0 a_21211_n1943.t7 dvdd.t57 dvdd.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X311 xout.t22 vbreg.t18 xout.t21 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X312 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X313 a_2132_n16918.t0 a_18932_n16752.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X314 dvss vg2.t3 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X315 a_16055_n2791.t0 a_15705_n2791.t4 a_15960_n2791.t0 dvdd.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X316 dvss dvss dvss sky130_fd_pr__res_xhigh_po_0p35 l=75
X317 avss.t1 x3.in_b.t3 ena_33.t0 avss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X318 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X319 dvss_ip x4.in_b.t17 dvss.t197 dvss.t196 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X320 a_18371_n2247.t1 ena_ip.t13 dvdd.t112 dvdd.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X321 a_2130_n21508.t1 a_24530_n21674.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X322 a_18371_n2247.t2 a_17747_n2241.t4 a_18263_n1869.t3 dvdd.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X323 vbreg.t7 vbreg.t6 avdd_ip.t18 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X324 a_16620_n2791.t3 a_15705_n2791.t5 a_16273_n2549.t3 dvss.t198 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X325 x7.x2.x4.Q.t0 a_21211_n2817.t5 dvdd.t154 dvdd.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X326 dvdd.t173 a_16620_n2791.t5 a_16795_n2817.t1 dvdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X327 dvss_ip x4.in_b.t18 dvss.t203 dvss.t202 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X328 a_2130_n22172.t1 a_24530_n22338.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X329 a_10620_n8338.t1 a_24220_n8504.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X330 dvdd.t81 x7.x1.x3.CLK.t2 a_17747_n2241.t0 dvdd.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X331 dvdd.t162 standby_ip.t11 dvdd_ip.t53 dvdd.t161 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X332 inv_in.t8 a_17576_n6897.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X333 a_2132_n16586.t1 a_18932_n16752.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X334 a_17913_n2791.t1 a_17747_n2791.t5 dvss.t81 dvss.t80 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X335 a_16055_n1869.t1 a_15539_n2241.t7 a_15960_n1881.t0 dvss.t238 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X336 x7.x2.x2.Q.t1 a_16795_n2817.t6 dvss.t207 dvss.t206 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X337 avdd_ip.t32 dvss sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X338 x7.x3.B2.t1 a_21775_n2247.t3 dvss.t47 dvss.t46 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X339 dvss vg2.t2 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X340 dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X341 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X342 a_20689_n2549.t1 a_20471_n2791.t4 dvss.t7 dvss.t6 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X343 dvss.t205 x4.in_b.t19 dvss_ip dvss.t204 sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X344 dvdd.t49 a_19003_n1943.t5 a_19567_n2247.t0 dvdd.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X345 dvdd_ip.t21 a_9120_n9346.t0 a_9120_n9346.t1 dvdd_ip.t20 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X346 dvdd.t133 a_21211_n2817.t6 a_21775_n2791.t1 dvdd.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X347 a_20376_n1881.t2 x7.x3.B2.t6 dvdd.t99 dvdd.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X348 a_18937_n1869.t1 a_17747_n2241.t5 a_18828_n1869.t3 dvss.t239 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X349 dvss xin.t21 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X350 dvdd_ip.t41 vbp.t12 tail.t5 dvdd_ip.t40 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X351 a_21211_n2817.t0 a_21036_n2791.t5 a_21390_n2791.t1 dvss.t11 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X352 tail.t4 vbp.t13 dvdd_ip.t39 dvdd_ip.t38 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X353 a_17913_n2241.t1 a_17747_n2241.t6 dvss.t244 dvss.t243 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X354 dvdd.t1 a_20689_n2549.t5 a_20579_n2425.t0 dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X355 dvdd_ip.t18 standby_ip.t12 dvdd.t97 dvdd.t96 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X356 a_20567_n1869.t1 a_20121_n2241.t4 a_20471_n1869.t3 dvss.t155 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X357 dvdd.t176 dvss.t181 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X358 dvss.t267 a_19003_n2817.t6 a_19567_n2791.t1 dvss.t266 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X359 a_18481_n2273.t2 a_18263_n1869.t5 dvss.t193 dvss.t192 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X360 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X361 dvss_ip vn.t3 vn.t4 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X362 a_2130_n18852.t1 a_24530_n19018.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X363 dvss.t235 x7.x2.x3.CLK.t4 a_17747_n2791.t1 dvss.t234 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X364 dvdd.t177 dvss.t72 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X365 avss.t28 avdd.t9 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X366 avss.t11 standby_ip.t13 x4.out_b.t1 avss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X367 icnode.t1 vg2.t8 dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X368 avdd_ip.t17 vbreg.t19 xout.t15 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X369 a_21211_n1943.t1 a_21036_n1869.t5 a_21390_n1881.t0 dvss.t38 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X370 a_15960_n2791.t3 x7.x2.x3.CLK.t5 dvss.t133 dvss.t132 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X371 a_11526_n12394.t0 icnode.t3 a_8268_n12482.t0 dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X372 dvss dvss dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X373 dvss.t271 a_19003_n1943.t6 a_19567_n2247.t1 dvss.t270 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X374 xout.t14 vbreg.t20 avdd_ip.t16 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X375 dvss.t156 a_4857_n1521.t3 standby_ip.t0 dvss.t1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X376 a_14009_n2404.t1 standby_ip.t14 dvss.t99 dvss.t98 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X377 inv_in.t9 a_17576_n6897.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X378 dvdd_ip.t37 vbp.t1 vbp.t2 dvdd_ip.t36 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X379 a_2132_n14594.t1 a_18932_n14760.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X380 a_16620_n2791.t2 a_15539_n2791.t5 a_16273_n2549.t1 dvdd.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X381 dvss.t261 x7.x1.x3.CLK.t3 a_17747_n2241.t1 dvss.t260 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X382 a_18263_n2791.t0 a_17913_n2791.t4 a_18168_n2791.t0 dvdd.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X383 dvdd.t3 a_16795_n2817.t7 a_17359_n2791.t0 dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X384 a_2971_n1521.t0 ena.t1 dvss.t95 dvss.t94 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X385 dvss.t51 x4.in_b.t20 a_20733_n2791.t1 dvss.t50 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X386 a_15960_n1881.t1 x7.x1.x3.CLK.t4 dvss.t85 dvss.t84 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X387 a_14035_n2281.t0 x7.x3.A2.t7 dvss.t168 dvss.t98 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X388 a_20579_n2425.t1 a_19955_n2791.t4 a_20471_n2791.t2 dvdd.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X389 a_21145_n2791.t1 a_19955_n2791.t5 a_21036_n2791.t3 dvss.t275 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X390 dvdd.t67 a_16273_n2549.t5 a_16163_n2425.t1 dvdd.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X391 a_16151_n1869.t1 a_15705_n2241.t4 a_16055_n1869.t3 dvss.t209 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X392 a_2130_n18852.t0 xout.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X393 dvdd.t64 a_18828_n2791.t5 a_19003_n2817.t0 dvdd.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X394 a_16782_n2247.t1 a_15705_n2241.t5 a_16620_n1869.t2 dvdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X395 ena_b_33.t1 ena_ip.t14 avss.t19 avss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X396 dvss.t214 a_14009_n2404.t5 x7.x5.TE_B.t1 dvss.t98 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X397 avss.t29 avdd.t8 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X398 dvdd.t71 standby_ip.t15 dvdd_ip.t11 dvdd.t70 sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X399 a_18481_n2549.t3 a_18263_n2791.t5 dvss.t259 dvss.t258 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X400 a_18359_n2791.t0 a_17913_n2791.t5 a_18263_n2791.t1 dvss.t208 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X401 avdd_ip.t6 ena_b_33.t7 avdd.t18 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X402 a_18263_n1869.t0 a_17747_n2241.t7 a_18168_n1881.t1 dvss.t34 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X403 dvss.t174 ena_ip.t15 a_20733_n1881.t1 dvss.t173 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X404 x7.x2.x3.Q.t1 a_19003_n2817.t7 dvss.t101 dvss.t100 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X405 xout.t13 vbreg.t21 avdd_ip.t15 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X406 dvss dvss dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X407 x7.x1.x3.Q.t0 a_19003_n1943.t7 dvdd.t171 dvdd.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X408 a_21036_n2791.t0 a_20121_n2791.t4 a_20689_n2549.t2 dvss.t162 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X409 dvss.t53 x4.in_b.t21 dvss_ip dvss.t52 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X410 avdd_ip.t33 icnode.t0 sky130_fd_pr__cap_mim_m3_1 l=20 w=20
X411 a_21211_n1943.t2 ena_ip.t16 dvdd.t110 dvdd.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X412 inv_in.t10 a_17576_n6897.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X413 inv_in.t11 a_17576_n6897.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X414 a_10620_n8006.t0 a_24220_n8172.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X415 avdd_ip.t14 vbreg.t22 xout.t12 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X416 a_2130_n21840.t0 a_24530_n21674.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X417 inv_in.t12 a_17576_n6897.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X418 a_10620_n8006.t1 a_24220_n7840.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X419 avdd.t7 ena_b_33.t8 avdd_ip.t1 avdd.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X420 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X421 avss.t17 ena_ip.t17 ena_b_33.t0 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X422 a_2132_n16254.t0 a_18932_n16420.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X423 a_16163_n2425.t0 a_15539_n2791.t6 a_16055_n2791.t3 dvdd.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X424 tail.t3 vbp.t14 dvdd_ip.t35 dvdd_ip.t34 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X425 a_8268_n12482.t0 a_8268_n12482.t1 dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X426 x7.x2.x3.Q.t0 a_19003_n2817.t8 dvdd.t85 dvdd.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X427 dvss.t42 a_14009_n2701.t2 a_14035_n2743.t1 dvss.t30 sky130_fd_pr__nfet_01v8 ad=0.07665 pd=0.785 as=0.0441 ps=0.63 w=0.42 l=0.15
X428 x7.x2.x2.CLK.t0 a_15000_n2791.t4 dvdd.t152 dvdd.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X429 dvdd_ip.t31 vbp.t15 dvdd_ip.t30 dvdd_ip.t29 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X430 a_21390_n2791.t0 x4.in_b.t22 dvss.t15 dvss.t14 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X431 dvss.t212 a_21211_n2817.t7 a_21145_n2791.t0 dvss.t211 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X432 vg1.t8 xin.t2 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X433 dvss_ip x4.in_b.t23 dvss.t17 dvss.t16 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X434 inv_in.t13 a_17576_n6897.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X435 a_16729_n2791.t1 a_15539_n2791.t7 a_16620_n2791.t1 dvss.t64 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X436 a_9120_n9346.t3 a_9120_n9346.t2 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X437 a_2130_n21176.t0 a_24530_n21010.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X438 a_2132_n17914.t1 vg1.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X439 a_15960_n1881.t3 x7.x1.x3.CLK.t5 dvdd.t163 dvdd.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X440 a_20121_n2791.t0 a_19955_n2791.t6 dvdd.t172 dvdd.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X441 dvdd.t157 a_21211_n2817.t8 a_21198_n2425.t1 dvdd.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X442 a_14357_n2743.t0 dout_ip.t10 dout_filt.t0 dvdd.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X443 a_2971_n1521.t1 ena.t2 dvdd.t148 dvdd.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X444 a_21390_n1881.t1 ena_ip.t18 dvss.t237 dvss.t236 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X445 x4.in_b standby_ip.t16 dvdd.t114 dvdd.t113 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X446 dvss_ip a_10658_n5446.t2 a_10658_n5446.t3 dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X447 a_18828_n2791.t2 a_17747_n2791.t6 a_18481_n2549.t1 dvdd.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X448 a_18168_n1881.t2 x7.x1.x4.CLK.t5 dvdd.t69 dvdd.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X449 dvdd.t178 dvss.t73 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X450 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X451 dvss.t117 a_21211_n1943.t8 a_21145_n1869.t1 dvss.t116 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X452 a_14285_n2281.t1 ena_ip.t19 a_14285_n2079.t1 dvdd.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X453 avdd_ip.t13 vbreg.t23 avdd_ip.t12 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X454 a_2132_n16254.t1 a_18932_n16088.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X455 a_20689_n2549.t0 a_20471_n2791.t5 dvdd.t7 dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X456 dvdd.t100 x7.x3.B2.t7 a_15000_n1881.t2 dvdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X457 dvdd.t142 x4.in_b.t24 a_14285_n2281.t3 dvdd.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X458 dvdd.t61 a_18481_n2549.t5 a_18371_n2425.t0 dvdd.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X459 dvdd_ip.t28 vbp.t16 tail.t2 dvdd_ip.t27 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X460 xout.t11 vbreg.t24 avdd_ip.t10 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X461 a_18990_n2247.t1 a_17913_n2241.t5 a_18828_n1869.t0 dvdd.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X462 a_20689_n2273.t1 a_20471_n1869.t5 dvdd.t128 dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X463 dvss_ip a_10658_n5446.t13 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X464 vg1.t9 xin.t1 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X465 dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X466 a_2132_n17914.t0 a_18932_n17748.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X467 a_2132_n14262.t1 a_18932_n14428.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X468 a_21198_n2425.t0 a_20121_n2791.t5 a_21036_n2791.t1 dvdd.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X469 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X470 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X471 dvss.t4 a_16795_n2817.t8 a_16729_n2791.t0 dvss.t3 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X472 inv_in.t14 a_17576_n6897.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X473 dvdd_ip.t26 vbp.t17 dvdd_ip.t25 dvdd_ip.t24 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X474 dvss ena_33.t7 avss.t9 avss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X475 dvdd_ip.t19 standby_ip.t17 dvdd.t116 dvdd.t115 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X476 dvss vg2.t1 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X477 a_2132_n15922.t1 a_18932_n16088.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X478 a_18371_n2425.t2 x4.in_b.t25 dvdd.t143 dvdd.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X479 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X480 a_18371_n2425.t1 a_17747_n2791.t7 a_18263_n2791.t3 dvdd.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X481 a_10658_n5446.t1 a_10658_n5446.t0 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X482 dvss.t106 a_16795_n1943.t7 a_16729_n1869.t0 dvss.t105 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X483 dout.t0 dout_filt.t4 dvdd_ip.t1 dvdd_ip.t0 sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X484 a_2132_n14262.t0 vg2.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
X485 dvdd.t72 a_16795_n1943.t8 a_16782_n2247.t0 dvdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X486 avdd_ip.t9 vbreg.t25 avdd_ip.t8 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X487 xout.t26 avdd_ip.t4 sky130_fd_pr__diode_pd2nw_05v5 perim=1.8e+06 area=2.025e+11
X488 a_20471_n2791.t3 a_19955_n2791.t7 a_20376_n2791.t3 dvss.t276 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X489 x7.x1.x3.CLK.t1 a_17359_n2247.t3 dvss.t10 dvss.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X490 a_20471_n1869.t2 a_20121_n2241.t5 a_20376_n1881.t1 dvdd.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X491 avss.t15 ena_33.t8 dvss avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X492 dvdd.t74 standby_ip.t18 dvdd_ip.t14 dvdd.t73 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X493 a_2130_n21508.t0 a_24530_n21342.t0 dvss sky130_fd_pr__res_xhigh_po_0p35 l=110
X494 a_10620_n7674.t0 inv_in.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X495 dvdd.t153 a_19003_n1943.t8 a_18990_n2247.t0 dvdd.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X496 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X497 a_18168_n2791.t2 x7.x2.x4.CLK.t5 dvss.t97 dvss.t96 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X498 vrb.t1 vg2.t9 vbreg.t3 dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X499 a_2132_n15922.t0 a_18932_n15756.t1 dvss sky130_fd_pr__res_xhigh_po_0p35 l=82
R0 a_15705_n2241.t0 a_15705_n2241.n3 370.026
R1 a_15705_n2241.n0 a_15705_n2241.t2 351.356
R2 a_15705_n2241.n1 a_15705_n2241.t4 334.717
R3 a_15705_n2241.n3 a_15705_n2241.t1 325.971
R4 a_15705_n2241.n1 a_15705_n2241.t3 309.935
R5 a_15705_n2241.n0 a_15705_n2241.t5 305.683
R6 a_15705_n2241.n2 a_15705_n2241.n0 16.879
R7 a_15705_n2241.n3 a_15705_n2241.n2 10.8867
R8 a_15705_n2241.n2 a_15705_n2241.n1 9.3005
R9 a_16273_n2273.n3 a_16273_n2273.n2 647.119
R10 a_16273_n2273.n1 a_16273_n2273.t4 350.253
R11 a_16273_n2273.n2 a_16273_n2273.n0 260.339
R12 a_16273_n2273.n2 a_16273_n2273.n1 246.119
R13 a_16273_n2273.n1 a_16273_n2273.t5 189.588
R14 a_16273_n2273.n3 a_16273_n2273.t1 89.1195
R15 a_16273_n2273.n0 a_16273_n2273.t2 63.3338
R16 a_16273_n2273.t3 a_16273_n2273.n3 41.0422
R17 a_16273_n2273.n0 a_16273_n2273.t0 31.9797
R18 a_16620_n1869.n3 a_16620_n1869.n2 636.953
R19 a_16620_n1869.n1 a_16620_n1869.t4 366.856
R20 a_16620_n1869.n2 a_16620_n1869.n0 300.2
R21 a_16620_n1869.n2 a_16620_n1869.n1 225.036
R22 a_16620_n1869.n1 a_16620_n1869.t5 174.056
R23 a_16620_n1869.n0 a_16620_n1869.t1 70.0005
R24 a_16620_n1869.t0 a_16620_n1869.n3 68.0124
R25 a_16620_n1869.n3 a_16620_n1869.t2 63.3219
R26 a_16620_n1869.n0 a_16620_n1869.t3 61.6672
R27 dvss.n521 dvss.n520 184280
R28 dvss.n522 dvss.n521 123547
R29 dvss.n521 dvss.n123 10946.5
R30 dvss.n50 dvss.n16 8366.71
R31 dvss.n50 dvss.n17 8366.71
R32 dvss.n46 dvss.n17 8366.71
R33 dvss.n46 dvss.n16 8366.71
R34 dvss.n113 dvss.n112 7123.23
R35 dvss.n112 dvss.n111 5697.48
R36 dvss.n35 dvss.n30 4247.09
R37 dvss.n42 dvss.n30 4247.09
R38 dvss.n35 dvss.n31 4247.09
R39 dvss.n42 dvss.n31 4247.09
R40 dvss.n191 dvss.n185 4247.09
R41 dvss.n196 dvss.n185 4247.09
R42 dvss.n191 dvss.n186 4247.09
R43 dvss.n196 dvss.n186 4247.09
R44 dvss.n84 dvss.n14 2798.56
R45 dvss.n524 dvss.n14 2798.56
R46 dvss.n84 dvss.n15 2798.56
R47 dvss.n524 dvss.n15 2798.56
R48 dvss.n121 dvss.n53 2798.56
R49 dvss.n114 dvss.n53 2798.56
R50 dvss.n121 dvss.n54 2798.56
R51 dvss.n114 dvss.n54 2798.56
R52 dvss.n45 dvss.n43 2575.49
R53 dvss.n387 dvss.n386 2387.64
R54 dvss.n123 dvss.n122 2025.4
R55 dvss.n123 dvss.n51 2021.82
R56 dvss.n112 dvss.n85 1754.3
R57 dvss.n388 dvss.n387 1680.95
R58 dvss.n92 dvss.n87 1407.97
R59 dvss.n109 dvss.n87 1407.97
R60 dvss.n109 dvss.n88 1407.97
R61 dvss.n65 dvss.n62 1407.97
R62 dvss.n65 dvss.n63 1407.97
R63 dvss.n66 dvss.n62 1407.97
R64 dvss.n66 dvss.n63 1407.97
R65 dvss.n552 dvss.n0 1212.38
R66 dvss.n81 dvss.n80 1198.25
R67 dvss.n198 dvss.n7 1198.25
R68 dvss.n386 dvss.n385 1198.25
R69 dvss.n221 dvss.n202 1198.25
R70 dvss.n336 dvss.n222 1198.25
R71 dvss.n296 dvss.n239 1198.25
R72 dvss.n256 dvss.n124 1198.25
R73 dvss.n519 dvss.n518 1198.25
R74 dvss.n188 dvss.n143 1198.25
R75 dvss.n189 dvss.n160 1198.25
R76 dvss.n399 dvss.n179 1198.25
R77 dvss.n389 dvss.n388 1198.25
R78 dvss.n104 dvss.n86 1198.25
R79 dvss.n552 dvss.n551 1175.19
R80 dvss.t171 dvss.t247 935.78
R81 dvss.t273 dvss.t243 935.78
R82 dvss.t84 dvss.t268 935.78
R83 dvss.n49 dvss.n48 784.03
R84 dvss.n24 dvss.n23 783.962
R85 dvss.n48 dvss.n47 783.75
R86 dvss.n29 dvss.n24 783.683
R87 dvss.n221 dvss.t107 748.625
R88 dvss.t123 dvss.t166 717.851
R89 dvss.t80 dvss.t96 717.851
R90 dvss.t132 dvss.t164 717.851
R91 dvss.t223 dvss.t228 689.909
R92 dvss.t38 dvss.t223 689.909
R93 dvss.t270 dvss.t102 689.909
R94 dvss.t102 dvss.t23 689.909
R95 dvss.t142 dvss.t48 689.909
R96 dvss.t48 dvss.t8 689.909
R97 dvss.n523 dvss.n522 640.604
R98 dvss.n85 dvss.t175 620.187
R99 dvss.n523 dvss.t175 620.187
R100 dvss.t155 dvss.t41 609.174
R101 dvss.t140 dvss.t119 609.174
R102 dvss.t65 dvss.t209 609.174
R103 dvss.t56 dvss.n179 574.28
R104 dvss.t46 dvss.n124 554.129
R105 dvss.n239 dvss.t218 554.129
R106 dvss.n222 dvss.t9 554.129
R107 dvss.t116 dvss.t236 546.789
R108 dvss.t215 dvss.t177 546.789
R109 dvss.t220 dvss.t105 546.789
R110 dvss.t225 dvss.t68 529.24
R111 dvss.t11 dvss.t225 529.24
R112 dvss.t100 dvss.t266 529.24
R113 dvss.t86 dvss.t100 529.24
R114 dvss.t206 dvss.t112 529.24
R115 dvss.t289 dvss.t206 529.24
R116 dvss.t173 dvss.t262 484.404
R117 dvss.t192 dvss.t190 484.404
R118 dvss.t188 dvss.t182 484.404
R119 dvss.t217 dvss.t5 467.307
R120 dvss.t208 dvss.t148 467.307
R121 dvss.t45 dvss.t169 467.307
R122 dvss.t107 dvss.t245 447.707
R123 dvss.n387 dvss.n198 426.382
R124 dvss.n519 dvss.t35 425.08
R125 dvss.t54 dvss.n188 425.08
R126 dvss.t82 dvss.n189 425.08
R127 dvss.t211 dvss.t14 419.45
R128 dvss.t138 dvss.t146 419.45
R129 dvss.t3 dvss.t144 419.45
R130 dvss.n110 dvss.n86 419.18
R131 dvss.t227 dvss.t170 400
R132 dvss.t239 dvss.t125 400
R133 dvss.t272 dvss.t210 400
R134 dvss.n92 dvss.n91 390.825
R135 dvss.t50 dvss.t6 371.594
R136 dvss.t114 dvss.t258 371.594
R137 dvss.t251 dvss.t66 371.594
R138 dvss.n522 dvss.t62 366.435
R139 dvss.t262 dvss.t227 363.303
R140 dvss.t125 dvss.t192 363.303
R141 dvss.t210 dvss.t188 363.303
R142 dvss.t228 dvss.t46 355.964
R143 dvss.t218 dvss.t270 355.964
R144 dvss.t9 dvss.t142 355.964
R145 dvss.t170 dvss.t116 352.295
R146 dvss.t149 dvss.t155 352.295
R147 dvss.t177 dvss.t239 352.295
R148 dvss.t119 dvss.t34 352.295
R149 dvss.t105 dvss.t272 352.295
R150 dvss.t209 dvss.t238 352.295
R151 dvss.t247 dvss.t149 348.625
R152 dvss.t34 dvss.t273 348.625
R153 dvss.t238 dvss.t84 348.625
R154 dvss.n111 dvss.n110 344.228
R155 dvss.t134 dvss.t56 343.442
R156 dvss.t236 dvss.t38 333.945
R157 dvss.t23 dvss.t215 333.945
R158 dvss.t8 dvss.t220 333.945
R159 dvss.n520 dvss.n124 308.257
R160 dvss.t91 dvss.t171 308.257
R161 dvss.t243 dvss.t260 308.257
R162 dvss.t268 dvss.t184 308.257
R163 dvss.n86 dvss 308.139
R164 dvss.n205 dvss.t85 307.536
R165 dvss.n330 dvss.t274 307.536
R166 dvss.n290 dvss.t248 307.536
R167 dvss.n140 dvss.t167 307.536
R168 dvss.n157 dvss.t97 307.536
R169 dvss.n405 dvss.t133 307.536
R170 dvss.t162 dvss.t275 306.846
R171 dvss.t118 dvss.t255 306.846
R172 dvss.t198 dvss.t64 306.846
R173 dvss.n63 dvss.n61 292.5
R174 dvss.n63 dvss.n58 292.5
R175 dvss.n67 dvss.n66 292.5
R176 dvss.n66 dvss.t0 292.5
R177 dvss.n62 dvss.n60 292.5
R178 dvss.n62 dvss.n52 292.5
R179 dvss.n65 dvss.n64 292.5
R180 dvss.t0 dvss.n65 292.5
R181 dvss.n90 dvss.n88 292.5
R182 dvss.n109 dvss.n108 292.5
R183 dvss.n110 dvss.n109 292.5
R184 dvss.n89 dvss.n87 292.5
R185 dvss.n87 dvss.t93 292.5
R186 dvss.n93 dvss.n92 292.5
R187 dvss.t88 dvss 289.909
R188 dvss.t6 dvss.t162 278.695
R189 dvss.t258 dvss.t118 278.695
R190 dvss.t66 dvss.t198 278.695
R191 dvss.n195 dvss.n193 276.286
R192 dvss.n239 dvss 275.229
R193 dvss dvss.n222 275.229
R194 dvss dvss.n221 275.229
R195 dvss.n386 dvss 275.229
R196 dvss.t256 dvss.n0 273.678
R197 dvss.n43 dvss.t256 273.678
R198 dvss.t68 dvss.t35 273.065
R199 dvss.t266 dvss.t54 273.065
R200 dvss.t112 dvss.t82 273.065
R201 dvss.t275 dvss.t211 270.25
R202 dvss.t276 dvss.t217 270.25
R203 dvss.t255 dvss.t138 270.25
R204 dvss.t179 dvss.t208 270.25
R205 dvss.t64 dvss.t3 270.25
R206 dvss.t166 dvss.t276 267.435
R207 dvss.t96 dvss.t179 267.435
R208 dvss.t163 dvss.t132 267.435
R209 dvss.t41 dvss.t173 264.221
R210 dvss.t190 dvss.t140 264.221
R211 dvss.t182 dvss.t65 264.221
R212 dvss.t245 dvss.t88 264.221
R213 dvss.t14 dvss.t11 256.175
R214 dvss.t146 dvss.t86 256.175
R215 dvss.t144 dvss.t289 256.175
R216 dvss.n45 dvss.t204 255.168
R217 dvss.n51 dvss.t150 255.168
R218 dvss.n215 dvss.t49 246.817
R219 dvss.n303 dvss.t103 246.817
R220 dvss.n263 dvss.t224 246.817
R221 dvss.n130 dvss.t226 246.817
R222 dvss.n470 dvss.t101 246.817
R223 dvss.n431 dvss.t207 246.817
R224 dvss.t94 dvss.t62 244.291
R225 dvss dvss.t91 238.532
R226 dvss.t260 dvss 238.532
R227 dvss.t184 dvss 238.532
R228 dvss.n520 dvss.n519 236.469
R229 dvss.t24 dvss.t123 236.469
R230 dvss.t234 dvss.t80 236.469
R231 dvss.t164 dvss.t58 236.469
R232 dvss.n122 dvss.n52 231.216
R233 dvss.n409 dvss.t33 229.185
R234 dvss.n32 dvss.t257 219.8
R235 dvss.n41 dvss.n33 217.329
R236 dvss.n193 dvss.n192 217.225
R237 dvss.n218 dvss.n217 214.742
R238 dvss.n236 dvss.n235 214.742
R239 dvss.n253 dvss.n252 214.742
R240 dvss.n129 dvss.n128 214.742
R241 dvss.n476 dvss.n145 214.742
R242 dvss.n437 dvss.n162 214.742
R243 dvss.n188 dvss 211.132
R244 dvss.n189 dvss 211.132
R245 dvss dvss.n179 211.132
R246 dvss.n388 dvss 211.132
R247 dvss.n213 dvss.n212 209.254
R248 dvss.n310 dvss.n232 209.254
R249 dvss.n270 dvss.n249 209.254
R250 dvss.n133 dvss.n132 209.254
R251 dvss.n151 dvss.n150 209.254
R252 dvss.n168 dvss.n167 209.254
R253 dvss.t204 dvss.t196 208.894
R254 dvss.t196 dvss.t152 208.894
R255 dvss.t152 dvss.t16 208.894
R256 dvss.t16 dvss.t52 208.894
R257 dvss.t60 dvss.t249 208.894
R258 dvss.t249 dvss.t202 208.894
R259 dvss.t202 dvss.t194 208.894
R260 dvss.t194 dvss.t150 208.894
R261 dvss.t5 dvss.t50 202.688
R262 dvss.t148 dvss.t114 202.688
R263 dvss.t169 dvss.t251 202.688
R264 dvss.t87 dvss.t134 202.688
R265 dvss.n537 dvss.n6 202.067
R266 dvss.n3 dvss.n2 200.516
R267 dvss.n76 dvss.n75 199.739
R268 dvss.n371 dvss.n204 199.739
R269 dvss.n358 dvss.n209 199.739
R270 dvss.n224 dvss.n223 199.739
R271 dvss.n318 dvss.n317 199.739
R272 dvss.n241 dvss.n240 199.739
R273 dvss.n278 dvss.n277 199.739
R274 dvss.n496 dvss.n137 199.739
R275 dvss.n483 dvss.n142 199.739
R276 dvss.n457 dvss.n154 199.739
R277 dvss.n444 dvss.n159 199.739
R278 dvss.n418 dvss.n171 199.739
R279 dvss.n178 dvss.n177 199.739
R280 dvss.n101 dvss.n100 199.739
R281 dvss.n41 dvss.n40 198.024
R282 dvss.t28 dvss.n52 188.078
R283 dvss.n379 dvss.n378 185
R284 dvss.n184 dvss.n183 185
R285 dvss.n550 dvss.n549 185
R286 dvss dvss.t24 182.982
R287 dvss dvss.t234 182.982
R288 dvss.n83 dvss.n11 181.835
R289 dvss.n83 dvss.n82 181.835
R290 dvss.n115 dvss.n57 181.835
R291 dvss.n116 dvss.n115 181.835
R292 dvss.n91 dvss.n88 174.962
R293 dvss.n190 dvss.t163 166.091
R294 dvss.n197 dvss.t87 154.831
R295 dvss.n33 dvss.n30 148.029
R296 dvss.n196 dvss.n195 146.25
R297 dvss.n197 dvss.n196 146.25
R298 dvss.n192 dvss.n191 146.25
R299 dvss.n191 dvss.n190 146.25
R300 dvss.n34 dvss.n31 146.25
R301 dvss.n31 dvss.t256 146.25
R302 dvss.n30 dvss.t256 146.25
R303 dvss.n36 dvss.n33 143.809
R304 dvss dvss.t1 141.49
R305 dvss.t58 dvss.t32 140.756
R306 dvss dvss.t30 140.144
R307 dvss.n195 dvss.n194 127.487
R308 dvss.n113 dvss.n81 122.51
R309 dvss.n115 dvss.n114 117.001
R310 dvss.n114 dvss.n113 117.001
R311 dvss.n116 dvss.n54 117.001
R312 dvss.t28 dvss.n54 117.001
R313 dvss.n121 dvss.n120 117.001
R314 dvss.n122 dvss.n121 117.001
R315 dvss.n57 dvss.n53 117.001
R316 dvss.t28 dvss.n53 117.001
R317 dvss.n525 dvss.n524 117.001
R318 dvss.n524 dvss.n523 117.001
R319 dvss.n15 dvss.n11 117.001
R320 dvss.t175 dvss.n15 117.001
R321 dvss.n84 dvss.n83 117.001
R322 dvss.n85 dvss.n84 117.001
R323 dvss.n82 dvss.n14 117.001
R324 dvss.t175 dvss.n14 117.001
R325 dvss.t52 dvss.n44 104.448
R326 dvss.n44 dvss.t60 104.448
R327 dvss.n190 dvss.t45 104.159
R328 dvss.n525 dvss.n12 102.025
R329 dvss.n526 dvss.n525 102.025
R330 dvss.n120 dvss.n55 102.025
R331 dvss.n120 dvss.n119 102.025
R332 dvss.n212 dvss.t221 100.001
R333 dvss.n232 dvss.t216 100.001
R334 dvss.n249 dvss.t237 100.001
R335 dvss.n132 dvss.t15 100.001
R336 dvss.n150 dvss.t147 100.001
R337 dvss.n167 dvss.t145 100.001
R338 dvss.n64 dvss.n61 91.4829
R339 dvss.n93 dvss.n89 91.4829
R340 dvss.n70 dvss.t29 83.7183
R341 dvss.n95 dvss.t176 83.7183
R342 dvss.n91 dvss.t93 81.1932
R343 dvss dvss.t94 80.5052
R344 dvss.n526 dvss.n11 79.8123
R345 dvss.n82 dvss.n12 79.8123
R346 dvss.n57 dvss.n55 79.8123
R347 dvss.n119 dvss.n116 79.8123
R348 dvss.n378 dvss.t108 72.8576
R349 dvss.n209 dvss.t183 72.8576
R350 dvss.n317 dvss.t191 72.8576
R351 dvss.n277 dvss.t174 72.8576
R352 dvss.n183 dvss.t57 72.8576
R353 dvss.n137 dvss.t51 72.8576
R354 dvss.n154 dvss.t115 72.8576
R355 dvss.n171 dvss.t252 72.8576
R356 dvss.n212 dvss.t106 70.0005
R357 dvss.n232 dvss.t178 70.0005
R358 dvss.n249 dvss.t117 70.0005
R359 dvss.n132 dvss.t212 70.0005
R360 dvss.n150 dvss.t139 70.0005
R361 dvss.n167 dvss.t4 70.0005
R362 dvss.n67 dvss.n61 69.6045
R363 dvss.n108 dvss.n89 69.0306
R364 dvss.t0 dvss 69.0201
R365 dvss.n187 dvss.n175 68.8106
R366 dvss dvss.n197 67.5629
R367 dvss.n64 dvss.n60 66.3131
R368 dvss.n94 dvss.n93 65.475
R369 dvss.n209 dvss.t189 60.5809
R370 dvss.n317 dvss.t193 60.5809
R371 dvss.n277 dvss.t263 60.5809
R372 dvss.n137 dvss.t7 60.5809
R373 dvss.n154 dvss.t259 60.5809
R374 dvss.n171 dvss.t67 60.5809
R375 dvss.n378 dvss.t246 58.5719
R376 dvss.n183 dvss.t135 58.5719
R377 dvss.n217 dvss.t143 57.1434
R378 dvss.n235 dvss.t271 57.1434
R379 dvss.n252 dvss.t229 57.1434
R380 dvss.n128 dvss.t69 57.1434
R381 dvss.n145 dvss.t267 57.1434
R382 dvss.n162 dvss.t113 57.1434
R383 dvss.n549 dvss.t42 52.8576
R384 dvss.n549 dvss.t31 51.4291
R385 dvss.t32 dvss 42.227
R386 dvss.n194 dvss.n186 41.7862
R387 dvss.t32 dvss.n186 41.7862
R388 dvss.n193 dvss.n185 41.7862
R389 dvss.t32 dvss.n185 41.7862
R390 dvss.n42 dvss.n41 41.7862
R391 dvss.n43 dvss.n42 41.7862
R392 dvss.n36 dvss.n35 41.7862
R393 dvss.n35 dvss.n0 41.7862
R394 dvss.n50 dvss.n49 41.7862
R395 dvss.n51 dvss.n50 41.7862
R396 dvss.n47 dvss.n46 41.7862
R397 dvss.n46 dvss.n45 41.7862
R398 dvss.n548 dvss.n547 40.0735
R399 dvss.n204 dvss.t269 38.5719
R400 dvss.n204 dvss.t185 38.5719
R401 dvss.n223 dvss.t244 38.5719
R402 dvss.n223 dvss.t261 38.5719
R403 dvss.n240 dvss.t172 38.5719
R404 dvss.n240 dvss.t92 38.5719
R405 dvss.n142 dvss.t124 38.5719
R406 dvss.n142 dvss.t25 38.5719
R407 dvss.n159 dvss.t81 38.5719
R408 dvss.n159 dvss.t235 38.5719
R409 dvss.n177 dvss.t165 38.5719
R410 dvss.n177 dvss.t59 38.5719
R411 dvss.n107 dvss.n90 37.6894
R412 dvss.n69 dvss.n68 37.4862
R413 dvss.t0 dvss.t28 36.2358
R414 dvss.n81 dvss.n58 36.2358
R415 dvss.n6 dvss.t141 36.0005
R416 dvss.n541 dvss.n5 34.6358
R417 dvss.n542 dvss.n541 34.6358
R418 dvss.n543 dvss.n542 34.6358
R419 dvss.n384 dvss.n200 34.6358
R420 dvss.n377 dvss.n376 34.6358
R421 dvss.n360 dvss.n359 34.6358
R422 dvss.n360 dvss.n207 34.6358
R423 dvss.n364 dvss.n207 34.6358
R424 dvss.n365 dvss.n364 34.6358
R425 dvss.n366 dvss.n365 34.6358
R426 dvss.n352 dvss.n351 34.6358
R427 dvss.n353 dvss.n352 34.6358
R428 dvss.n353 dvss.n210 34.6358
R429 dvss.n357 dvss.n210 34.6358
R430 dvss.n338 dvss.n337 34.6358
R431 dvss.n342 dvss.n341 34.6358
R432 dvss.n343 dvss.n342 34.6358
R433 dvss.n347 dvss.n346 34.6358
R434 dvss.n348 dvss.n347 34.6358
R435 dvss.n323 dvss.n228 34.6358
R436 dvss.n324 dvss.n323 34.6358
R437 dvss.n325 dvss.n324 34.6358
R438 dvss.n325 dvss.n226 34.6358
R439 dvss.n329 dvss.n226 34.6358
R440 dvss.n311 dvss.n230 34.6358
R441 dvss.n315 dvss.n230 34.6358
R442 dvss.n316 dvss.n315 34.6358
R443 dvss.n319 dvss.n316 34.6358
R444 dvss.n298 dvss.n297 34.6358
R445 dvss.n302 dvss.n301 34.6358
R446 dvss.n304 dvss.n302 34.6358
R447 dvss.n308 dvss.n233 34.6358
R448 dvss.n309 dvss.n308 34.6358
R449 dvss.n283 dvss.n245 34.6358
R450 dvss.n284 dvss.n283 34.6358
R451 dvss.n285 dvss.n284 34.6358
R452 dvss.n285 dvss.n243 34.6358
R453 dvss.n289 dvss.n243 34.6358
R454 dvss.n271 dvss.n247 34.6358
R455 dvss.n275 dvss.n247 34.6358
R456 dvss.n276 dvss.n275 34.6358
R457 dvss.n279 dvss.n276 34.6358
R458 dvss.n258 dvss.n257 34.6358
R459 dvss.n262 dvss.n261 34.6358
R460 dvss.n264 dvss.n262 34.6358
R461 dvss.n268 dvss.n250 34.6358
R462 dvss.n269 dvss.n268 34.6358
R463 dvss.n517 dvss.n126 34.6358
R464 dvss.n513 dvss.n512 34.6358
R465 dvss.n512 dvss.n511 34.6358
R466 dvss.n508 dvss.n507 34.6358
R467 dvss.n507 dvss.n506 34.6358
R468 dvss.n503 dvss.n502 34.6358
R469 dvss.n502 dvss.n501 34.6358
R470 dvss.n501 dvss.n135 34.6358
R471 dvss.n497 dvss.n135 34.6358
R472 dvss.n495 dvss.n494 34.6358
R473 dvss.n494 dvss.n138 34.6358
R474 dvss.n490 dvss.n138 34.6358
R475 dvss.n490 dvss.n489 34.6358
R476 dvss.n489 dvss.n488 34.6358
R477 dvss.n478 dvss.n477 34.6358
R478 dvss.n475 dvss.n146 34.6358
R479 dvss.n471 dvss.n146 34.6358
R480 dvss.n469 dvss.n468 34.6358
R481 dvss.n468 dvss.n148 34.6358
R482 dvss.n464 dvss.n463 34.6358
R483 dvss.n463 dvss.n462 34.6358
R484 dvss.n462 dvss.n152 34.6358
R485 dvss.n458 dvss.n152 34.6358
R486 dvss.n456 dvss.n455 34.6358
R487 dvss.n455 dvss.n155 34.6358
R488 dvss.n451 dvss.n155 34.6358
R489 dvss.n451 dvss.n450 34.6358
R490 dvss.n450 dvss.n449 34.6358
R491 dvss.n439 dvss.n438 34.6358
R492 dvss.n436 dvss.n163 34.6358
R493 dvss.n432 dvss.n163 34.6358
R494 dvss.n430 dvss.n429 34.6358
R495 dvss.n429 dvss.n165 34.6358
R496 dvss.n425 dvss.n424 34.6358
R497 dvss.n424 dvss.n169 34.6358
R498 dvss.n420 dvss.n169 34.6358
R499 dvss.n420 dvss.n419 34.6358
R500 dvss.n417 dvss.n172 34.6358
R501 dvss.n413 dvss.n172 34.6358
R502 dvss.n413 dvss.n412 34.6358
R503 dvss.n412 dvss.n174 34.6358
R504 dvss.n406 dvss.n174 34.6358
R505 dvss.n398 dvss.n181 34.6358
R506 dvss.n393 dvss.n392 34.6358
R507 dvss.n75 dvss.t2 33.462
R508 dvss.n75 dvss.t156 33.462
R509 dvss.n100 dvss.t95 33.462
R510 dvss.n100 dvss.t63 33.462
R511 dvss.n2 dvss.t214 33.2313
R512 dvss.n341 dvss.n218 31.2476
R513 dvss.n301 dvss.n236 31.2476
R514 dvss.n261 dvss.n253 31.2476
R515 dvss.n513 dvss.n129 31.2476
R516 dvss.n476 dvss.n475 31.2476
R517 dvss.n437 dvss.n436 31.2476
R518 dvss.t98 dvss.t30 30.4092
R519 dvss dvss.n552 30.4092
R520 dvss.n370 dvss.n205 29.7417
R521 dvss.n331 dvss.n330 29.7417
R522 dvss.n291 dvss.n290 29.7417
R523 dvss.n484 dvss.n140 29.7417
R524 dvss.n445 dvss.n157 29.7417
R525 dvss.n405 dvss.n404 29.7417
R526 dvss.n346 dvss.n215 27.8593
R527 dvss.n303 dvss.n233 27.8593
R528 dvss.n263 dvss.n250 27.8593
R529 dvss.n508 dvss.n130 27.8593
R530 dvss.n470 dvss.n469 27.8593
R531 dvss.n431 dvss.n430 27.8593
R532 dvss.n547 dvss.n3 25.977
R533 dvss.n217 dvss.t10 25.4291
R534 dvss.n235 dvss.t219 25.4291
R535 dvss.n252 dvss.t47 25.4291
R536 dvss.n128 dvss.t36 25.4291
R537 dvss.n145 dvss.t55 25.4291
R538 dvss.n162 dvss.t83 25.4291
R539 dvss.n2 dvss.t168 24.9236
R540 dvss.n6 dvss.t99 24.9236
R541 dvss.n24 dvss.n16 24.3755
R542 dvss.n44 dvss.n16 24.3755
R543 dvss.n48 dvss.n17 24.3755
R544 dvss.n44 dvss.n17 24.3755
R545 dvss.n380 dvss.n200 23.7737
R546 dvss.n394 dvss.n393 23.7737
R547 dvss.n80 dvss.n79 23.7181
R548 dvss.n536 dvss.n7 23.7181
R549 dvss.n385 dvss.n384 23.7181
R550 dvss.n376 dvss.n202 23.7181
R551 dvss.n372 dvss.n202 23.7181
R552 dvss.n337 dvss.n336 23.7181
R553 dvss.n336 dvss.n335 23.7181
R554 dvss.n297 dvss.n296 23.7181
R555 dvss.n296 dvss.n295 23.7181
R556 dvss.n257 dvss.n256 23.7181
R557 dvss.n518 dvss.n517 23.7181
R558 dvss.n482 dvss.n143 23.7181
R559 dvss.n478 dvss.n143 23.7181
R560 dvss.n443 dvss.n160 23.7181
R561 dvss.n439 dvss.n160 23.7181
R562 dvss.n400 dvss.n399 23.7181
R563 dvss.n399 dvss.n398 23.7181
R564 dvss.n392 dvss.n389 23.7181
R565 dvss.n104 dvss.n103 23.7181
R566 dvss.n537 dvss.n5 22.9652
R567 dvss.n371 dvss.n370 22.9652
R568 dvss.n331 dvss.n224 22.9652
R569 dvss.n291 dvss.n241 22.9652
R570 dvss.n484 dvss.n483 22.9652
R571 dvss.n445 dvss.n444 22.9652
R572 dvss.n404 dvss.n178 22.9652
R573 dvss.n537 dvss.n536 21.4593
R574 dvss.n372 dvss.n371 21.4593
R575 dvss.n335 dvss.n224 21.4593
R576 dvss.n295 dvss.n241 21.4593
R577 dvss.n483 dvss.n482 21.4593
R578 dvss.n444 dvss.n443 21.4593
R579 dvss.n400 dvss.n178 21.4593
R580 dvss.n551 dvss.n550 21.4265
R581 dvss.n47 dvss.t205 21.1687
R582 dvss.n49 dvss.t151 21.1687
R583 dvss.n198 dvss.t98 21.1543
R584 dvss.n379 dvss.n377 20.9718
R585 dvss.n184 dvss.n181 20.9718
R586 dvss.n32 dvss.n8 19.9405
R587 dvss.n22 dvss.n18 18.4515
R588 dvss.n21 dvss.n19 18.4515
R589 dvss.n27 dvss.n26 18.4515
R590 dvss.n28 dvss.n25 18.4515
R591 dvss.n543 dvss.n3 18.4476
R592 dvss.n348 dvss.n213 17.6946
R593 dvss.n310 dvss.n309 17.6946
R594 dvss.n270 dvss.n269 17.6946
R595 dvss.n506 dvss.n133 17.6946
R596 dvss.n151 dvss.n148 17.6946
R597 dvss.n168 dvss.n165 17.6946
R598 dvss.n111 dvss.t93 16.6567
R599 dvss.n76 dvss 15.0593
R600 dvss.n101 dvss 15.0593
R601 dvss.n366 dvss.n205 14.6829
R602 dvss.n330 dvss.n329 14.6829
R603 dvss.n290 dvss.n289 14.6829
R604 dvss.n488 dvss.n140 14.6829
R605 dvss.n449 dvss.n157 14.6829
R606 dvss.n406 dvss.n405 14.6829
R607 dvss.t1 dvss.n58 13.8044
R608 dvss.n39 dvss.n8 13.3461
R609 dvss.n38 dvss.n37 13.0158
R610 dvss.n33 dvss.n32 11.7338
R611 dvss.n40 dvss.n39 10.1755
R612 dvss.n119 dvss 9.488
R613 dvss.n79 dvss.n78 9.3005
R614 dvss.n80 dvss.n59 9.3005
R615 dvss.n390 dvss.n389 9.3005
R616 dvss.n408 dvss.n174 9.3005
R617 dvss.n407 dvss.n406 9.3005
R618 dvss.n405 dvss.n176 9.3005
R619 dvss.n404 dvss.n403 9.3005
R620 dvss.n402 dvss.n178 9.3005
R621 dvss.n401 dvss.n400 9.3005
R622 dvss.n399 dvss.n180 9.3005
R623 dvss.n398 dvss.n397 9.3005
R624 dvss.n396 dvss.n181 9.3005
R625 dvss.n395 dvss.n394 9.3005
R626 dvss.n393 dvss.n182 9.3005
R627 dvss.n392 dvss.n391 9.3005
R628 dvss.n518 dvss.n125 9.3005
R629 dvss.n517 dvss.n516 9.3005
R630 dvss.n515 dvss.n126 9.3005
R631 dvss.n514 dvss.n513 9.3005
R632 dvss.n512 dvss.n127 9.3005
R633 dvss.n511 dvss.n510 9.3005
R634 dvss.n509 dvss.n508 9.3005
R635 dvss.n507 dvss.n131 9.3005
R636 dvss.n506 dvss.n505 9.3005
R637 dvss.n504 dvss.n503 9.3005
R638 dvss.n502 dvss.n134 9.3005
R639 dvss.n501 dvss.n500 9.3005
R640 dvss.n499 dvss.n135 9.3005
R641 dvss.n498 dvss.n497 9.3005
R642 dvss.n495 dvss.n136 9.3005
R643 dvss.n494 dvss.n493 9.3005
R644 dvss.n492 dvss.n138 9.3005
R645 dvss.n491 dvss.n490 9.3005
R646 dvss.n489 dvss.n139 9.3005
R647 dvss.n488 dvss.n487 9.3005
R648 dvss.n486 dvss.n140 9.3005
R649 dvss.n485 dvss.n484 9.3005
R650 dvss.n483 dvss.n141 9.3005
R651 dvss.n482 dvss.n481 9.3005
R652 dvss.n480 dvss.n143 9.3005
R653 dvss.n479 dvss.n478 9.3005
R654 dvss.n477 dvss.n144 9.3005
R655 dvss.n475 dvss.n474 9.3005
R656 dvss.n473 dvss.n146 9.3005
R657 dvss.n472 dvss.n471 9.3005
R658 dvss.n469 dvss.n147 9.3005
R659 dvss.n468 dvss.n467 9.3005
R660 dvss.n466 dvss.n148 9.3005
R661 dvss.n465 dvss.n464 9.3005
R662 dvss.n463 dvss.n149 9.3005
R663 dvss.n462 dvss.n461 9.3005
R664 dvss.n460 dvss.n152 9.3005
R665 dvss.n459 dvss.n458 9.3005
R666 dvss.n456 dvss.n153 9.3005
R667 dvss.n455 dvss.n454 9.3005
R668 dvss.n453 dvss.n155 9.3005
R669 dvss.n452 dvss.n451 9.3005
R670 dvss.n450 dvss.n156 9.3005
R671 dvss.n449 dvss.n448 9.3005
R672 dvss.n447 dvss.n157 9.3005
R673 dvss.n446 dvss.n445 9.3005
R674 dvss.n444 dvss.n158 9.3005
R675 dvss.n443 dvss.n442 9.3005
R676 dvss.n441 dvss.n160 9.3005
R677 dvss.n440 dvss.n439 9.3005
R678 dvss.n438 dvss.n161 9.3005
R679 dvss.n436 dvss.n435 9.3005
R680 dvss.n434 dvss.n163 9.3005
R681 dvss.n433 dvss.n432 9.3005
R682 dvss.n430 dvss.n164 9.3005
R683 dvss.n429 dvss.n428 9.3005
R684 dvss.n427 dvss.n165 9.3005
R685 dvss.n426 dvss.n425 9.3005
R686 dvss.n424 dvss.n423 9.3005
R687 dvss.n422 dvss.n169 9.3005
R688 dvss.n421 dvss.n420 9.3005
R689 dvss.n419 dvss.n170 9.3005
R690 dvss.n417 dvss.n416 9.3005
R691 dvss.n415 dvss.n172 9.3005
R692 dvss.n414 dvss.n413 9.3005
R693 dvss.n412 dvss.n411 9.3005
R694 dvss.n256 dvss.n255 9.3005
R695 dvss.n257 dvss.n254 9.3005
R696 dvss.n259 dvss.n258 9.3005
R697 dvss.n261 dvss.n260 9.3005
R698 dvss.n262 dvss.n251 9.3005
R699 dvss.n265 dvss.n264 9.3005
R700 dvss.n266 dvss.n250 9.3005
R701 dvss.n268 dvss.n267 9.3005
R702 dvss.n269 dvss.n248 9.3005
R703 dvss.n272 dvss.n271 9.3005
R704 dvss.n273 dvss.n247 9.3005
R705 dvss.n275 dvss.n274 9.3005
R706 dvss.n276 dvss.n246 9.3005
R707 dvss.n280 dvss.n279 9.3005
R708 dvss.n281 dvss.n245 9.3005
R709 dvss.n283 dvss.n282 9.3005
R710 dvss.n284 dvss.n244 9.3005
R711 dvss.n286 dvss.n285 9.3005
R712 dvss.n287 dvss.n243 9.3005
R713 dvss.n289 dvss.n288 9.3005
R714 dvss.n290 dvss.n242 9.3005
R715 dvss.n292 dvss.n291 9.3005
R716 dvss.n293 dvss.n241 9.3005
R717 dvss.n295 dvss.n294 9.3005
R718 dvss.n296 dvss.n238 9.3005
R719 dvss.n297 dvss.n237 9.3005
R720 dvss.n299 dvss.n298 9.3005
R721 dvss.n301 dvss.n300 9.3005
R722 dvss.n302 dvss.n234 9.3005
R723 dvss.n305 dvss.n304 9.3005
R724 dvss.n306 dvss.n233 9.3005
R725 dvss.n308 dvss.n307 9.3005
R726 dvss.n309 dvss.n231 9.3005
R727 dvss.n312 dvss.n311 9.3005
R728 dvss.n313 dvss.n230 9.3005
R729 dvss.n315 dvss.n314 9.3005
R730 dvss.n316 dvss.n229 9.3005
R731 dvss.n320 dvss.n319 9.3005
R732 dvss.n321 dvss.n228 9.3005
R733 dvss.n323 dvss.n322 9.3005
R734 dvss.n324 dvss.n227 9.3005
R735 dvss.n326 dvss.n325 9.3005
R736 dvss.n327 dvss.n226 9.3005
R737 dvss.n329 dvss.n328 9.3005
R738 dvss.n330 dvss.n225 9.3005
R739 dvss.n332 dvss.n331 9.3005
R740 dvss.n333 dvss.n224 9.3005
R741 dvss.n335 dvss.n334 9.3005
R742 dvss.n336 dvss.n220 9.3005
R743 dvss.n337 dvss.n219 9.3005
R744 dvss.n339 dvss.n338 9.3005
R745 dvss.n341 dvss.n340 9.3005
R746 dvss.n342 dvss.n216 9.3005
R747 dvss.n344 dvss.n343 9.3005
R748 dvss.n346 dvss.n345 9.3005
R749 dvss.n347 dvss.n214 9.3005
R750 dvss.n349 dvss.n348 9.3005
R751 dvss.n351 dvss.n350 9.3005
R752 dvss.n352 dvss.n211 9.3005
R753 dvss.n354 dvss.n353 9.3005
R754 dvss.n355 dvss.n210 9.3005
R755 dvss.n357 dvss.n356 9.3005
R756 dvss.n359 dvss.n208 9.3005
R757 dvss.n361 dvss.n360 9.3005
R758 dvss.n362 dvss.n207 9.3005
R759 dvss.n364 dvss.n363 9.3005
R760 dvss.n365 dvss.n206 9.3005
R761 dvss.n367 dvss.n366 9.3005
R762 dvss.n368 dvss.n205 9.3005
R763 dvss.n370 dvss.n369 9.3005
R764 dvss.n371 dvss.n203 9.3005
R765 dvss.n373 dvss.n372 9.3005
R766 dvss.n374 dvss.n202 9.3005
R767 dvss.n376 dvss.n375 9.3005
R768 dvss.n377 dvss.n201 9.3005
R769 dvss.n381 dvss.n380 9.3005
R770 dvss.n382 dvss.n200 9.3005
R771 dvss.n384 dvss.n383 9.3005
R772 dvss.n385 dvss.n199 9.3005
R773 dvss.n534 dvss.n7 9.3005
R774 dvss.n538 dvss.n537 9.3005
R775 dvss.n544 dvss.n543 9.3005
R776 dvss.n542 dvss.n4 9.3005
R777 dvss.n541 dvss.n540 9.3005
R778 dvss.n539 dvss.n5 9.3005
R779 dvss.n536 dvss.n535 9.3005
R780 dvss.n545 dvss.n3 9.3005
R781 dvss.n547 dvss.n546 9.3005
R782 dvss.n105 dvss.n104 9.3005
R783 dvss.n103 dvss.n102 9.3005
R784 dvss.n97 dvss.n12 9.3005
R785 dvss.n527 dvss.n526 9.3005
R786 dvss.n72 dvss.n55 9.3005
R787 dvss.n108 dvss.n107 8.88939
R788 dvss.n68 dvss.n67 8.77764
R789 dvss.n359 dvss.n358 7.90638
R790 dvss.n318 dvss.n228 7.90638
R791 dvss.n278 dvss.n245 7.90638
R792 dvss.n496 dvss.n495 7.90638
R793 dvss.n457 dvss.n456 7.90638
R794 dvss.n418 dvss.n417 7.90638
R795 dvss.n102 dvss.n101 7.18226
R796 dvss.n77 dvss.n76 7.17078
R797 dvss.n79 dvss 7.15344
R798 dvss.n103 dvss 7.15344
R799 dvss.n343 dvss.n215 6.77697
R800 dvss.n304 dvss.n303 6.77697
R801 dvss.n264 dvss.n263 6.77697
R802 dvss.n511 dvss.n130 6.77697
R803 dvss.n471 dvss.n470 6.77697
R804 dvss.n432 dvss.n431 6.77697
R805 dvss.n194 dvss.n175 6.7005
R806 dvss.n550 dvss.n548 6.56103
R807 dvss.n40 dvss.n34 5.66204
R808 dvss.n38 dvss.n34 5.19708
R809 dvss.n18 dvss.t203 4.3505
R810 dvss.n18 dvss.t195 4.3505
R811 dvss.n19 dvss.t61 4.3505
R812 dvss.n19 dvss.t250 4.3505
R813 dvss.n26 dvss.t17 4.3505
R814 dvss.n26 dvss.t53 4.3505
R815 dvss.n25 dvss.t197 4.3505
R816 dvss.n25 dvss.t153 4.3505
R817 dvss.n338 dvss.n218 3.38874
R818 dvss.n298 dvss.n236 3.38874
R819 dvss.n258 dvss.n253 3.38874
R820 dvss.n129 dvss.n126 3.38874
R821 dvss.n477 dvss.n476 3.38874
R822 dvss.n438 dvss.n437 3.38874
R823 dvss.n537 dvss 3.29747
R824 dvss.n551 dvss.n1 3.21038
R825 dvss.n74 dvss.n69 3.17391
R826 dvss.n351 dvss.n213 2.63579
R827 dvss.n311 dvss.n310 2.63579
R828 dvss.n271 dvss.n270 2.63579
R829 dvss.n503 dvss.n133 2.63579
R830 dvss.n464 dvss.n151 2.63579
R831 dvss.n425 dvss.n168 2.63579
R832 dvss.n39 dvss.n38 2.50662
R833 dvss.n106 dvss.n94 2.44193
R834 dvss.n68 dvss.n59 2.41042
R835 dvss.n107 dvss.n106 2.3255
R836 dvss.n533 dvss 2.30337
R837 dvss.n548 dvss.n1 1.93239
R838 dvss.n358 dvss.n357 1.88285
R839 dvss.n319 dvss.n318 1.88285
R840 dvss.n279 dvss.n278 1.88285
R841 dvss.n497 dvss.n496 1.88285
R842 dvss.n458 dvss.n457 1.88285
R843 dvss.n419 dvss.n418 1.88285
R844 dvss.n37 dvss.n36 1.85983
R845 dvss.n23 dvss.n22 1.57196
R846 dvss.n29 dvss.n28 1.57139
R847 dvss.n187 dvss.n173 1.5505
R848 dvss.n69 dvss.n60 1.46336
R849 dvss.n525 dvss.n13 1.32907
R850 dvss.n120 dvss.n56 1.32907
R851 dvss.n410 dvss.n175 1.11858
R852 dvss.n192 dvss.n187 0.649775
R853 dvss dvss.n118 0.637219
R854 dvss.n380 dvss.n379 0.630008
R855 dvss.n394 dvss.n184 0.630008
R856 dvss.t180 dvss.n529 0.474702
R857 dvss.n529 dvss 0.36436
R858 dvss.n529 dvss.n528 0.357983
R859 dvss.n37 dvss 0.326572
R860 dvss.n534 dvss.n533 0.286958
R861 dvss.n99 dvss.n98 0.260009
R862 dvss.n166 dvss.t73 0.189075
R863 dvss.n73 dvss 0.178871
R864 dvss.n94 dvss.n90 0.178278
R865 dvss.n255 dvss 0.165648
R866 dvss.n533 dvss.n532 0.160391
R867 dvss.n528 dvss.n527 0.148545
R868 dvss.n71 dvss 0.145311
R869 dvss.n409 dvss 0.142307
R870 dvss.n98 dvss 0.140381
R871 dvss.n527 dvss.n10 0.136163
R872 dvss.n532 dvss.n531 0.13579
R873 dvss.n408 dvss.n407 0.120292
R874 dvss.n407 dvss.n176 0.120292
R875 dvss.n403 dvss.n176 0.120292
R876 dvss.n403 dvss.n402 0.120292
R877 dvss.n402 dvss.n401 0.120292
R878 dvss.n397 dvss.n396 0.120292
R879 dvss.n396 dvss.n395 0.120292
R880 dvss.n395 dvss.n182 0.120292
R881 dvss.n391 dvss.n182 0.120292
R882 dvss.n539 dvss.n538 0.120292
R883 dvss.n540 dvss.n539 0.120292
R884 dvss.n540 dvss.n4 0.120292
R885 dvss.n544 dvss.n4 0.120292
R886 dvss.n545 dvss.n544 0.120292
R887 dvss.n546 dvss.n545 0.120292
R888 dvss.n96 dvss 0.115052
R889 dvss.n118 dvss.n117 0.109875
R890 dvss.n74 dvss.n73 0.109468
R891 dvss.n410 dvss 0.0999624
R892 dvss.n538 dvss 0.0968542
R893 dvss.n99 dvss 0.0959969
R894 dvss.n77 dvss 0.080434
R895 dvss.n78 dvss.n77 0.0777204
R896 dvss.t72 dvss.t181 0.070611
R897 dvss.n49 dvss.n23 0.0678684
R898 dvss.n530 dvss.t180 0.0675999
R899 dvss.n47 dvss.n29 0.0671667
R900 dvss.n532 dvss.n8 0.0664942
R901 dvss dvss.n125 0.0652681
R902 dvss.n20 dvss 0.0633141
R903 dvss.n117 dvss.n56 0.0606266
R904 dvss.n528 dvss 0.060557
R905 dvss.n531 dvss.t73 0.060491
R906 dvss.n180 dvss 0.0603958
R907 dvss.n397 dvss 0.0603958
R908 dvss dvss.n390 0.0603958
R909 dvss.n535 dvss 0.0603958
R910 dvss.n71 dvss.n70 0.0603629
R911 dvss.n1 dvss 0.0525833
R912 dvss.n13 dvss.n10 0.0495635
R913 dvss.n106 dvss.n105 0.0482484
R914 dvss.n96 dvss.n95 0.0467134
R915 dvss.n28 dvss.n27 0.0457733
R916 dvss.n409 dvss.n408 0.0447708
R917 dvss.n117 dvss 0.0421667
R918 dvss.n530 dvss.n9 0.0405094
R919 dvss.n22 dvss 0.0346686
R920 dvss dvss.n534 0.0343542
R921 dvss dvss.n99 0.0335285
R922 dvss dvss.n180 0.0330521
R923 dvss.n390 dvss 0.0330521
R924 dvss.n10 dvss 0.0300195
R925 dvss.n73 dvss.n72 0.028566
R926 dvss.n102 dvss 0.0248902
R927 dvss.n535 dvss 0.0239375
R928 dvss.n27 dvss.n9 0.0228519
R929 dvss.n401 dvss 0.0226354
R930 dvss.n391 dvss 0.0226354
R931 dvss.n74 dvss 0.0215598
R932 dvss.n98 dvss.n97 0.0208358
R933 dvss.n118 dvss 0.0193397
R934 dvss.n21 dvss.n20 0.0184385
R935 dvss dvss.n59 0.0174837
R936 dvss.n516 dvss.n515 0.015957
R937 dvss.n515 dvss.n514 0.015957
R938 dvss.n514 dvss.n127 0.015957
R939 dvss.n510 dvss.n127 0.015957
R940 dvss.n510 dvss.n509 0.015957
R941 dvss.n509 dvss.n131 0.015957
R942 dvss.n505 dvss.n131 0.015957
R943 dvss.n505 dvss.n504 0.015957
R944 dvss.n504 dvss.n134 0.015957
R945 dvss.n500 dvss.n134 0.015957
R946 dvss.n500 dvss.n499 0.015957
R947 dvss.n499 dvss.n498 0.015957
R948 dvss.n498 dvss.n136 0.015957
R949 dvss.n493 dvss.n136 0.015957
R950 dvss.n493 dvss.n492 0.015957
R951 dvss.n492 dvss.n491 0.015957
R952 dvss.n491 dvss.n139 0.015957
R953 dvss.n487 dvss.n139 0.015957
R954 dvss.n487 dvss.n486 0.015957
R955 dvss.n486 dvss.n485 0.015957
R956 dvss.n485 dvss.n141 0.015957
R957 dvss.n481 dvss.n141 0.015957
R958 dvss.n479 dvss.n144 0.015957
R959 dvss.n474 dvss.n144 0.015957
R960 dvss.n474 dvss.n473 0.015957
R961 dvss.n473 dvss.n472 0.015957
R962 dvss.n472 dvss.n147 0.015957
R963 dvss.n467 dvss.n147 0.015957
R964 dvss.n467 dvss.n466 0.015957
R965 dvss.n466 dvss.n465 0.015957
R966 dvss.n465 dvss.n149 0.015957
R967 dvss.n461 dvss.n149 0.015957
R968 dvss.n461 dvss.n460 0.015957
R969 dvss.n460 dvss.n459 0.015957
R970 dvss.n459 dvss.n153 0.015957
R971 dvss.n454 dvss.n153 0.015957
R972 dvss.n454 dvss.n453 0.015957
R973 dvss.n453 dvss.n452 0.015957
R974 dvss.n452 dvss.n156 0.015957
R975 dvss.n448 dvss.n156 0.015957
R976 dvss.n448 dvss.n447 0.015957
R977 dvss.n447 dvss.n446 0.015957
R978 dvss.n446 dvss.n158 0.015957
R979 dvss.n442 dvss.n158 0.015957
R980 dvss.n440 dvss.n161 0.015957
R981 dvss.n435 dvss.n161 0.015957
R982 dvss.n435 dvss.n434 0.015957
R983 dvss.n434 dvss.n433 0.015957
R984 dvss.n433 dvss.n164 0.015957
R985 dvss.n428 dvss.n164 0.015957
R986 dvss.n428 dvss.n427 0.015957
R987 dvss.n427 dvss.n426 0.015957
R988 dvss.n423 dvss.n422 0.015957
R989 dvss.n422 dvss.n421 0.015957
R990 dvss.n421 dvss.n170 0.015957
R991 dvss.n416 dvss.n170 0.015957
R992 dvss.n416 dvss.n415 0.015957
R993 dvss.n415 dvss.n414 0.015957
R994 dvss.n410 dvss.n409 0.0141555
R995 dvss.n259 dvss.n254 0.0125293
R996 dvss.n260 dvss.n259 0.0125293
R997 dvss.n260 dvss.n251 0.0125293
R998 dvss.n265 dvss.n251 0.0125293
R999 dvss.n266 dvss.n265 0.0125293
R1000 dvss.n267 dvss.n266 0.0125293
R1001 dvss.n267 dvss.n248 0.0125293
R1002 dvss.n272 dvss.n248 0.0125293
R1003 dvss.n273 dvss.n272 0.0125293
R1004 dvss.n274 dvss.n273 0.0125293
R1005 dvss.n274 dvss.n246 0.0125293
R1006 dvss.n280 dvss.n246 0.0125293
R1007 dvss.n281 dvss.n280 0.0125293
R1008 dvss.n282 dvss.n281 0.0125293
R1009 dvss.n282 dvss.n244 0.0125293
R1010 dvss.n286 dvss.n244 0.0125293
R1011 dvss.n287 dvss.n286 0.0125293
R1012 dvss.n288 dvss.n287 0.0125293
R1013 dvss.n288 dvss.n242 0.0125293
R1014 dvss.n292 dvss.n242 0.0125293
R1015 dvss.n293 dvss.n292 0.0125293
R1016 dvss.n294 dvss.n293 0.0125293
R1017 dvss.n299 dvss.n237 0.0125293
R1018 dvss.n300 dvss.n299 0.0125293
R1019 dvss.n300 dvss.n234 0.0125293
R1020 dvss.n305 dvss.n234 0.0125293
R1021 dvss.n306 dvss.n305 0.0125293
R1022 dvss.n307 dvss.n306 0.0125293
R1023 dvss.n307 dvss.n231 0.0125293
R1024 dvss.n312 dvss.n231 0.0125293
R1025 dvss.n313 dvss.n312 0.0125293
R1026 dvss.n314 dvss.n313 0.0125293
R1027 dvss.n314 dvss.n229 0.0125293
R1028 dvss.n320 dvss.n229 0.0125293
R1029 dvss.n321 dvss.n320 0.0125293
R1030 dvss.n322 dvss.n321 0.0125293
R1031 dvss.n322 dvss.n227 0.0125293
R1032 dvss.n326 dvss.n227 0.0125293
R1033 dvss.n327 dvss.n326 0.0125293
R1034 dvss.n328 dvss.n327 0.0125293
R1035 dvss.n328 dvss.n225 0.0125293
R1036 dvss.n332 dvss.n225 0.0125293
R1037 dvss.n333 dvss.n332 0.0125293
R1038 dvss.n334 dvss.n333 0.0125293
R1039 dvss.n339 dvss.n219 0.0125293
R1040 dvss.n340 dvss.n339 0.0125293
R1041 dvss.n340 dvss.n216 0.0125293
R1042 dvss.n344 dvss.n216 0.0125293
R1043 dvss.n345 dvss.n344 0.0125293
R1044 dvss.n345 dvss.n214 0.0125293
R1045 dvss.n349 dvss.n214 0.0125293
R1046 dvss.n350 dvss.n349 0.0125293
R1047 dvss.n350 dvss.n211 0.0125293
R1048 dvss.n354 dvss.n211 0.0125293
R1049 dvss.n355 dvss.n354 0.0125293
R1050 dvss.n356 dvss.n355 0.0125293
R1051 dvss.n356 dvss.n208 0.0125293
R1052 dvss.n361 dvss.n208 0.0125293
R1053 dvss.n362 dvss.n361 0.0125293
R1054 dvss.n363 dvss.n362 0.0125293
R1055 dvss.n363 dvss.n206 0.0125293
R1056 dvss.n367 dvss.n206 0.0125293
R1057 dvss.n368 dvss.n367 0.0125293
R1058 dvss.n369 dvss.n368 0.0125293
R1059 dvss.n369 dvss.n203 0.0125293
R1060 dvss.n373 dvss.n203 0.0125293
R1061 dvss.n375 dvss.n201 0.0125293
R1062 dvss.n381 dvss.n201 0.0125293
R1063 dvss.n382 dvss.n381 0.0125293
R1064 dvss.n383 dvss.n382 0.0125293
R1065 dvss.n423 dvss.n166 0.0122608
R1066 dvss.n99 dvss 0.012146
R1067 dvss dvss.n21 0.0110353
R1068 dvss.n78 dvss.n74 0.0106902
R1069 dvss.n531 dvss.t72 0.0106199
R1070 dvss.n105 dvss 0.0105932
R1071 dvss.n411 dvss.n173 0.0099086
R1072 dvss.n546 dvss.n1 0.0083125
R1073 dvss.n516 dvss 0.00822849
R1074 dvss dvss.n480 0.00822849
R1075 dvss dvss.n479 0.00822849
R1076 dvss dvss.n441 0.00822849
R1077 dvss dvss.n440 0.00822849
R1078 dvss.n72 dvss.n71 0.00733962
R1079 dvss.n414 dvss.n173 0.00654839
R1080 dvss dvss.n254 0.00651464
R1081 dvss dvss.n238 0.00651464
R1082 dvss dvss.n237 0.00651464
R1083 dvss dvss.n220 0.00651464
R1084 dvss dvss.n219 0.00651464
R1085 dvss.n374 dvss 0.00651464
R1086 dvss.n375 dvss 0.00651464
R1087 dvss dvss.n199 0.00651464
R1088 dvss.n97 dvss.n96 0.00591045
R1089 dvss dvss.n1 0.00570833
R1090 dvss.n20 dvss.n9 0.00519818
R1091 dvss dvss.n125 0.00470027
R1092 dvss.n480 dvss 0.00470027
R1093 dvss.n441 dvss 0.00470027
R1094 dvss.n426 dvss.n166 0.00419624
R1095 dvss.n255 dvss 0.00376883
R1096 dvss.n238 dvss 0.00376883
R1097 dvss.n220 dvss 0.00376883
R1098 dvss dvss.n374 0.00376883
R1099 dvss.n199 dvss 0.00376883
R1100 dvss.t181 dvss.n530 0.00351108
R1101 dvss.n481 dvss 0.00335618
R1102 dvss.n442 dvss 0.00335618
R1103 dvss.n294 dvss 0.0027228
R1104 dvss.n334 dvss 0.0027228
R1105 dvss dvss.n373 0.0027228
R1106 dvss.n383 dvss 0.0027228
R1107 dvss.n411 dvss.n410 0.00150806
R1108 dvss.n70 dvss.n56 0.000763713
R1109 dvss.n95 dvss.n13 0.000703583
R1110 x7.x3.A2.n7 x7.x3.A2.t1 373.866
R1111 x7.x3.A2.n5 x7.x3.A2.t6 333.651
R1112 x7.x3.A2.n5 x7.x3.A2.t2 297.233
R1113 x7.x3.A2.n0 x7.x3.A2.t5 241.536
R1114 x7.x3.A2 x7.x3.A2.t0 237.101
R1115 x7.x3.A2.n3 x7.x3.A2.t3 207.423
R1116 x7.x3.A2.n2 x7.x3.A2.t4 202.133
R1117 x7.x3.A2 x7.x3.A2.n5 195.701
R1118 x7.x3.A2.n0 x7.x3.A2.t7 169.237
R1119 x7.x3.A2.n4 x7.x3.A2.n3 159.758
R1120 x7.x3.A2.n2 x7.x3.A2 154.91
R1121 x7.x3.A2.n1 x7.x3.A2.n0 152
R1122 x7.x3.A2.n3 x7.x3.A2.n2 36.8275
R1123 x7.x3.A2 x7.x3.A2.n7 26.7478
R1124 x7.x3.A2.n6 x7.x3.A2 15.8995
R1125 x7.x3.A2.n6 x7.x3.A2 15.7806
R1126 x7.x3.A2 x7.x3.A2.n1 14.8117
R1127 x7.x3.A2 x7.x3.A2.n4 13.8784
R1128 x7.x3.A2.n7 x7.x3.A2.n6 3.1005
R1129 x7.x3.A2.n4 x7.x3.A2 2.52171
R1130 x7.x3.A2.n1 x7.x3.A2 1.9205
R1131 dvdd.n294 dvdd.n285 5128.23
R1132 dvdd.n294 dvdd.n286 5128.23
R1133 dvdd.n292 dvdd.n286 5128.23
R1134 dvdd.n292 dvdd.n285 5128.23
R1135 dvdd.n42 dvdd.n5 1736.47
R1136 dvdd.n45 dvdd.n4 1736.47
R1137 dvdd.n30 dvdd.n27 1736.47
R1138 dvdd.n33 dvdd.n29 1736.47
R1139 dvdd.n254 dvdd.t142 838.817
R1140 dvdd.n67 dvdd.t170 806.511
R1141 dvdd.n67 dvdd.t122 806.511
R1142 dvdd.n88 dvdd.t107 806.511
R1143 dvdd.n88 dvdd.t80 806.511
R1144 dvdd.n109 dvdd.t128 806.511
R1145 dvdd.n109 dvdd.t7 806.511
R1146 dvdd.n291 dvdd.n283 787.447
R1147 dvdd.n291 dvdd.n284 786.827
R1148 dvdd.n56 dvdd.t53 668.683
R1149 dvdd.n56 dvdd.t118 668.683
R1150 dvdd.n225 dvdd.t163 667.778
R1151 dvdd.n225 dvdd.t124 667.778
R1152 dvdd.n187 dvdd.t69 667.778
R1153 dvdd.n187 dvdd.t160 667.778
R1154 dvdd.n149 dvdd.t99 667.778
R1155 dvdd.n149 dvdd.t15 667.778
R1156 dvdd.n295 dvdd.n283 604.574
R1157 dvdd.n71 dvdd.n69 604.457
R1158 dvdd.n71 dvdd.n70 604.457
R1159 dvdd.n92 dvdd.n90 604.457
R1160 dvdd.n92 dvdd.n91 604.457
R1161 dvdd.n113 dvdd.n111 604.457
R1162 dvdd.n113 dvdd.n112 604.457
R1163 dvdd.n230 dvdd.n59 604.394
R1164 dvdd.n230 dvdd.n60 604.394
R1165 dvdd.n192 dvdd.n80 604.394
R1166 dvdd.n192 dvdd.n81 604.394
R1167 dvdd.n154 dvdd.n101 604.394
R1168 dvdd.n154 dvdd.n102 604.394
R1169 dvdd.n218 dvdd.n65 601.679
R1170 dvdd.n218 dvdd.n66 601.679
R1171 dvdd.n180 dvdd.n86 601.679
R1172 dvdd.n180 dvdd.n87 601.679
R1173 dvdd.n142 dvdd.n107 601.679
R1174 dvdd.n142 dvdd.n108 601.679
R1175 dvdd.n259 dvdd.n258 585
R1176 dvdd.t158 dvdd.t141 556.386
R1177 dvdd.n245 dvdd 538.664
R1178 dvdd.n18 dvdd 535.705
R1179 dvdd.n11 dvdd 535.705
R1180 dvdd.t130 dvdd 473.521
R1181 dvdd.t14 dvdd.t145 448.146
R1182 dvdd.t68 dvdd.t20 448.146
R1183 dvdd.t123 dvdd.t24 448.146
R1184 dvdd.n295 dvdd.n284 423.062
R1185 dvdd.t132 dvdd.t56 367.579
R1186 dvdd.t48 dvdd.t84 367.579
R1187 dvdd.t2 dvdd.t101 367.579
R1188 dvdd.n273 dvdd.t16 360.005
R1189 dvdd.t6 dvdd.t134 330.654
R1190 dvdd.t79 dvdd.t111 330.654
R1191 dvdd.t121 dvdd.t91 330.654
R1192 dvdd.n43 dvdd.n4 314.781
R1193 dvdd.n44 dvdd.n5 314.781
R1194 dvdd.n31 dvdd.n29 314.781
R1195 dvdd.n32 dvdd.n27 314.781
R1196 dvdd.n23 dvdd.n17 312.053
R1197 dvdd.n9 dvdd.n8 312.051
R1198 dvdd.n265 dvdd.n255 312.051
R1199 dvdd.t39 dvdd.t37 304.829
R1200 dvdd.t141 dvdd.t10 284.113
R1201 dvdd.t56 dvdd.t50 275.265
R1202 dvdd.t84 dvdd.t63 275.265
R1203 dvdd.t101 dvdd.t8 275.265
R1204 dvdd.t10 dvdd.t130 275.235
R1205 dvdd.n270 dvdd.t82 261.837
R1206 dvdd.t32 dvdd.t137 260.437
R1207 dvdd.t147 dvdd.t41 260.437
R1208 dvdd.n205 dvdd.n74 259.707
R1209 dvdd.n205 dvdd.n73 259.707
R1210 dvdd.n167 dvdd.n95 259.707
R1211 dvdd.n167 dvdd.n94 259.707
R1212 dvdd.n129 dvdd.n116 259.707
R1213 dvdd.n129 dvdd.n115 259.707
R1214 dvdd.t82 dvdd.t12 258.481
R1215 dvdd.n272 dvdd.t108 253.446
R1216 dvdd.n271 dvdd.t4 253.446
R1217 dvdd.t19 dvdd.t98 248.599
R1218 dvdd.t98 dvdd.t158 248.599
R1219 dvdd.n199 dvdd.n78 242.607
R1220 dvdd.n161 dvdd.n99 242.607
R1221 dvdd.n123 dvdd.n121 242.607
R1222 dvdd.n199 dvdd.n77 242.607
R1223 dvdd.n161 dvdd.n98 242.607
R1224 dvdd.n123 dvdd.n120 242.607
R1225 dvdd.t0 dvdd.t103 234.982
R1226 dvdd.t60 dvdd.t36 234.982
R1227 dvdd.t43 dvdd.t89 234.982
R1228 dvdd dvdd.n269 232.445
R1229 dvdd.n0 dvdd.t114 228.215
R1230 dvdd.n0 dvdd.t126 228.215
R1231 dvdd.n238 dvdd.n236 215.123
R1232 dvdd.n238 dvdd.n237 215.123
R1233 dvdd.t37 dvdd.t62 213.084
R1234 dvdd.n41 dvdd.n3 185.225
R1235 dvdd.n46 dvdd.n3 185.225
R1236 dvdd.n34 dvdd.n28 185.225
R1237 dvdd.n28 dvdd.n26 185.225
R1238 dvdd.t30 dvdd.t54 181.273
R1239 dvdd.t94 dvdd.t86 181.273
R1240 dvdd.t65 dvdd.t58 181.273
R1241 dvdd.t144 dvdd.t6 166.167
R1242 dvdd.t103 dvdd.t105 166.167
R1243 dvdd.t34 dvdd.t79 166.167
R1244 dvdd.t36 dvdd.t18 166.167
R1245 dvdd.t104 dvdd.t121 166.167
R1246 dvdd.t89 dvdd.t136 166.167
R1247 dvdd.t16 dvdd.t132 162.81
R1248 dvdd.t134 dvdd.t0 162.81
R1249 dvdd.t108 dvdd.t48 162.81
R1250 dvdd.t111 dvdd.t60 162.81
R1251 dvdd.t4 dvdd.t2 162.81
R1252 dvdd.t91 dvdd.t43 162.81
R1253 dvdd.t70 dvdd.n292 161.316
R1254 dvdd.n294 dvdd.t164 161.316
R1255 dvdd.t105 dvdd.t14 154.417
R1256 dvdd.t18 dvdd.t68 154.417
R1257 dvdd.t136 dvdd.t123 154.417
R1258 dvdd.t12 dvdd.t52 147.703
R1259 dvdd.n73 dvdd.t9 147.111
R1260 dvdd.n74 dvdd.t173 147.111
R1261 dvdd.n94 dvdd.t156 147.111
R1262 dvdd.n95 dvdd.t64 147.111
R1263 dvdd.n115 dvdd.t159 147.111
R1264 dvdd.n116 dvdd.t51 147.111
R1265 dvdd.t106 dvdd.t144 144.346
R1266 dvdd.t45 dvdd.t34 144.346
R1267 dvdd.t26 dvdd.t104 144.346
R1268 dvdd.t50 dvdd.t30 140.989
R1269 dvdd.t54 dvdd.t106 140.989
R1270 dvdd.t145 dvdd.t119 140.989
R1271 dvdd.t63 dvdd.t94 140.989
R1272 dvdd.t86 dvdd.t45 140.989
R1273 dvdd.t20 dvdd.t46 140.989
R1274 dvdd.t8 dvdd.t65 140.989
R1275 dvdd.t58 dvdd.t26 140.989
R1276 dvdd.t24 dvdd.t28 140.989
R1277 dvdd.t52 dvdd 132.597
R1278 dvdd dvdd.n272 125.883
R1279 dvdd dvdd.n271 125.883
R1280 dvdd dvdd.n270 125.883
R1281 dvdd.t77 dvdd.t70 121.245
R1282 dvdd.t75 dvdd.t77 121.245
R1283 dvdd.t96 dvdd.t75 121.245
R1284 dvdd.t161 dvdd.t96 121.245
R1285 dvdd.t73 dvdd.t166 121.245
R1286 dvdd.t115 dvdd.t73 121.245
R1287 dvdd.t22 dvdd.t115 121.245
R1288 dvdd.t164 dvdd.t22 121.245
R1289 dvdd.n69 dvdd.t72 119.608
R1290 dvdd.n70 dvdd.t59 119.608
R1291 dvdd.n90 dvdd.t153 119.608
R1292 dvdd.n91 dvdd.t87 119.608
R1293 dvdd.n111 dvdd.t55 119.608
R1294 dvdd.n112 dvdd.t157 119.608
R1295 dvdd.t119 dvdd 109.1
R1296 dvdd.t46 dvdd 109.1
R1297 dvdd.t28 dvdd 109.1
R1298 dvdd.n73 dvdd.t102 108.413
R1299 dvdd.n74 dvdd.t140 108.413
R1300 dvdd.n94 dvdd.t171 108.413
R1301 dvdd.n95 dvdd.t85 108.413
R1302 dvdd.n115 dvdd.t57 108.413
R1303 dvdd.n116 dvdd.t154 108.413
R1304 dvdd.n270 dvdd.n55 106.559
R1305 dvdd.n271 dvdd.n54 106.559
R1306 dvdd.n272 dvdd.n53 106.559
R1307 dvdd.n47 dvdd.n2 105.412
R1308 dvdd.n40 dvdd.n2 105.412
R1309 dvdd.n37 dvdd.n36 105.412
R1310 dvdd.n36 dvdd.n35 105.412
R1311 dvdd dvdd.t39 100.624
R1312 dvdd.n65 dvdd.t44 93.81
R1313 dvdd.n66 dvdd.t67 93.81
R1314 dvdd.n86 dvdd.t168 93.81
R1315 dvdd.n87 dvdd.t61 93.81
R1316 dvdd.n107 dvdd.t174 93.81
R1317 dvdd.n108 dvdd.t1 93.81
R1318 dvdd dvdd.t32 91.745
R1319 dvdd dvdd.t147 91.745
R1320 dvdd dvdd.t19 88.7855
R1321 dvdd.n258 dvdd.t40 86.7743
R1322 dvdd.n47 dvdd.n46 79.8123
R1323 dvdd.n41 dvdd.n40 79.8123
R1324 dvdd.n35 dvdd.n34 79.8123
R1325 dvdd.n37 dvdd.n26 79.8123
R1326 dvdd.n236 dvdd.t100 74.7554
R1327 dvdd.n237 dvdd.t13 74.7554
R1328 dvdd.n65 dvdd.t92 63.3219
R1329 dvdd.n66 dvdd.t93 63.3219
R1330 dvdd.n69 dvdd.t90 63.3219
R1331 dvdd.n70 dvdd.t66 63.3219
R1332 dvdd.n86 dvdd.t112 63.3219
R1333 dvdd.n87 dvdd.t143 63.3219
R1334 dvdd.n90 dvdd.t150 63.3219
R1335 dvdd.n91 dvdd.t95 63.3219
R1336 dvdd.n107 dvdd.t135 63.3219
R1337 dvdd.n108 dvdd.t139 63.3219
R1338 dvdd.n111 dvdd.t110 63.3219
R1339 dvdd.n112 dvdd.t31 63.3219
R1340 dvdd.n77 dvdd.t27 61.9829
R1341 dvdd.n98 dvdd.t49 61.9829
R1342 dvdd.n120 dvdd.t151 61.9829
R1343 dvdd.n78 dvdd.t3 61.9826
R1344 dvdd.n99 dvdd.t88 61.9826
R1345 dvdd.n121 dvdd.t133 61.9826
R1346 dvdd.n258 dvdd.t38 61.05
R1347 dvdd.n293 dvdd.t161 60.6225
R1348 dvdd.t166 dvdd.n293 60.6225
R1349 dvdd.n291 dvdd.t71 60.3236
R1350 dvdd.n295 dvdd.t165 60.3236
R1351 dvdd.n296 dvdd.n282 54.7085
R1352 dvdd.n297 dvdd.n281 54.7085
R1353 dvdd.n289 dvdd.n288 54.7085
R1354 dvdd.n290 dvdd.n287 54.7085
R1355 dvdd.n59 dvdd.t155 41.5552
R1356 dvdd.n59 dvdd.t127 41.5552
R1357 dvdd.n60 dvdd.t25 41.5552
R1358 dvdd.n60 dvdd.t29 41.5552
R1359 dvdd.n80 dvdd.t129 41.5552
R1360 dvdd.n80 dvdd.t81 41.5552
R1361 dvdd.n81 dvdd.t21 41.5552
R1362 dvdd.n81 dvdd.t47 41.5552
R1363 dvdd.n101 dvdd.t146 41.5552
R1364 dvdd.n101 dvdd.t169 41.5552
R1365 dvdd.n102 dvdd.t172 41.5552
R1366 dvdd.n102 dvdd.t120 41.5552
R1367 dvdd.n46 dvdd.n45 37.0005
R1368 dvdd.n42 dvdd.n41 37.0005
R1369 dvdd.n34 dvdd.n33 37.0005
R1370 dvdd.n30 dvdd.n26 37.0005
R1371 dvdd.n17 dvdd.t33 36.1587
R1372 dvdd.n17 dvdd.t138 36.1587
R1373 dvdd.n8 dvdd.t148 36.1587
R1374 dvdd.n8 dvdd.t42 36.1587
R1375 dvdd.n255 dvdd.t11 35.4605
R1376 dvdd.n249 dvdd.n248 34.6358
R1377 dvdd.n253 dvdd.n244 34.6358
R1378 dvdd.n264 dvdd.n256 34.6358
R1379 dvdd.n229 dvdd.n61 34.6358
R1380 dvdd.n219 dvdd.n63 34.6358
R1381 dvdd.n223 dvdd.n63 34.6358
R1382 dvdd.n224 dvdd.n223 34.6358
R1383 dvdd.n217 dvdd.n216 34.6358
R1384 dvdd.n211 dvdd.n210 34.6358
R1385 dvdd.n212 dvdd.n211 34.6358
R1386 dvdd.n198 dvdd.n197 34.6358
R1387 dvdd.n200 dvdd.n75 34.6358
R1388 dvdd.n204 dvdd.n75 34.6358
R1389 dvdd.n191 dvdd.n82 34.6358
R1390 dvdd.n181 dvdd.n84 34.6358
R1391 dvdd.n185 dvdd.n84 34.6358
R1392 dvdd.n186 dvdd.n185 34.6358
R1393 dvdd.n179 dvdd.n178 34.6358
R1394 dvdd.n173 dvdd.n172 34.6358
R1395 dvdd.n174 dvdd.n173 34.6358
R1396 dvdd.n160 dvdd.n159 34.6358
R1397 dvdd.n162 dvdd.n96 34.6358
R1398 dvdd.n166 dvdd.n96 34.6358
R1399 dvdd.n153 dvdd.n103 34.6358
R1400 dvdd.n143 dvdd.n105 34.6358
R1401 dvdd.n147 dvdd.n105 34.6358
R1402 dvdd.n148 dvdd.n147 34.6358
R1403 dvdd.n141 dvdd.n140 34.6358
R1404 dvdd.n135 dvdd.n134 34.6358
R1405 dvdd.n136 dvdd.n135 34.6358
R1406 dvdd.n122 dvdd.n52 34.6358
R1407 dvdd.n124 dvdd.n117 34.6358
R1408 dvdd.n128 dvdd.n117 34.6358
R1409 dvdd.n238 dvdd.n235 33.8829
R1410 dvdd.n225 dvdd.n224 32.377
R1411 dvdd.n187 dvdd.n186 32.377
R1412 dvdd.n149 dvdd.n148 32.377
R1413 dvdd.n212 dvdd.n67 32.0005
R1414 dvdd.n174 dvdd.n88 32.0005
R1415 dvdd.n136 dvdd.n109 32.0005
R1416 dvdd.n239 dvdd.n238 31.624
R1417 dvdd.n200 dvdd.n199 31.2476
R1418 dvdd.n162 dvdd.n161 31.2476
R1419 dvdd.n124 dvdd.n123 31.2476
R1420 dvdd.n5 dvdd.n3 30.8338
R1421 dvdd.n4 dvdd.n2 30.8338
R1422 dvdd.n36 dvdd.n27 30.8338
R1423 dvdd.n29 dvdd.n28 30.8338
R1424 dvdd.n77 dvdd.t5 30.1745
R1425 dvdd.n98 dvdd.t149 30.1745
R1426 dvdd.n120 dvdd.t17 30.1745
R1427 dvdd.n78 dvdd.t35 30.1738
R1428 dvdd.n99 dvdd.t109 30.1738
R1429 dvdd.n121 dvdd.t117 30.1738
R1430 dvdd.n206 dvdd.n71 30.1181
R1431 dvdd.n168 dvdd.n92 30.1181
R1432 dvdd.n130 dvdd.n113 30.1181
R1433 dvdd.n43 dvdd.n42 29.6618
R1434 dvdd.n45 dvdd.n44 29.6618
R1435 dvdd.n31 dvdd.n30 29.6618
R1436 dvdd.n33 dvdd.n32 29.6618
R1437 dvdd.n236 dvdd.t83 28.5349
R1438 dvdd.n237 dvdd.t152 28.5349
R1439 dvdd.n260 dvdd.n256 28.2952
R1440 dvdd dvdd.n244 27.8593
R1441 dvdd.n255 dvdd.t131 26.5955
R1442 dvdd.n259 dvdd.n257 25.2079
R1443 dvdd.n22 dvdd.n18 23.7181
R1444 dvdd.n11 dvdd.n10 23.7181
R1445 dvdd.n248 dvdd.n245 23.7181
R1446 dvdd.n231 dvdd.n55 23.7181
R1447 dvdd.n197 dvdd.n54 23.7181
R1448 dvdd.n193 dvdd.n54 23.7181
R1449 dvdd.n159 dvdd.n53 23.7181
R1450 dvdd.n155 dvdd.n53 23.7181
R1451 dvdd.n273 dvdd.n52 23.7181
R1452 dvdd.n235 dvdd.n55 23.7181
R1453 dvdd.n230 dvdd.n229 22.9652
R1454 dvdd.n192 dvdd.n191 22.9652
R1455 dvdd.n154 dvdd.n153 22.9652
R1456 dvdd.n266 dvdd.n254 22.5887
R1457 dvdd.n265 dvdd.n264 22.5887
R1458 dvdd.n266 dvdd.n265 21.8358
R1459 dvdd.n231 dvdd.n230 21.4593
R1460 dvdd.n193 dvdd.n192 21.4593
R1461 dvdd.n155 dvdd.n154 21.4593
R1462 dvdd.n210 dvdd.n71 20.3299
R1463 dvdd.n172 dvdd.n92 20.3299
R1464 dvdd.n134 dvdd.n113 20.3299
R1465 dvdd.n254 dvdd.n253 19.9534
R1466 dvdd.n239 dvdd.n56 19.577
R1467 dvdd.n269 dvdd.n56 18.4476
R1468 dvdd.n225 dvdd.n61 18.0711
R1469 dvdd.n187 dvdd.n82 18.0711
R1470 dvdd.n149 dvdd.n103 18.0711
R1471 dvdd.n23 dvdd 15.8123
R1472 dvdd dvdd.n9 15.8123
R1473 dvdd.n295 dvdd.n294 13.2148
R1474 dvdd.n292 dvdd.n291 13.2148
R1475 dvdd.n38 dvdd.n37 10.0436
R1476 dvdd.n35 dvdd.n1 9.59217
R1477 dvdd.n216 dvdd.n67 9.41227
R1478 dvdd.n178 dvdd.n88 9.41227
R1479 dvdd.n140 dvdd.n109 9.41227
R1480 dvdd.n19 dvdd.n18 9.3005
R1481 dvdd.n22 dvdd.n21 9.3005
R1482 dvdd.n10 dvdd.n6 9.3005
R1483 dvdd.n12 dvdd.n11 9.3005
R1484 dvdd.n40 dvdd.n39 9.3005
R1485 dvdd.n48 dvdd.n47 9.3005
R1486 dvdd.n261 dvdd.n260 9.3005
R1487 dvdd.n262 dvdd.n256 9.3005
R1488 dvdd.n264 dvdd.n263 9.3005
R1489 dvdd.n265 dvdd.n242 9.3005
R1490 dvdd.n254 dvdd.n243 9.3005
R1491 dvdd.n253 dvdd.n252 9.3005
R1492 dvdd.n251 dvdd.n244 9.3005
R1493 dvdd.n250 dvdd.n249 9.3005
R1494 dvdd.n248 dvdd.n247 9.3005
R1495 dvdd.n246 dvdd.n245 9.3005
R1496 dvdd.n269 dvdd.n268 9.3005
R1497 dvdd.n274 dvdd.n273 9.3005
R1498 dvdd.n118 dvdd.n52 9.3005
R1499 dvdd.n122 dvdd.n119 9.3005
R1500 dvdd.n125 dvdd.n124 9.3005
R1501 dvdd.n126 dvdd.n117 9.3005
R1502 dvdd.n128 dvdd.n127 9.3005
R1503 dvdd.n129 dvdd.n114 9.3005
R1504 dvdd.n131 dvdd.n130 9.3005
R1505 dvdd.n132 dvdd.n113 9.3005
R1506 dvdd.n134 dvdd.n133 9.3005
R1507 dvdd.n135 dvdd.n110 9.3005
R1508 dvdd.n137 dvdd.n136 9.3005
R1509 dvdd.n138 dvdd.n109 9.3005
R1510 dvdd.n140 dvdd.n139 9.3005
R1511 dvdd.n141 dvdd.n106 9.3005
R1512 dvdd.n144 dvdd.n143 9.3005
R1513 dvdd.n145 dvdd.n105 9.3005
R1514 dvdd.n147 dvdd.n146 9.3005
R1515 dvdd.n148 dvdd.n104 9.3005
R1516 dvdd.n150 dvdd.n149 9.3005
R1517 dvdd.n151 dvdd.n103 9.3005
R1518 dvdd.n153 dvdd.n152 9.3005
R1519 dvdd.n154 dvdd.n100 9.3005
R1520 dvdd.n156 dvdd.n155 9.3005
R1521 dvdd.n157 dvdd.n53 9.3005
R1522 dvdd.n159 dvdd.n158 9.3005
R1523 dvdd.n160 dvdd.n97 9.3005
R1524 dvdd.n163 dvdd.n162 9.3005
R1525 dvdd.n164 dvdd.n96 9.3005
R1526 dvdd.n166 dvdd.n165 9.3005
R1527 dvdd.n167 dvdd.n93 9.3005
R1528 dvdd.n169 dvdd.n168 9.3005
R1529 dvdd.n170 dvdd.n92 9.3005
R1530 dvdd.n172 dvdd.n171 9.3005
R1531 dvdd.n173 dvdd.n89 9.3005
R1532 dvdd.n175 dvdd.n174 9.3005
R1533 dvdd.n176 dvdd.n88 9.3005
R1534 dvdd.n178 dvdd.n177 9.3005
R1535 dvdd.n179 dvdd.n85 9.3005
R1536 dvdd.n182 dvdd.n181 9.3005
R1537 dvdd.n183 dvdd.n84 9.3005
R1538 dvdd.n185 dvdd.n184 9.3005
R1539 dvdd.n186 dvdd.n83 9.3005
R1540 dvdd.n188 dvdd.n187 9.3005
R1541 dvdd.n189 dvdd.n82 9.3005
R1542 dvdd.n191 dvdd.n190 9.3005
R1543 dvdd.n192 dvdd.n79 9.3005
R1544 dvdd.n194 dvdd.n193 9.3005
R1545 dvdd.n195 dvdd.n54 9.3005
R1546 dvdd.n197 dvdd.n196 9.3005
R1547 dvdd.n198 dvdd.n76 9.3005
R1548 dvdd.n201 dvdd.n200 9.3005
R1549 dvdd.n202 dvdd.n75 9.3005
R1550 dvdd.n204 dvdd.n203 9.3005
R1551 dvdd.n205 dvdd.n72 9.3005
R1552 dvdd.n207 dvdd.n206 9.3005
R1553 dvdd.n208 dvdd.n71 9.3005
R1554 dvdd.n210 dvdd.n209 9.3005
R1555 dvdd.n211 dvdd.n68 9.3005
R1556 dvdd.n213 dvdd.n212 9.3005
R1557 dvdd.n214 dvdd.n67 9.3005
R1558 dvdd.n216 dvdd.n215 9.3005
R1559 dvdd.n217 dvdd.n64 9.3005
R1560 dvdd.n220 dvdd.n219 9.3005
R1561 dvdd.n221 dvdd.n63 9.3005
R1562 dvdd.n223 dvdd.n222 9.3005
R1563 dvdd.n224 dvdd.n62 9.3005
R1564 dvdd.n226 dvdd.n225 9.3005
R1565 dvdd.n227 dvdd.n61 9.3005
R1566 dvdd.n229 dvdd.n228 9.3005
R1567 dvdd.n230 dvdd.n58 9.3005
R1568 dvdd.n232 dvdd.n231 9.3005
R1569 dvdd.n233 dvdd.n55 9.3005
R1570 dvdd.n235 dvdd.n234 9.3005
R1571 dvdd.n240 dvdd.n239 9.3005
R1572 dvdd.n241 dvdd.n56 9.3005
R1573 dvdd.n267 dvdd.n266 9.3005
R1574 dvdd.n206 dvdd.n205 9.03579
R1575 dvdd.n168 dvdd.n167 9.03579
R1576 dvdd.n130 dvdd.n129 9.03579
R1577 dvdd.n285 dvdd.n283 7.70883
R1578 dvdd.n293 dvdd.n285 7.70883
R1579 dvdd.n286 dvdd.n284 7.70883
R1580 dvdd.n293 dvdd.n286 7.70883
R1581 dvdd.n24 dvdd.n23 7.17001
R1582 dvdd.n9 dvdd.n7 7.15376
R1583 dvdd.n282 dvdd.t116 7.14175
R1584 dvdd.n282 dvdd.t23 7.14175
R1585 dvdd.n281 dvdd.t167 7.14175
R1586 dvdd.n281 dvdd.t74 7.14175
R1587 dvdd.n288 dvdd.t97 7.14175
R1588 dvdd.n288 dvdd.t162 7.14175
R1589 dvdd.n287 dvdd.t78 7.14175
R1590 dvdd.n287 dvdd.t76 7.14175
R1591 dvdd.n249 dvdd 6.77697
R1592 dvdd.n44 dvdd.t125 6.70818
R1593 dvdd.t125 dvdd.n43 6.70818
R1594 dvdd.n32 dvdd.t113 6.70818
R1595 dvdd.t113 dvdd.n31 6.70818
R1596 dvdd dvdd.n22 6.4005
R1597 dvdd.n10 dvdd 6.4005
R1598 dvdd.n219 dvdd.n218 6.02403
R1599 dvdd.n205 dvdd.n204 6.02403
R1600 dvdd.n181 dvdd.n180 6.02403
R1601 dvdd.n167 dvdd.n166 6.02403
R1602 dvdd.n143 dvdd.n142 6.02403
R1603 dvdd.n129 dvdd.n128 6.02403
R1604 dvdd.n238 dvdd.n57 4.62124
R1605 dvdd.n218 dvdd.n217 3.76521
R1606 dvdd.n180 dvdd.n179 3.76521
R1607 dvdd.n142 dvdd.n141 3.76521
R1608 dvdd.n199 dvdd.n198 3.38874
R1609 dvdd.n161 dvdd.n160 3.38874
R1610 dvdd.n123 dvdd.n122 3.38874
R1611 dvdd.n296 dvdd.n295 1.66909
R1612 dvdd.n275 dvdd.n274 1.6403
R1613 dvdd.n291 dvdd.n290 1.57188
R1614 dvdd.n246 dvdd.n51 1.3879
R1615 dvdd.n36 dvdd.n0 1.32907
R1616 dvdd.n2 dvdd.n0 1.32907
R1617 dvdd.n260 dvdd.n259 1.23559
R1618 dvdd.n51 dvdd 0.694944
R1619 dvdd dvdd.n267 0.438
R1620 dvdd.n50 dvdd.n49 0.432317
R1621 dvdd.n16 dvdd 0.42713
R1622 dvdd dvdd.n16 0.32387
R1623 dvdd.n267 dvdd 0.313
R1624 dvdd.n275 dvdd.n51 0.252941
R1625 dvdd.n7 dvdd 0.203706
R1626 dvdd.n234 dvdd.n57 0.180304
R1627 dvdd.n240 dvdd.n57 0.180304
R1628 dvdd.n13 dvdd 0.167167
R1629 dvdd.n19 dvdd 0.164848
R1630 dvdd.n257 dvdd 0.159538
R1631 dvdd.n38 dvdd.n15 0.141704
R1632 dvdd.n261 dvdd.n257 0.141672
R1633 dvdd.n38 dvdd.n25 0.139389
R1634 dvdd.n14 dvdd.n6 0.127236
R1635 dvdd.n263 dvdd.n242 0.120292
R1636 dvdd.n251 dvdd.n250 0.120292
R1637 dvdd.n252 dvdd.n251 0.120292
R1638 dvdd.n252 dvdd.n243 0.120292
R1639 dvdd.n119 dvdd.n118 0.120292
R1640 dvdd.n125 dvdd.n119 0.120292
R1641 dvdd.n126 dvdd.n125 0.120292
R1642 dvdd.n127 dvdd.n126 0.120292
R1643 dvdd.n127 dvdd.n114 0.120292
R1644 dvdd.n131 dvdd.n114 0.120292
R1645 dvdd.n132 dvdd.n131 0.120292
R1646 dvdd.n133 dvdd.n132 0.120292
R1647 dvdd.n133 dvdd.n110 0.120292
R1648 dvdd.n137 dvdd.n110 0.120292
R1649 dvdd.n138 dvdd.n137 0.120292
R1650 dvdd.n139 dvdd.n138 0.120292
R1651 dvdd.n139 dvdd.n106 0.120292
R1652 dvdd.n144 dvdd.n106 0.120292
R1653 dvdd.n145 dvdd.n144 0.120292
R1654 dvdd.n146 dvdd.n145 0.120292
R1655 dvdd.n146 dvdd.n104 0.120292
R1656 dvdd.n150 dvdd.n104 0.120292
R1657 dvdd.n151 dvdd.n150 0.120292
R1658 dvdd.n152 dvdd.n151 0.120292
R1659 dvdd.n152 dvdd.n100 0.120292
R1660 dvdd.n156 dvdd.n100 0.120292
R1661 dvdd.n158 dvdd.n97 0.120292
R1662 dvdd.n163 dvdd.n97 0.120292
R1663 dvdd.n164 dvdd.n163 0.120292
R1664 dvdd.n165 dvdd.n164 0.120292
R1665 dvdd.n165 dvdd.n93 0.120292
R1666 dvdd.n169 dvdd.n93 0.120292
R1667 dvdd.n170 dvdd.n169 0.120292
R1668 dvdd.n171 dvdd.n170 0.120292
R1669 dvdd.n171 dvdd.n89 0.120292
R1670 dvdd.n175 dvdd.n89 0.120292
R1671 dvdd.n176 dvdd.n175 0.120292
R1672 dvdd.n177 dvdd.n176 0.120292
R1673 dvdd.n177 dvdd.n85 0.120292
R1674 dvdd.n182 dvdd.n85 0.120292
R1675 dvdd.n183 dvdd.n182 0.120292
R1676 dvdd.n184 dvdd.n183 0.120292
R1677 dvdd.n184 dvdd.n83 0.120292
R1678 dvdd.n188 dvdd.n83 0.120292
R1679 dvdd.n189 dvdd.n188 0.120292
R1680 dvdd.n190 dvdd.n189 0.120292
R1681 dvdd.n190 dvdd.n79 0.120292
R1682 dvdd.n194 dvdd.n79 0.120292
R1683 dvdd.n196 dvdd.n76 0.120292
R1684 dvdd.n201 dvdd.n76 0.120292
R1685 dvdd.n202 dvdd.n201 0.120292
R1686 dvdd.n203 dvdd.n202 0.120292
R1687 dvdd.n203 dvdd.n72 0.120292
R1688 dvdd.n207 dvdd.n72 0.120292
R1689 dvdd.n208 dvdd.n207 0.120292
R1690 dvdd.n209 dvdd.n208 0.120292
R1691 dvdd.n209 dvdd.n68 0.120292
R1692 dvdd.n213 dvdd.n68 0.120292
R1693 dvdd.n214 dvdd.n213 0.120292
R1694 dvdd.n215 dvdd.n214 0.120292
R1695 dvdd.n215 dvdd.n64 0.120292
R1696 dvdd.n220 dvdd.n64 0.120292
R1697 dvdd.n221 dvdd.n220 0.120292
R1698 dvdd.n222 dvdd.n221 0.120292
R1699 dvdd.n222 dvdd.n62 0.120292
R1700 dvdd.n226 dvdd.n62 0.120292
R1701 dvdd.n227 dvdd.n226 0.120292
R1702 dvdd.n228 dvdd.n227 0.120292
R1703 dvdd.n228 dvdd.n58 0.120292
R1704 dvdd.n232 dvdd.n58 0.120292
R1705 dvdd.n241 dvdd.n240 0.120292
R1706 dvdd.n276 dvdd.n275 0.109494
R1707 dvdd.n15 dvdd.n14 0.109053
R1708 dvdd.n267 dvdd.n243 0.107271
R1709 dvdd.n14 dvdd 0.0983618
R1710 dvdd dvdd.n261 0.0981562
R1711 dvdd.n250 dvdd 0.0968542
R1712 dvdd.n280 dvdd.n279 0.0944312
R1713 dvdd.n277 dvdd.n276 0.0856755
R1714 dvdd.n278 dvdd.n277 0.0856755
R1715 dvdd dvdd.n6 0.0803611
R1716 dvdd.n279 dvdd.n278 0.0777774
R1717 dvdd.n14 dvdd.n7 0.070241
R1718 dvdd.n25 dvdd.n24 0.0685285
R1719 dvdd.n267 dvdd 0.063
R1720 dvdd.n263 dvdd 0.0603958
R1721 dvdd dvdd.n262 0.0603958
R1722 dvdd.n247 dvdd 0.0603958
R1723 dvdd.n118 dvdd 0.0603958
R1724 dvdd.n157 dvdd 0.0603958
R1725 dvdd.n158 dvdd 0.0603958
R1726 dvdd.n195 dvdd 0.0603958
R1727 dvdd.n196 dvdd 0.0603958
R1728 dvdd.n233 dvdd 0.0603958
R1729 dvdd.n234 dvdd 0.0603958
R1730 dvdd.n268 dvdd 0.0603958
R1731 dvdd dvdd.n13 0.0595278
R1732 dvdd.n21 dvdd.n16 0.0535523
R1733 dvdd.n12 dvdd 0.0508472
R1734 dvdd.n290 dvdd.n289 0.0456945
R1735 dvdd.n39 dvdd.n38 0.0456858
R1736 dvdd.n20 dvdd 0.0405
R1737 dvdd dvdd.n296 0.0385435
R1738 dvdd dvdd.n246 0.0382604
R1739 dvdd.n39 dvdd.n0 0.0379437
R1740 dvdd.n21 dvdd 0.0339302
R1741 dvdd.n13 dvdd.n12 0.0334861
R1742 dvdd.n274 dvdd 0.03175
R1743 dvdd dvdd.n157 0.03175
R1744 dvdd dvdd.n195 0.03175
R1745 dvdd dvdd.n233 0.03175
R1746 dvdd.n268 dvdd 0.03175
R1747 dvdd.n24 dvdd.n16 0.0300191
R1748 dvdd.n247 dvdd 0.0239375
R1749 dvdd.n49 dvdd.n0 0.0233041
R1750 dvdd.n262 dvdd 0.0226354
R1751 dvdd dvdd.n156 0.0226354
R1752 dvdd dvdd.n194 0.0226354
R1753 dvdd dvdd.n232 0.0226354
R1754 dvdd dvdd.n241 0.0226354
R1755 dvdd.n298 dvdd.n297 0.0219531
R1756 dvdd.n15 dvdd 0.0210592
R1757 dvdd.n20 dvdd.n19 0.0205
R1758 dvdd.n51 dvdd 0.0188824
R1759 dvdd.n48 dvdd.n1 0.0182365
R1760 dvdd.n25 dvdd 0.0179419
R1761 dvdd.n49 dvdd.n48 0.0151396
R1762 dvdd.n289 dvdd.n280 0.0150881
R1763 dvdd dvdd.n20 0.0121279
R1764 dvdd.n298 dvdd.n280 0.00936728
R1765 dvdd.n267 dvdd.n242 0.0083125
R1766 dvdd.n276 dvdd.t178 0.0083125
R1767 dvdd.n277 dvdd.t177 0.0083125
R1768 dvdd.n278 dvdd.t176 0.0083125
R1769 dvdd.n50 dvdd.t175 0.0083125
R1770 dvdd.n297 dvdd 0.00765103
R1771 dvdd.n279 dvdd.n50 0.00754239
R1772 dvdd.n1 dvdd 0.00176689
R1773 dvdd.n298 dvdd 0.001125
R1774 a_20376_n2791.n1 a_20376_n2791.n0 926.024
R1775 a_20376_n2791.n1 a_20376_n2791.t2 82.0838
R1776 a_20376_n2791.n0 a_20376_n2791.t3 63.3338
R1777 a_20376_n2791.t0 a_20376_n2791.n1 63.3219
R1778 a_20376_n2791.n0 a_20376_n2791.t1 29.7268
R1779 a_19955_n2241.n1 a_19955_n2241.t7 530.01
R1780 a_19955_n2241.t1 a_19955_n2241.n5 421.021
R1781 a_19955_n2241.n0 a_19955_n2241.t2 337.142
R1782 a_19955_n2241.n3 a_19955_n2241.t0 280.223
R1783 a_19955_n2241.n4 a_19955_n2241.t3 263.173
R1784 a_19955_n2241.n4 a_19955_n2241.t5 227.826
R1785 a_19955_n2241.n0 a_19955_n2241.t4 199.762
R1786 a_19955_n2241.n2 a_19955_n2241.n1 170.81
R1787 a_19955_n2241.n2 a_19955_n2241.n0 167.321
R1788 a_19955_n2241.n5 a_19955_n2241.n4 152
R1789 a_19955_n2241.n1 a_19955_n2241.t6 141.923
R1790 a_19955_n2241.n3 a_19955_n2241.n2 10.8376
R1791 a_19955_n2241.n5 a_19955_n2241.n3 2.50485
R1792 a_20689_n2273.n3 a_20689_n2273.n2 647.119
R1793 a_20689_n2273.n1 a_20689_n2273.t4 350.253
R1794 a_20689_n2273.n2 a_20689_n2273.n0 260.339
R1795 a_20689_n2273.n2 a_20689_n2273.n1 246.119
R1796 a_20689_n2273.n1 a_20689_n2273.t5 189.588
R1797 a_20689_n2273.n3 a_20689_n2273.t0 89.1195
R1798 a_20689_n2273.n0 a_20689_n2273.t2 63.3338
R1799 a_20689_n2273.t1 a_20689_n2273.n3 41.0422
R1800 a_20689_n2273.n0 a_20689_n2273.t3 31.9797
R1801 a_21036_n1869.n3 a_21036_n1869.n2 636.953
R1802 a_21036_n1869.n1 a_21036_n1869.t5 366.856
R1803 a_21036_n1869.n2 a_21036_n1869.n0 300.2
R1804 a_21036_n1869.n2 a_21036_n1869.n1 225.036
R1805 a_21036_n1869.n1 a_21036_n1869.t4 174.056
R1806 a_21036_n1869.n0 a_21036_n1869.t2 70.0005
R1807 a_21036_n1869.t0 a_21036_n1869.n3 68.0124
R1808 a_21036_n1869.n3 a_21036_n1869.t3 63.3219
R1809 a_21036_n1869.n0 a_21036_n1869.t1 61.6672
R1810 a_10620_n8338.t0 a_10620_n8338.t1 83.9243
R1811 a_24220_n8172.t0 a_24220_n8172.t1 83.56
R1812 a_16620_n2791.n3 a_16620_n2791.n2 636.953
R1813 a_16620_n2791.n1 a_16620_n2791.t4 366.856
R1814 a_16620_n2791.n2 a_16620_n2791.n0 300.2
R1815 a_16620_n2791.n2 a_16620_n2791.n1 225.036
R1816 a_16620_n2791.n1 a_16620_n2791.t5 174.056
R1817 a_16620_n2791.n0 a_16620_n2791.t3 70.0005
R1818 a_16620_n2791.n3 a_16620_n2791.t2 68.0124
R1819 a_16620_n2791.t0 a_16620_n2791.n3 63.3219
R1820 a_16620_n2791.n0 a_16620_n2791.t1 61.6672
R1821 a_16974_n2791.t0 a_16974_n2791.t1 87.1434
R1822 a_16795_n2817.n4 a_16795_n2817.n0 746.659
R1823 a_16795_n2817.n5 a_16795_n2817.t3 389.183
R1824 a_16795_n2817.n1 a_16795_n2817.t7 256.988
R1825 a_16795_n2817.n6 a_16795_n2817.n5 251.167
R1826 a_16795_n2817.t0 a_16795_n2817.n6 223.571
R1827 a_16795_n2817.n3 a_16795_n2817.t5 212.081
R1828 a_16795_n2817.n4 a_16795_n2817.n3 181.942
R1829 a_16795_n2817.n5 a_16795_n2817.t8 174.891
R1830 a_16795_n2817.n1 a_16795_n2817.t4 163.803
R1831 a_16795_n2817.n2 a_16795_n2817.t6 139.78
R1832 a_16795_n2817.n2 a_16795_n2817.n1 129.264
R1833 a_16795_n2817.n0 a_16795_n2817.t1 63.3219
R1834 a_16795_n2817.n0 a_16795_n2817.t2 63.3219
R1835 a_16795_n2817.n6 a_16795_n2817.n4 24.6993
R1836 a_16795_n2817.n3 a_16795_n2817.n2 22.6399
R1837 ena_ip.t1 ena_ip.n1 744.115
R1838 ena_ip ena_ip.t1 732.75
R1839 ena_ip.n16 ena_ip.t7 408.63
R1840 ena_ip.n12 ena_ip.t13 408.63
R1841 ena_ip.n8 ena_ip.t4 408.63
R1842 ena_ip.n13 ena_ip.t6 347.577
R1843 ena_ip.n9 ena_ip.t8 347.577
R1844 ena_ip.n5 ena_ip.t16 347.577
R1845 ena_ip.n3 ena_ip.t14 332.752
R1846 ena_ip.t14 ena_ip.n2 332.752
R1847 ena_ip.n3 ena_ip.t17 332.411
R1848 ena_ip.t17 ena_ip.n2 332.411
R1849 ena_ip.n17 ena_ip.t19 239.505
R1850 ena_ip ena_ip.t0 216.155
R1851 ena_ip.n13 ena_ip.t9 193.337
R1852 ena_ip.n9 ena_ip.t10 193.337
R1853 ena_ip.n5 ena_ip.t18 193.337
R1854 ena_ip.n17 ena_ip.t11 167.204
R1855 ena_ip ena_ip.n16 165.089
R1856 ena_ip ena_ip.n12 165.089
R1857 ena_ip ena_ip.n8 165.089
R1858 ena_ip ena_ip.n17 157.12
R1859 ena_ip.n14 ena_ip.n13 152
R1860 ena_ip.n10 ena_ip.n9 152
R1861 ena_ip.n6 ena_ip.n5 152
R1862 ena_ip.n16 ena_ip.t3 132.282
R1863 ena_ip.n12 ena_ip.t5 132.282
R1864 ena_ip.n8 ena_ip.t15 132.282
R1865 ena_ip.n0 ena_ip.t2 59.9857
R1866 ena_ip ena_ip.t12 59.0936
R1867 ena_ip.n1 ena_ip 57.4755
R1868 ena_ip ena_ip.n18 13.8078
R1869 ena_ip.n18 ena_ip 9.82907
R1870 ena_ip ena_ip.n7 9.3005
R1871 ena_ip ena_ip.n11 9.3005
R1872 ena_ip ena_ip.n15 9.3005
R1873 ena_ip ena_ip.n19 8.84514
R1874 ena_ip.n18 ena_ip 5.71479
R1875 ena_ip.n4 ena_ip.n2 5.53161
R1876 ena_ip.n14 ena_ip 4.67077
R1877 ena_ip.n10 ena_ip 4.67077
R1878 ena_ip.n6 ena_ip 4.67077
R1879 ena_ip.n4 ena_ip.n3 4.67076
R1880 ena_ip.n19 ena_ip 4.17561
R1881 ena_ip.n1 ena_ip 3.62625
R1882 ena_ip.n0 ena_ip.n4 3.51723
R1883 ena_ip.n15 ena_ip 2.94104
R1884 ena_ip.n11 ena_ip 2.94104
R1885 ena_ip.n7 ena_ip 2.94104
R1886 ena_ip.n15 ena_ip.n14 2.76807
R1887 ena_ip.n11 ena_ip.n10 2.76807
R1888 ena_ip.n7 ena_ip.n6 2.76807
R1889 ena_ip ena_ip.n0 1.97628
R1890 ena_ip.n19 ena_ip 1.86127
R1891 x3.in_b.n1 x3.in_b.n0 3.2348
R1892 x3.in_b.n1 x3.in_b.t3 166.376
R1893 x3.in_b.n1 x3.in_b.t2 166.207
R1894 x3.in_b.n0 x3.in_b.t0 228.429
R1895 x3.in_b.n0 x3.in_b.t1 83.9309
R1896 a_21211_n1943.n6 a_21211_n1943.n5 746.659
R1897 a_21211_n1943.n0 a_21211_n1943.t6 389.183
R1898 a_21211_n1943.n2 a_21211_n1943.t4 256.988
R1899 a_21211_n1943.n1 a_21211_n1943.n0 251.167
R1900 a_21211_n1943.n1 a_21211_n1943.t1 223.571
R1901 a_21211_n1943.n4 a_21211_n1943.t7 212.081
R1902 a_21211_n1943.n5 a_21211_n1943.n4 181.942
R1903 a_21211_n1943.n0 a_21211_n1943.t8 174.891
R1904 a_21211_n1943.n2 a_21211_n1943.t5 163.803
R1905 a_21211_n1943.n3 a_21211_n1943.t3 139.78
R1906 a_21211_n1943.n3 a_21211_n1943.n2 129.264
R1907 a_21211_n1943.t0 a_21211_n1943.n6 63.3219
R1908 a_21211_n1943.n6 a_21211_n1943.t2 63.3219
R1909 a_21211_n1943.n5 a_21211_n1943.n1 24.6993
R1910 a_21211_n1943.n4 a_21211_n1943.n3 22.6399
R1911 a_17913_n2791.t0 a_17913_n2791.n3 370.026
R1912 a_17913_n2791.n0 a_17913_n2791.t2 351.356
R1913 a_17913_n2791.n1 a_17913_n2791.t5 334.717
R1914 a_17913_n2791.n3 a_17913_n2791.t1 325.971
R1915 a_17913_n2791.n1 a_17913_n2791.t4 309.935
R1916 a_17913_n2791.n0 a_17913_n2791.t3 305.683
R1917 a_17913_n2791.n2 a_17913_n2791.n0 16.879
R1918 a_17913_n2791.n3 a_17913_n2791.n2 10.8867
R1919 a_17913_n2791.n2 a_17913_n2791.n1 9.3005
R1920 a_18481_n2549.n3 a_18481_n2549.n2 647.119
R1921 a_18481_n2549.n1 a_18481_n2549.t4 350.253
R1922 a_18481_n2549.n2 a_18481_n2549.n0 260.339
R1923 a_18481_n2549.n2 a_18481_n2549.n1 246.119
R1924 a_18481_n2549.n1 a_18481_n2549.t5 189.588
R1925 a_18481_n2549.n3 a_18481_n2549.t1 89.1195
R1926 a_18481_n2549.n0 a_18481_n2549.t0 63.3338
R1927 a_18481_n2549.t2 a_18481_n2549.n3 41.0422
R1928 a_18481_n2549.n0 a_18481_n2549.t3 31.9797
R1929 a_18828_n2791.n3 a_18828_n2791.n2 636.953
R1930 a_18828_n2791.n1 a_18828_n2791.t4 366.856
R1931 a_18828_n2791.n2 a_18828_n2791.n0 300.2
R1932 a_18828_n2791.n2 a_18828_n2791.n1 225.036
R1933 a_18828_n2791.n1 a_18828_n2791.t5 174.056
R1934 a_18828_n2791.n0 a_18828_n2791.t0 70.0005
R1935 a_18828_n2791.n3 a_18828_n2791.t2 68.0124
R1936 a_18828_n2791.t1 a_18828_n2791.n3 63.3219
R1937 a_18828_n2791.n0 a_18828_n2791.t3 61.6672
R1938 a_2130_n19848.t0 a_2130_n19848.t1 82.0028
R1939 a_24530_n20014.t0 a_24530_n20014.t1 81.9478
R1940 icnode.t1 icnode 84.0284
R1941 icnode icnode.n3 0.00744444
R1942 icnode icnode.n3 0.00851282
R1943 icnode.n3 icnode.n2 0.0822308
R1944 icnode icnode.n2 0.0585357
R1945 icnode.n2 icnode.t0 1.17945
R1946 icnode icnode.n2 0.224859
R1947 icnode.n2 icnode.n1 1.59826
R1948 icnode icnode.n1 1.42175
R1949 icnode.n1 icnode.n0 0.463625
R1950 icnode.n0 icnode.t2 6.12107
R1951 icnode.n0 icnode.t3 5.08419
R1952 a_11526_n12394.t0 a_11526_n12394.t1 78.7148
R1953 vbreg.n7 vbreg.t0 245.107
R1954 vbreg.n55 vbreg.n50 202.542
R1955 vbreg.n44 vbreg.n2 201.036
R1956 vbreg.n36 vbreg.n15 200.282
R1957 vbreg.n7 vbreg.t3 22.4293
R1958 vbreg.t2 vbreg.n6 21.8369
R1959 vbreg.n46 vbreg.n27 179.953
R1960 vbreg.n39 vbreg.n2 179.201
R1961 vbreg.n50 vbreg.n27 178.447
R1962 vbreg.n39 vbreg.n15 176.941
R1963 vbreg.n46 vbreg.n10 1.98197
R1964 vbreg.n39 vbreg.n20 116.609
R1965 vbreg.n39 vbreg.n16 116.609
R1966 vbreg.n34 vbreg.n2 116.609
R1967 vbreg.n18 vbreg.n2 116.609
R1968 vbreg.n48 vbreg.n27 116.609
R1969 vbreg.n61 vbreg.n27 116.609
R1970 vbreg.n58 vbreg.n50 116.609
R1971 vbreg.n50 vbreg.n28 116.609
R1972 vbreg.n19 vbreg.n15 116.609
R1973 vbreg.n17 vbreg.n15 116.609
R1974 vbreg.n46 vbreg.n29 115.162
R1975 vbreg.t13 vbreg.n24 86.3125
R1976 vbreg.n37 vbreg.t10 86.3125
R1977 vbreg.n19 vbreg.t14 86.3125
R1978 vbreg.t12 vbreg.n17 86.3125
R1979 vbreg.t23 vbreg.n53 86.3125
R1980 vbreg.n56 vbreg.t25 86.3125
R1981 vbreg.t17 vbreg.n42 86.3125
R1982 vbreg.n31 vbreg.t18 86.3125
R1983 vbreg.n16 vbreg.t9 86.3125
R1984 vbreg.n20 vbreg.t11 86.3125
R1985 vbreg.n41 vbreg.t15 86.3125
R1986 vbreg.n33 vbreg.t16 86.3125
R1987 vbreg.n62 vbreg.t6 86.3125
R1988 vbreg.n47 vbreg.t20 86.3125
R1989 vbreg.n60 vbreg.t19 86.3125
R1990 vbreg.n59 vbreg.t22 86.3125
R1991 vbreg.n52 vbreg.t21 86.3125
R1992 vbreg.n57 vbreg.t24 86.3125
R1993 vbreg.n17 vbreg.n37 72.5338
R1994 vbreg.n42 vbreg.n41 72.5338
R1995 vbreg.n53 vbreg.n52 72.5338
R1996 vbreg.n19 vbreg.n24 72.5338
R1997 vbreg.n33 vbreg.n31 72.5338
R1998 vbreg.n57 vbreg.n56 72.5338
R1999 vbreg.n16 vbreg.n18 71.7809
R2000 vbreg.n62 vbreg.n61 71.7809
R2001 vbreg.n20 vbreg.n34 71.7809
R2002 vbreg.n31 vbreg.n29 71.7809
R2003 vbreg.n48 vbreg.n47 71.7809
R2004 vbreg.n17 vbreg.n14 2.62088
R2005 vbreg.n13 vbreg.n19 2.62088
R2006 vbreg.n60 vbreg.n28 71.2789
R2007 vbreg.n59 vbreg.n58 71.2789
R2008 vbreg.n4 vbreg.t7 60.1061
R2009 vbreg.n42 vbreg.n9 2.20744
R2010 vbreg.n35 vbreg.t13 55.9125
R2011 vbreg.n35 vbreg.t10 55.9125
R2012 vbreg.t14 vbreg.n38 55.9125
R2013 vbreg.n38 vbreg.t12 55.9125
R2014 vbreg.n54 vbreg.t23 55.9125
R2015 vbreg.n54 vbreg.t25 55.9125
R2016 vbreg.n43 vbreg.t17 55.9125
R2017 vbreg.n43 vbreg.t18 55.9125
R2018 vbreg.t9 vbreg.n40 55.9125
R2019 vbreg.n40 vbreg.t11 55.9125
R2020 vbreg.n30 vbreg.t15 55.9125
R2021 vbreg.t16 vbreg.n30 55.9125
R2022 vbreg.n45 vbreg.t6 55.9125
R2023 vbreg.n45 vbreg.t20 55.9125
R2024 vbreg.n49 vbreg.t19 55.9125
R2025 vbreg.t22 vbreg.n49 55.9125
R2026 vbreg.t21 vbreg.n51 55.9125
R2027 vbreg.n51 vbreg.t24 55.9125
R2028 vbreg.n36 vbreg.n35 30.4005
R2029 vbreg.n55 vbreg.n54 30.4005
R2030 vbreg.n40 vbreg.n39 30.4005
R2031 vbreg.n30 vbreg.n2 30.4005
R2032 vbreg.n44 vbreg.n43 30.4005
R2033 vbreg.n46 vbreg.n45 30.4005
R2034 vbreg.n49 vbreg.n27 30.4005
R2035 vbreg.n51 vbreg.n50 30.4005
R2036 vbreg.n38 vbreg.n15 30.4005
R2037 vbreg.n11 vbreg.t8 20.967
R2038 vbreg.n11 vbreg.t5 21.221
R2039 vbreg.n26 vbreg.t1 21.2773
R2040 vbreg.n10 vbreg.n4 0.049973
R2041 vbreg.n4 vbreg.n9 0.0436067
R2042 vbreg.n44 vbreg.n10 2.89594
R2043 vbreg.n25 vbreg.n24 2.80002
R2044 vbreg.n56 vbreg.n23 2.74579
R2045 vbreg.n23 vbreg.n55 2.3255
R2046 vbreg.n21 vbreg.n27 2.3255
R2047 vbreg.n22 vbreg.n50 2.3255
R2048 vbreg.n60 vbreg.n8 2.3255
R2049 vbreg.n53 vbreg.n23 2.3255
R2050 vbreg.n52 vbreg.n8 2.3255
R2051 vbreg.n12 vbreg.n59 2.3255
R2052 vbreg.n57 vbreg.n12 2.3255
R2053 vbreg.n25 vbreg.n36 2.3255
R2054 vbreg.n37 vbreg.n25 2.3255
R2055 vbreg.n39 vbreg.n0 2.3255
R2056 vbreg.n41 vbreg.n3 2.3255
R2057 vbreg.n3 vbreg.n2 2.3255
R2058 vbreg.n33 vbreg.n32 2.3255
R2059 vbreg.n31 vbreg.n5 2.3255
R2060 vbreg.n47 vbreg.n5 2.3255
R2061 vbreg.n9 vbreg.n62 2.10407
R2062 vbreg.n5 vbreg.n4 1.77403
R2063 vbreg.n4 vbreg.n7 1.69472
R2064 vbreg.n52 vbreg.n28 1.2554
R2065 vbreg.n58 vbreg.n57 1.2554
R2066 vbreg.t4 vbreg.n26 21.2177
R2067 vbreg.n20 vbreg.n13 2.62088
R2068 vbreg.n1 vbreg.n13 0.429184
R2069 vbreg.n14 vbreg.n16 2.62088
R2070 vbreg.n32 vbreg.n3 1.38145
R2071 vbreg.n4 vbreg.n8 1.3464
R2072 vbreg.n21 vbreg.n12 1.22472
R2073 vbreg.n32 vbreg.n5 1.22324
R2074 vbreg.n1 vbreg.n0 0.325142
R2075 vbreg.n8 vbreg.n22 1.17859
R2076 vbreg.n3 vbreg.n0 1.02185
R2077 vbreg.n8 vbreg.n23 0.922356
R2078 vbreg.n25 vbreg.n0 0.915412
R2079 vbreg.n7 vbreg.n6 0.00467336
R2080 vbreg.n26 vbreg.n7 0.845047
R2081 vbreg.n11 vbreg.n6 0.800043
R2082 vbreg.n14 vbreg.n0 0.795018
R2083 vbreg.n41 vbreg.n18 0.753441
R2084 vbreg.n61 vbreg.n60 0.753441
R2085 vbreg.n34 vbreg.n33 0.753441
R2086 vbreg.n47 vbreg.n29 0.753441
R2087 vbreg.n59 vbreg.n48 0.753441
R2088 vbreg.n8 vbreg.n21 0.690976
R2089 vbreg.n22 vbreg.n12 0.690976
R2090 vbreg.n1 vbreg.n15 2.50917
R2091 a_15000_n2791.n2 a_15000_n2791.n1 682.193
R2092 a_15000_n2791.n0 a_15000_n2791.t4 279.142
R2093 a_15000_n2791.n1 a_15000_n2791.t1 250.526
R2094 a_15000_n2791.n0 a_15000_n2791.t3 145.958
R2095 a_15000_n2791.n1 a_15000_n2791.n0 118.642
R2096 a_15000_n2791.n2 a_15000_n2791.t2 70.3576
R2097 a_15000_n2791.t0 a_15000_n2791.n2 65.6672
R2098 x7.x2.x2.CLK x7.x2.x2.CLK.t0 721.571
R2099 x7.x2.x2.CLK.n2 x7.x2.x2.CLK.t0 707.66
R2100 x7.x2.x2.CLK.n0 x7.x2.x2.CLK.t2 294.557
R2101 x7.x2.x2.CLK.n1 x7.x2.x2.CLK.t1 271.777
R2102 x7.x2.x2.CLK.n0 x7.x2.x2.CLK.t3 211.01
R2103 x7.x2.x2.CLK x7.x2.x2.CLK.n0 152
R2104 x7.x2.x2.CLK.n2 x7.x2.x2.CLK.n1 38.2982
R2105 x7.x2.x2.CLK.n1 x7.x2.x2.CLK 32.5125
R2106 x7.x2.x2.CLK x7.x2.x2.CLK.n2 3.76521
R2107 x7.x1.x4.CLK.n3 x7.x1.x4.CLK.t1 372.361
R2108 x7.x1.x4.CLK.n2 x7.x1.x4.CLK.t2 333.651
R2109 x7.x1.x4.CLK.n2 x7.x1.x4.CLK.t5 297.233
R2110 x7.x1.x4.CLK.n0 x7.x1.x4.CLK.t3 294.557
R2111 x7.x1.x4.CLK.n4 x7.x1.x4.CLK.t0 231.921
R2112 x7.x1.x4.CLK.n0 x7.x1.x4.CLK.t4 211.01
R2113 x7.x1.x4.CLK x7.x1.x4.CLK.n2 195.701
R2114 x7.x1.x4.CLK.n1 x7.x1.x4.CLK.n0 152
R2115 x7.x1.x4.CLK.n4 x7.x1.x4.CLK.n1 41.5091
R2116 x7.x1.x4.CLK.n3 x7.x1.x4.CLK 25.2781
R2117 x7.x1.x4.CLK.n4 x7.x1.x4.CLK.n3 18.1966
R2118 x7.x1.x4.CLK.n1 x7.x1.x4.CLK 4.20621
R2119 x7.x1.x4.CLK x7.x1.x4.CLK.n4 2.5605
R2120 a_18168_n1881.n1 a_18168_n1881.n0 926.024
R2121 a_18168_n1881.t0 a_18168_n1881.n1 82.0838
R2122 a_18168_n1881.n0 a_18168_n1881.t1 63.3338
R2123 a_18168_n1881.n1 a_18168_n1881.t2 63.3219
R2124 a_18168_n1881.n0 a_18168_n1881.t3 29.7268
R2125 vbp vbp.t11 150.532
R2126 vbp.n1 vbp.n0 24.4313
R2127 vbp.n8 vbp 145.601
R2128 vbp vbp.t2 111.784
R2129 vbp vbp.t12 64.09
R2130 vbp.n3 vbp.t6 21.3499
R2131 vbp.n2 vbp.t13 21.3436
R2132 vbp.n3 vbp.n0 8.69141
R2133 vbp.n5 vbp 70.6788
R2134 vbp vbp.t1 68.2084
R2135 vbp vbp.t3 62.2125
R2136 vbp.t10 vbp.n0 62.2125
R2137 vbp vbp.t14 62.2125
R2138 vbp vbp.t4 62.2125
R2139 vbp vbp.t7 62.2125
R2140 vbp.t9 vbp.n6 62.2125
R2141 vbp.n0 vbp.n2 8.19623
R2142 vbp.n6 vbp 54.6138
R2143 vbp.n6 vbp 54.6138
R2144 vbp.n5 vbp 44.5222
R2145 vbp vbp.t0 40.0025
R2146 vbp.n3 vbp.t16 20.9636
R2147 vbp.t3 vbp.n10 31.8125
R2148 vbp.n10 vbp.t10 31.8125
R2149 vbp.t14 vbp.n9 31.8125
R2150 vbp.n9 vbp.t4 31.8125
R2151 vbp.n7 vbp.t7 31.8125
R2152 vbp.t12 vbp.n7 31.8125
R2153 vbp.n8 vbp.t17 31.8125
R2154 vbp.t11 vbp.n8 31.8125
R2155 vbp.n11 vbp.t1 31.8125
R2156 vbp.n11 vbp.t9 31.8125
R2157 vbp.t8 vbp.n2 20.9685
R2158 vbp.n1 vbp.t15 31.8136
R2159 vbp.n7 vbp 30.4005
R2160 vbp.n9 vbp 30.4005
R2161 vbp.n5 vbp.n11 30.4005
R2162 vbp.n10 vbp 30.4005
R2163 vbp.n4 vbp.n6 1.72982
R2164 vbp.n4 vbp.n5 5.41061
R2165 vbp.t17 vbp 65.2042
R2166 vbp.n4 vbp 17.0614
R2167 vbp.n0 vbp 11.5581
R2168 vbp.n1 vbp.t5 16.8504
R2169 dvdd_ip.n8 dvdd_ip.n6 12175.6
R2170 dvdd_ip.n7 dvdd_ip.n6 12175.6
R2171 dvdd_ip.n70 dvdd_ip.n8 2.31015
R2172 dvdd_ip.n8 dvdd_ip.n10 12175.6
R2173 dvdd_ip.n7 dvdd_ip.n10 12175.6
R2174 dvdd_ip.n71 dvdd_ip.n7 2.31015
R2175 dvdd_ip.n103 dvdd_ip.n33 10440
R2176 dvdd_ip.n105 dvdd_ip.n33 10440
R2177 dvdd_ip.n105 dvdd_ip.n34 10440
R2178 dvdd_ip.n103 dvdd_ip.n34 10440
R2179 dvdd_ip.n64 dvdd_ip.n9 4516.33
R2180 dvdd_ip.n71 dvdd_ip.n9 4243.24
R2181 dvdd_ip.n62 dvdd_ip.n61 4030.59
R2182 dvdd_ip.n59 dvdd_ip.n57 4030.59
R2183 dvdd_ip.n91 dvdd_ip.n48 4030.59
R2184 dvdd_ip.n94 dvdd_ip.n47 4030.59
R2185 dvdd_ip.n53 dvdd_ip.n20 3741.35
R2186 dvdd_ip.n70 dvdd_ip.n53 3618.82
R2187 dvdd_ip.n96 dvdd_ip.n43 3190.03
R2188 dvdd_ip.n98 dvdd_ip.n43 3190.03
R2189 dvdd_ip.n98 dvdd_ip.n44 3190.03
R2190 dvdd_ip.n96 dvdd_ip.n44 3190.03
R2191 dvdd_ip.n73 dvdd_ip.n24 2795.29
R2192 dvdd_ip.n76 dvdd_ip.n52 2795.29
R2193 dvdd_ip.n84 dvdd_ip.n50 2417.65
R2194 dvdd_ip.n84 dvdd_ip.n51 2417.65
R2195 dvdd_ip.n82 dvdd_ip.n51 2417.65
R2196 dvdd_ip.n82 dvdd_ip.n50 2417.65
R2197 dvdd_ip.n93 dvdd_ip.n48 1199.77
R2198 dvdd_ip.n92 dvdd_ip.n47 1199.77
R2199 dvdd_ip.n75 dvdd_ip.n24 703.912
R2200 dvdd_ip.n74 dvdd_ip.n52 703.912
R2201 dvdd_ip.n64 dvdd_ip.n63 654.165
R2202 dvdd_ip.n49 dvdd_ip.t13 642.13
R2203 dvdd_ip.n26 dvdd_ip.t21 642.383
R2204 dvdd_ip.n46 dvdd_ip.t7 642.13
R2205 dvdd_ip.t56 dvdd_ip.n78 594.953
R2206 dvdd_ip.t56 dvdd_ip.n79 594.301
R2207 dvdd_ip.n58 dvdd_ip.n55 429.93
R2208 dvdd_ip.n63 dvdd_ip.n55 429.93
R2209 dvdd_ip.t40 dvdd_ip.t24 397.805
R2210 dvdd_ip.t34 dvdd_ip.t40 397.805
R2211 dvdd_ip.t36 dvdd_ip.t34 397.805
R2212 dvdd_ip.t27 dvdd_ip.t42 397.805
R2213 dvdd_ip.t38 dvdd_ip.t27 397.805
R2214 dvdd_ip.t29 dvdd_ip.t38 397.805
R2215 dvdd_ip.n58 dvdd_ip.n54 340.42
R2216 dvdd_ip.t2 dvdd_ip.n82 327.8
R2217 dvdd_ip.n84 dvdd_ip.t4 327.8
R2218 dvdd_ip.t9 dvdd_ip.t22 312.123
R2219 dvdd_ip.t10 dvdd_ip.t23 312.123
R2220 dvdd_ip.t22 dvdd_ip.n96 259.716
R2221 dvdd_ip.n98 dvdd_ip.t10 259.716
R2222 dvdd_ip.t24 dvdd_ip.n103 250.107
R2223 dvdd_ip.n105 dvdd_ip.t29 250.107
R2224 dvdd_ip.n95 dvdd_ip.n19 221.308
R2225 dvdd_ip.n104 dvdd_ip.t36 198.903
R2226 dvdd_ip.t42 dvdd_ip.n104 198.903
R2227 dvdd_ip.n83 dvdd_ip.t2 159.988
R2228 dvdd_ip.t4 dvdd_ip.n83 159.988
R2229 dvdd_ip.n97 dvdd_ip.t9 156.062
R2230 dvdd_ip.t23 dvdd_ip.n97 156.062
R2231 dvdd_ip.n29 dvdd_ip.n32 146.071
R2232 dvdd_ip.n102 dvdd_ip.n99 138.667
R2233 dvdd_ip.n100 dvdd_ip.n32 135.279
R2234 dvdd_ip.n1 dvdd_ip.t41 113.606
R2235 dvdd_ip.n0 dvdd_ip.t47 113.606
R2236 dvdd_ip.n15 dvdd_ip.t28 113.594
R2237 dvdd_ip.n16 dvdd_ip.t48 113.594
R2238 dvdd_ip.n39 dvdd_ip.t37 113.562
R2239 dvdd_ip.n39 dvdd_ip.t51 113.562
R2240 dvdd_ip.n2 dvdd_ip.t45 113.562
R2241 dvdd_ip.n2 dvdd_ip.t35 113.562
R2242 dvdd_ip.n15 dvdd_ip.t52 113.531
R2243 dvdd_ip.n31 dvdd_ip.t31 111.784
R2244 dvdd_ip.n36 dvdd_ip.t26 111.784
R2245 dvdd_ip.n35 dvdd_ip.t25 111.784
R2246 dvdd_ip.n38 dvdd_ip.t33 111.784
R2247 dvdd_ip.n37 dvdd_ip.t32 111.784
R2248 dvdd_ip.n41 dvdd_ip.t44 111.784
R2249 dvdd_ip.n40 dvdd_ip.t43 111.784
R2250 dvdd_ip.n62 dvdd_ip.n56 106.282
R2251 dvdd_ip.n60 dvdd_ip.n59 106.282
R2252 dvdd_ip.n30 dvdd_ip.n29 102.18
R2253 dvdd_ip.n45 dvdd_ip.n42 89.4643
R2254 dvdd_ip.n17 dvdd_ip.n102 64.1367
R2255 dvdd_ip.n72 dvdd_ip.t1 60.3236
R2256 dvdd_ip.n79 dvdd_ip.t3 57.1305
R2257 dvdd_ip.n79 dvdd_ip.t12 57.1305
R2258 dvdd_ip.n78 dvdd_ip.t17 57.1305
R2259 dvdd_ip.n78 dvdd_ip.t5 57.1305
R2260 dvdd_ip.n86 dvdd_ip.n22 55.1223
R2261 dvdd_ip.n14 dvdd_ip.n69 54.7105
R2262 dvdd_ip.n14 dvdd_ip.n66 54.7105
R2263 dvdd_ip.n14 dvdd_ip.n68 54.7085
R2264 dvdd_ip.n14 dvdd_ip.n67 54.7085
R2265 dvdd_ip.n14 dvdd_ip.n65 54.7085
R2266 dvdd_ip.n80 dvdd_ip.n49 53.6981
R2267 dvdd_ip.n3 dvdd_ip.n26 7.75105
R2268 dvdd_ip.n87 dvdd_ip.n47 46.2505
R2269 dvdd_ip.n88 dvdd_ip.n48 46.2505
R2270 dvdd_ip.n57 dvdd_ip.n54 46.2505
R2271 dvdd_ip.n61 dvdd_ip.n55 46.2505
R2272 dvdd_ip.n57 dvdd_ip.n56 44.5206
R2273 dvdd_ip.n61 dvdd_ip.n60 44.5206
R2274 dvdd_ip.n89 dvdd_ip.n88 37.2058
R2275 dvdd_ip.n52 dvdd_ip.n13 37.0005
R2276 dvdd_ip.n20 dvdd_ip.n24 37.0005
R2277 dvdd_ip.n86 dvdd_ip.n85 33.5615
R2278 dvdd_ip.n5 dvdd_ip.n21 1.04644
R2279 dvdd_ip.n89 dvdd_ip.n45 31.3351
R2280 dvdd_ip.n82 dvdd_ip.n13 26.4291
R2281 dvdd_ip.n85 dvdd_ip.n84 26.4291
R2282 dvdd_ip.n94 dvdd_ip.n5 12.8793
R2283 dvdd_ip.n3 dvdd_ip.n64 23.3225
R2284 dvdd_ip.n90 dvdd_ip.n89 22.576
R2285 dvdd_ip.n50 dvdd_ip.n22 20.5561
R2286 dvdd_ip.n83 dvdd_ip.n50 20.5561
R2287 dvdd_ip.n81 dvdd_ip.n51 20.5561
R2288 dvdd_ip.n83 dvdd_ip.n51 20.5561
R2289 dvdd_ip.n81 dvdd_ip.n80 19.0763
R2290 dvdd_ip.n99 dvdd_ip.n19 18.9635
R2291 dvdd_ip.n85 dvdd_ip.n49 17.7956
R2292 dvdd_ip.n77 dvdd_ip.n20 17.833
R2293 dvdd_ip.n23 dvdd_ip.n77 17.5685
R2294 dvdd_ip.n36 dvdd_ip.n35 14.6565
R2295 dvdd_ip.n38 dvdd_ip.n37 14.6565
R2296 dvdd_ip.t30 dvdd_ip.n31 14.6565
R2297 dvdd_ip.t50 dvdd_ip.t49 14.6565
R2298 dvdd_ip.n5 dvdd_ip.n11 2.19457
R2299 dvdd_ip.n41 dvdd_ip.n40 14.299
R2300 dvdd_ip.n72 dvdd_ip.t56 0.604318
R2301 dvdd_ip.n23 dvdd_ip.n22 13.4443
R2302 dvdd_ip.n77 dvdd_ip.n76 13.2148
R2303 dvdd_ip.n73 dvdd_ip.n72 13.2148
R2304 dvdd_ip.n96 dvdd_ip.n11 12.3338
R2305 dvdd_ip.n99 dvdd_ip.n98 12.3338
R2306 dvdd_ip.n103 dvdd_ip.n19 11.563
R2307 dvdd_ip.n29 dvdd_ip.n105 11.563
R2308 dvdd_ip.n88 dvdd_ip.n11 11.1792
R2309 dvdd_ip.n71 dvdd_ip.n25 5.53168
R2310 dvdd_ip.n5 dvdd_ip.n45 11.0012
R2311 dvdd_ip.n101 dvdd_ip.n100 10.7927
R2312 dvdd_ip.n76 dvdd_ip.n75 9.84115
R2313 dvdd_ip.n74 dvdd_ip.n73 9.84115
R2314 dvdd_ip.n49 dvdd_ip.n5 9.4314
R2315 dvdd_ip.n5 dvdd_ip.n46 9.30175
R2316 dvdd_ip.n100 dvdd_ip.n4 9.3005
R2317 dvdd_ip.n17 dvdd_ip.n42 8.03454
R2318 dvdd_ip.n33 dvdd_ip.n18 15.3082
R2319 dvdd_ip.n91 dvdd_ip.n90 7.4005
R2320 dvdd_ip.n59 dvdd_ip.n58 7.4005
R2321 dvdd_ip.n63 dvdd_ip.n62 7.4005
R2322 dvdd_ip.n69 dvdd_ip.t15 7.14175
R2323 dvdd_ip.n69 dvdd_ip.t18 7.14175
R2324 dvdd_ip.n68 dvdd_ip.t14 7.14175
R2325 dvdd_ip.n68 dvdd_ip.t19 7.14175
R2326 dvdd_ip.n67 dvdd_ip.t8 7.14175
R2327 dvdd_ip.n67 dvdd_ip.t54 7.14175
R2328 dvdd_ip.n66 dvdd_ip.t53 7.14175
R2329 dvdd_ip.n66 dvdd_ip.t55 7.14175
R2330 dvdd_ip.n65 dvdd_ip.t11 7.14175
R2331 dvdd_ip.n65 dvdd_ip.t16 7.14175
R2332 dvdd_ip.n29 dvdd_ip.n28 1.82386
R2333 dvdd_ip.n95 dvdd_ip.n43 6.37981
R2334 dvdd_ip.n97 dvdd_ip.n43 6.37981
R2335 dvdd_ip.n44 dvdd_ip.n42 6.37981
R2336 dvdd_ip.n97 dvdd_ip.n44 6.37981
R2337 dvdd_ip.n87 dvdd_ip.n86 5.51614
R2338 dvdd_ip.n94 dvdd_ip.n93 5.18874
R2339 dvdd_ip.n92 dvdd_ip.n91 5.18874
R2340 dvdd_ip.t56 dvdd_ip.n81 3.8204
R2341 dvdd_ip.n75 dvdd_ip.t0 3.32862
R2342 dvdd_ip.t0 dvdd_ip.n74 3.32862
R2343 dvdd_ip.t56 dvdd_ip.n25 1.8903
R2344 dvdd_ip.n86 dvdd_ip.n5 3.14232
R2345 dvdd_ip.n35 dvdd_ip.n4 1.23063
R2346 dvdd_ip.n27 dvdd_ip.n101 8.0274
R2347 dvdd_ip.n29 dvdd_ip.t50 3.1045
R2348 dvdd_ip.n104 dvdd_ip.n33 2.76169
R2349 dvdd_ip.n34 dvdd_ip.n32 2.76169
R2350 dvdd_ip.n104 dvdd_ip.n34 2.76169
R2351 dvdd_ip.n21 dvdd_ip.n87 2.74244
R2352 dvdd_ip.n12 dvdd_ip.t56 0.384439
R2353 dvdd_ip.t6 dvdd_ip.n92 2.20373
R2354 dvdd_ip.n93 dvdd_ip.t6 2.20373
R2355 dvdd_ip.n70 dvdd_ip.n3 5.23222
R2356 dvdd_ip.n3 dvdd_ip.n40 2.01844
R2357 dvdd_ip.n102 dvdd_ip.n101 1.95955
R2358 dvdd_ip.n21 dvdd_ip.n80 9.20625
R2359 dvdd_ip.n37 dvdd_ip.n27 0.701705
R2360 dvdd_ip.n28 dvdd_ip.n3 1.0491
R2361 dvdd_ip.t50 dvdd_ip.n3 1.8605
R2362 dvdd_ip.n1 dvdd_ip.n36 1.8245
R2363 dvdd_ip.n0 dvdd_ip.n38 1.8245
R2364 dvdd_ip.t46 dvdd_ip.t30 1.7925
R2365 dvdd_ip.t49 dvdd_ip.t39 1.7925
R2366 dvdd_ip.n16 dvdd_ip.n41 1.74879
R2367 dvdd_ip.n4 dvdd_ip.n18 1.42286
R2368 dvdd_ip.n54 dvdd_ip.n26 1.22276
R2369 dvdd_ip.n18 dvdd_ip.n30 0.319081
R2370 dvdd_ip.n4 dvdd_ip.n39 1.343
R2371 dvdd_ip.n3 dvdd_ip.n30 1.2342
R2372 dvdd_ip.n5 dvdd_ip.n95 83.6014
R2373 dvdd_ip.n17 dvdd_ip.n5 1.7115
R2374 dvdd_ip.n4 dvdd_ip.n27 1.68015
R2375 dvdd_ip.n12 dvdd_ip.n13 0.973956
R2376 dvdd_ip.n3 dvdd_ip.n15 1.61215
R2377 dvdd_ip.n10 dvdd_ip.n9 1.53577
R2378 dvdd_ip.n53 dvdd_ip.n6 1.53577
R2379 dvdd_ip.n20 dvdd_ip.n25 1.39615
R2380 dvdd_ip.n19 dvdd_ip.n4 0.881757
R2381 dvdd_ip.n4 dvdd_ip.n17 1.26747
R2382 dvdd_ip.n28 dvdd_ip.n31 0.516501
R2383 dvdd_ip.n60 dvdd_ip.t20 1.22055
R2384 dvdd_ip.t20 dvdd_ip.n56 1.22055
R2385 dvdd_ip.n4 dvdd_ip.n3 1.12387
R2386 dvdd_ip.n90 dvdd_ip.n5 1.02666
R2387 dvdd_ip.n3 dvdd_ip.n14 0.974166
R2388 dvdd_ip.n3 dvdd_ip.n16 0.930808
R2389 dvdd_ip.n4 dvdd_ip.n1 0.9305
R2390 dvdd_ip.n4 dvdd_ip.n0 0.9305
R2391 dvdd_ip.n4 dvdd_ip.n2 0.9305
R2392 dvdd_ip.n3 dvdd_ip.t46 0.9305
R2393 dvdd_ip.t39 dvdd_ip.n3 0.9305
R2394 dvdd_ip.t56 dvdd_ip.n5 0.868735
R2395 dvdd_ip.n88 dvdd_ip.n46 0.83013
R2396 dvdd_ip.n12 dvdd_ip.n23 1.21666
R2397 tail.n4 tail.t4 113.562
R2398 tail.n4 tail.t9 113.562
R2399 tail.n3 tail.t7 113.562
R2400 tail.n3 tail.t2 113.562
R2401 tail.n5 tail.t11 113.562
R2402 tail.n5 tail.t6 113.562
R2403 tail.n7 tail.t3 113.562
R2404 tail.n7 tail.t8 113.562
R2405 tail.n6 tail.t5 113.562
R2406 tail.n6 tail.t10 113.562
R2407 tail.n2 tail.n1 53.5531
R2408 tail.n1 tail.t0 6.92425
R2409 tail.n1 tail.t1 6.92425
R2410 tail tail.n2 3.613
R2411 tail tail.n5 1.3055
R2412 tail.n0 tail.n4 1.1139
R2413 tail.n0 tail.n3 1.04033
R2414 tail.n6 tail 1.10604
R2415 tail.n2 tail 0.471179
R2416 tail.n7 tail 1.04408
R2417 tail tail.n0 1.02446
R2418 a_16273_n2549.n3 a_16273_n2549.n2 647.119
R2419 a_16273_n2549.n1 a_16273_n2549.t4 350.253
R2420 a_16273_n2549.n2 a_16273_n2549.n0 260.339
R2421 a_16273_n2549.n2 a_16273_n2549.n1 246.119
R2422 a_16273_n2549.n1 a_16273_n2549.t5 189.588
R2423 a_16273_n2549.n3 a_16273_n2549.t1 89.1195
R2424 a_16273_n2549.n0 a_16273_n2549.t3 63.3338
R2425 a_16273_n2549.t2 a_16273_n2549.n3 41.0422
R2426 a_16273_n2549.n0 a_16273_n2549.t0 31.9797
R2427 a_16151_n2791.t1 a_16151_n2791.t0 198.571
R2428 a_16317_n2791.t0 a_16317_n2791.t1 60.0005
R2429 x4.in_b.n5 x4.in_b.t14 408.63
R2430 x4.in_b.n7 x4.in_b.t25 408.63
R2431 x4.in_b.n9 x4.in_b.t11 408.63
R2432 x4.in_b.n0 x4.in_b.t19 187.875
R2433 x4.in_b.t16 x4.in_b.n1 188.125
R2434 x4.in_b.n0 x4.in_b.n1 0.276071
R2435 x4.in_b.t18 x4.in_b.n1 187.659
R2436 x4.in_b.t0 x4.in_b.n2 187.724
R2437 x4.in_b.n2 x4.in_b.t3 187.722
R2438 x4.in_b.n2 x4.in_b.n0 2.14521
R2439 x4.in_b.t23 x4.in_b.n3 187.724
R2440 x4.in_b.t17 x4.in_b.n0 187.716
R2441 x4.in_b.n13 x4.in_b.t13 347.577
R2442 x4.in_b.n12 x4.in_b.t15 347.577
R2443 x4.in_b.n11 x4.in_b.t2 347.577
R2444 x4.in_b.n4 x4.in_b.t12 332.752
R2445 x4.in_b.t12 x4.in_b 332.752
R2446 x4.in_b.n4 x4.in_b.t4 332.411
R2447 x4.in_b.t4 x4.in_b 332.411
R2448 x4.in_b.n14 x4.in_b.t24 236.552
R2449 x4.in_b.n13 x4.in_b.t8 193.337
R2450 x4.in_b.n12 x4.in_b.t9 193.337
R2451 x4.in_b.n11 x4.in_b.t22 193.337
R2452 x4.in_b x4.in_b.n5 165.089
R2453 x4.in_b x4.in_b.n7 165.089
R2454 x4.in_b x4.in_b.n9 165.089
R2455 x4.in_b.n14 x4.in_b.t10 164.251
R2456 x4.in_b x4.in_b.n14 154.47
R2457 x4.in_b x4.in_b.n13 152
R2458 x4.in_b x4.in_b.n12 152
R2459 x4.in_b x4.in_b.n11 152
R2460 x4.in_b.n5 x4.in_b.t1 132.282
R2461 x4.in_b.n7 x4.in_b.t5 132.282
R2462 x4.in_b.n9 x4.in_b.t20 132.282
R2463 x4.in_b.t6 x4.in_b.n0 187.133
R2464 x4.in_b.t7 x4.in_b.n0 187.724
R2465 x4.in_b.t21 x4.in_b.n3 187.722
R2466 x4.in_b.n6 x4.in_b 16.7098
R2467 x4.in_b x4.in_b.n6 14.0185
R2468 x4.in_b x4.in_b.n8 14.0185
R2469 x4.in_b x4.in_b.n10 14.0185
R2470 x4.in_b.n6 x4.in_b 11.4672
R2471 x4.in_b.n8 x4.in_b 11.4672
R2472 x4.in_b.n10 x4.in_b 11.4672
R2473 x4.in_b x4.in_b.n4 11.1417
R2474 x4.in_b x4.in_b.n0 10.4718
R2475 x4.in_b.n0 x4.in_b 10.4505
R2476 x4.in_b.n3 x4.in_b.n0 10.356
R2477 x4.in_b.n10 x4.in_b 9.3005
R2478 x4.in_b.n8 x4.in_b 9.3005
R2479 a_9120_n9346.n1 a_9120_n9346.t1 651.505
R2480 a_9120_n9346.n0 a_9120_n9346.t3 229.508
R2481 a_9120_n9346.t4 a_9120_n9346.n1 44.6806
R2482 a_9120_n9346.n1 a_9120_n9346.t0 5.54227
R2483 a_9120_n9346.n0 a_9120_n9346.t2 5.09877
R2484 a_9120_n9346.n1 a_9120_n9346.n0 0.631058
R2485 a_24220_n9832.t0 a_24220_n9832.t1 83.56
R2486 a_16974_n1881.t0 a_16974_n1881.t1 87.1434
R2487 a_16795_n1943.n6 a_16795_n1943.n5 746.659
R2488 a_16795_n1943.n0 a_16795_n1943.t8 389.183
R2489 a_16795_n1943.n2 a_16795_n1943.t4 256.988
R2490 a_16795_n1943.n1 a_16795_n1943.n0 251.167
R2491 a_16795_n1943.n1 a_16795_n1943.t1 223.571
R2492 a_16795_n1943.n4 a_16795_n1943.t5 212.081
R2493 a_16795_n1943.n5 a_16795_n1943.n4 181.942
R2494 a_16795_n1943.n0 a_16795_n1943.t7 174.891
R2495 a_16795_n1943.n2 a_16795_n1943.t6 163.803
R2496 a_16795_n1943.n3 a_16795_n1943.t3 139.78
R2497 a_16795_n1943.n3 a_16795_n1943.n2 129.264
R2498 a_16795_n1943.t0 a_16795_n1943.n6 63.3219
R2499 a_16795_n1943.n6 a_16795_n1943.t2 63.3219
R2500 a_16795_n1943.n5 a_16795_n1943.n1 24.6993
R2501 a_16795_n1943.n4 a_16795_n1943.n3 22.6399
R2502 a_21775_n2247.t0 a_21775_n2247.n1 386.31
R2503 a_21775_n2247.n1 a_21775_n2247.t1 249.956
R2504 a_21775_n2247.n0 a_21775_n2247.t2 239.04
R2505 a_21775_n2247.n1 a_21775_n2247.n0 175.661
R2506 a_21775_n2247.n0 a_21775_n2247.t3 166.739
R2507 x7.x3.B2.n8 x7.x3.B2.t0 373.866
R2508 x7.x3.B2.n6 x7.x3.B2.t5 333.651
R2509 x7.x3.B2.n6 x7.x3.B2.t6 297.233
R2510 x7.x3.B2 x7.x3.B2.t1 247.159
R2511 x7.x3.B2.n0 x7.x3.B2.t3 241.536
R2512 x7.x3.B2.n2 x7.x3.B2.t4 207.423
R2513 x7.x3.B2.n3 x7.x3.B2.t7 202.133
R2514 x7.x3.B2 x7.x3.B2.n6 195.701
R2515 x7.x3.B2.n0 x7.x3.B2.t2 169.237
R2516 x7.x3.B2.n5 x7.x3.B2.n2 159.758
R2517 x7.x3.B2.n1 x7.x3.B2.n0 155.84
R2518 x7.x3.B2.n4 x7.x3.B2.n3 152
R2519 x7.x3.B2.n3 x7.x3.B2.n2 36.8275
R2520 x7.x3.B2 x7.x3.B2.n8 16.6907
R2521 x7.x3.B2.n7 x7.x3.B2 15.8995
R2522 x7.x3.B2.n7 x7.x3.B2 15.6656
R2523 x7.x3.B2 x7.x3.B2.n5 13.8109
R2524 x7.x3.B2 x7.x3.B2.n1 12.822
R2525 x7.x3.B2.n5 x7.x3.B2.n4 5.4308
R2526 x7.x3.B2.n4 x7.x3.B2 3.68535
R2527 x7.x3.B2.n1 x7.x3.B2 3.2005
R2528 x7.x3.B2.n8 x7.x3.B2.n7 3.1005
R2529 a_20121_n2241.t0 a_20121_n2241.n3 370.026
R2530 a_20121_n2241.n0 a_20121_n2241.t2 351.356
R2531 a_20121_n2241.n1 a_20121_n2241.t4 334.717
R2532 a_20121_n2241.n3 a_20121_n2241.t1 325.971
R2533 a_20121_n2241.n1 a_20121_n2241.t5 309.935
R2534 a_20121_n2241.n0 a_20121_n2241.t3 305.683
R2535 a_20121_n2241.n2 a_20121_n2241.n0 16.879
R2536 a_20121_n2241.n3 a_20121_n2241.n2 10.8867
R2537 a_20121_n2241.n2 a_20121_n2241.n1 9.3005
R2538 a_2130_n21176.t0 a_2130_n21176.t1 82.0028
R2539 a_24530_n21342.t0 a_24530_n21342.t1 81.9492
R2540 standby_33.n0 standby_33.t0 227.886
R2541 standby_33 standby_33.t3 216.05
R2542 standby_33.n0 standby_33.n1 25.0903
R2543 standby_33.n0 standby_33.t4 12.7763
R2544 standby_33.n1 standby_33.t2 5.5105
R2545 standby_33.n1 standby_33.t1 5.5105
R2546 standby_33.n0 standby_33 1.67737
R2547 ibias.n7 ibias.n1 1544.9
R2548 ibias.n4 ibias.n3 1544.9
R2549 ibias.n2 ibias.n0 300.425
R2550 ibias.n8 ibias.n2 300.425
R2551 ibias.n9 ibias.n0 177.746
R2552 ibias.n9 ibias.n8 177.746
R2553 ibias.n5 ibias.n1 139.143
R2554 ibias.n6 ibias.n3 139.143
R2555 ibias.n9 ibias.t1 60.1061
R2556 ibias.n4 ibias.n0 46.2505
R2557 ibias.n8 ibias.n7 46.2505
R2558 ibias.n5 ibias.n4 40.8622
R2559 ibias.n7 ibias.n6 40.8622
R2560 ibias.n3 ibias.n2 12.3338
R2561 ibias.n9 ibias.n1 12.3338
R2562 ibias.n6 ibias.t0 4.16651
R2563 ibias.t0 ibias.n5 4.16651
R2564 ibias ibias.n9 1.58676
R2565 a_10658_n5446.t10 a_10658_n5446.n0 64.1378
R2566 a_10658_n5446.n0 a_10658_n5446.t13 31.8313
R2567 a_10658_n5446.t6 a_10658_n5446.n0 31.4637
R2568 a_10658_n5446.n0 a_10658_n5446.t2 31.4635
R2569 a_10658_n5446.t12 a_10658_n5446.n0 31.5048
R2570 a_10658_n5446.n0 a_10658_n5446.t7 40.9588
R2571 a_10658_n5446.n0 a_10658_n5446.t3 40.9588
R2572 a_10658_n5446.n0 a_10658_n5446.t1 40.9588
R2573 a_10658_n5446.n0 a_10658_n5446.t9 40.9588
R2574 a_10658_n5446.n0 a_10658_n5446.t5 40.9588
R2575 a_10658_n5446.n0 a_10658_n5446.t0 32.5193
R2576 a_10658_n5446.n0 a_10658_n5446.t11 31.8633
R2577 a_10658_n5446.n0 a_10658_n5446.t8 31.4953
R2578 a_10658_n5446.n0 a_10658_n5446.t4 31.4953
R2579 avdd_ip.n59 avdd_ip.n5 58547.9
R2580 avdd_ip.n61 avdd_ip.n5 58547.9
R2581 avdd_ip.n60 avdd_ip.n59 58547.9
R2582 avdd_ip.n61 avdd_ip.n60 58547.9
R2583 avdd_ip.n83 avdd_ip.n82 50887.3
R2584 avdd_ip.n58 avdd_ip.n3 28978.4
R2585 avdd_ip.n62 avdd_ip.n3 28978.4
R2586 avdd_ip.n58 avdd_ip.n4 28978.4
R2587 avdd_ip.n62 avdd_ip.n4 28978.4
R2588 avdd_ip.n53 avdd_ip.n45 7296
R2589 avdd_ip.n51 avdd_ip.n45 7296
R2590 avdd_ip.n53 avdd_ip.n46 7296
R2591 avdd_ip.n51 avdd_ip.n46 7296
R2592 avdd_ip.n63 avdd_ip.n2 6735.06
R2593 avdd_ip.n57 avdd_ip.n2 6735.06
R2594 avdd_ip.n57 avdd_ip.n56 3209.98
R2595 avdd_ip.n92 avdd_ip.n63 2921.68
R2596 avdd_ip.n85 avdd_ip.n84 857.648
R2597 avdd_ip.n87 avdd_ip.n79 857.648
R2598 avdd_ip.n84 avdd_ip.n79 857.648
R2599 avdd_ip.n73 avdd_ip.n66 857.648
R2600 avdd_ip.n70 avdd_ip.n67 857.648
R2601 avdd_ip.n83 avdd_ip.t2 337.433
R2602 avdd_ip.n71 avdd_ip.n70 267.182
R2603 avdd_ip.n73 avdd_ip.n72 267.182
R2604 avdd_ip.n87 avdd_ip.n86 267.182
R2605 avdd_ip.n47 avdd_ip.n1 212.464
R2606 avdd_ip.n50 avdd_ip.n49 203.02
R2607 avdd_ip.n93 avdd_ip.n1 201.294
R2608 avdd_ip.n49 avdd_ip.n6 134.407
R2609 avdd_ip.n56 avdd_ip.n6 110.358
R2610 avdd_ip.t7 avdd_ip.n45 105.665
R2611 avdd_ip.t11 avdd_ip.n46 105.665
R2612 avdd_ip.n70 avdd_ip.n69 92.5005
R2613 avdd_ip.n66 avdd_ip.n65 92.5005
R2614 avdd_ip.n74 avdd_ip.n73 92.5005
R2615 avdd_ip.n68 avdd_ip.n67 92.5005
R2616 avdd_ip.n84 avdd_ip.n81 92.5005
R2617 avdd_ip.n84 avdd_ip.n83 92.5005
R2618 avdd_ip.n80 avdd_ip.n79 92.5005
R2619 avdd_ip.t2 avdd_ip.n79 92.5005
R2620 avdd_ip.n88 avdd_ip.n87 92.5005
R2621 avdd_ip.n85 avdd_ip.n78 92.5005
R2622 avdd_ip.n69 avdd_ip.n65 91.4872
R2623 avdd_ip.n81 avdd_ip.n78 91.4829
R2624 avdd_ip.n52 avdd_ip.t7 79.5673
R2625 avdd_ip.n52 avdd_ip.t11 79.5673
R2626 avdd_ip.n93 avdd_ip.n92 75.3225
R2627 avdd_ip.n69 avdd_ip.n68 66.8331
R2628 avdd_ip.n81 avdd_ip.n80 66.3131
R2629 avdd_ip.n75 avdd_ip.n65 63.936
R2630 avdd_ip.n89 avdd_ip.n78 63.936
R2631 avdd_ip.n15 avdd_ip.t1 61.8276
R2632 avdd_ip.n33 avdd_ip.t24 61.1199
R2633 avdd_ip.n30 avdd_ip.t23 61.0882
R2634 avdd_ip.n31 avdd_ip.t25 60.1061
R2635 avdd_ip.n29 avdd_ip.t21 60.1061
R2636 avdd_ip.n7 avdd_ip.t20 60.1061
R2637 avdd_ip.n49 avdd_ip.t15 60.1061
R2638 avdd_ip.n49 avdd_ip.t12 60.1061
R2639 avdd_ip.n49 avdd_ip.t13 60.1061
R2640 avdd_ip.n47 avdd_ip.t10 60.1061
R2641 avdd_ip.n47 avdd_ip.t8 60.1061
R2642 avdd_ip.n47 avdd_ip.t9 60.1061
R2643 avdd_ip.n38 avdd_ip.t16 60.1061
R2644 avdd_ip.n38 avdd_ip.t14 60.1061
R2645 avdd_ip.n37 avdd_ip.t18 60.1061
R2646 avdd_ip.n37 avdd_ip.t17 60.1061
R2647 avdd_ip.n11 avdd_ip.t27 60.1061
R2648 avdd_ip.n11 avdd_ip.t19 60.1061
R2649 avdd_ip.n10 avdd_ip.t28 60.1061
R2650 avdd_ip.n10 avdd_ip.t22 60.1061
R2651 avdd_ip.n32 avdd_ip.t26 60.1061
R2652 avdd_ip.n86 avdd_ip.n85 57.4849
R2653 avdd_ip.n71 avdd_ip.n66 57.4849
R2654 avdd_ip.n72 avdd_ip.n67 57.4849
R2655 avdd_ip.n16 avdd_ip.n14 55.1707
R2656 avdd_ip.n16 avdd_ip.n13 54.9038
R2657 avdd_ip.n42 avdd_ip.n9 44.6614
R2658 avdd_ip.n74 avdd_ip.n64 43.3376
R2659 avdd_ip.n88 avdd_ip.n77 43.3376
R2660 avdd_ip.n44 avdd_ip.n43 30.1747
R2661 avdd_ip.n72 avdd_ip.t4 28.8172
R2662 avdd_ip.t4 avdd_ip.n71 28.8172
R2663 avdd_ip.n86 avdd_ip.t2 28.8172
R2664 avdd_ip.n50 avdd_ip.n47 10.9739
R2665 avdd_ip.n26 avdd_ip.n8 9.3005
R2666 avdd_ip.n56 avdd_ip.n55 8.37369
R2667 avdd_ip.n29 avdd_ip.n7 7.25561
R2668 avdd_ip.n32 avdd_ip.n31 7.25561
R2669 avdd_ip.n13 avdd_ip.t5 6.92425
R2670 avdd_ip.n13 avdd_ip.t3 6.92425
R2671 avdd_ip.n14 avdd_ip.t0 6.92425
R2672 avdd_ip.n14 avdd_ip.t6 6.92425
R2673 avdd_ip.n51 avdd_ip.n50 6.37981
R2674 avdd_ip.n52 avdd_ip.n51 6.37981
R2675 avdd_ip.n54 avdd_ip.n53 6.37981
R2676 avdd_ip.n53 avdd_ip.n52 6.37981
R2677 avdd_ip.n55 avdd_ip.n54 5.31953
R2678 avdd_ip.n68 avdd_ip.n64 4.38907
R2679 avdd_ip.n80 avdd_ip.n77 4.38907
R2680 avdd_ip.n54 avdd_ip.n8 3.70667
R2681 avdd_ip.n43 avdd_ip.n1 3.6009
R2682 avdd_ip.n90 avdd_ip.n77 2.4925
R2683 avdd_ip.n76 avdd_ip.n64 2.44611
R2684 avdd_ip.n46 avdd_ip.n6 2.43471
R2685 avdd_ip.n45 avdd_ip.n44 2.43471
R2686 avdd_ip.n75 avdd_ip.n74 2.37764
R2687 avdd_ip.n89 avdd_ip.n88 2.37764
R2688 avdd_ip.n76 avdd_ip.n75 2.3255
R2689 avdd_ip.n90 avdd_ip.n89 2.3255
R2690 avdd_ip avdd_ip.n93 2.08167
R2691 avdd_ip.n27 avdd_ip.n9 1.57905
R2692 avdd_ip.n18 avdd_ip.n17 1.18871
R2693 avdd_ip.n4 avdd_ip.n2 1.05764
R2694 avdd_ip.n60 avdd_ip.n4 1.05764
R2695 avdd_ip.n43 avdd_ip.n3 1.05764
R2696 avdd_ip.n5 avdd_ip.n3 1.05764
R2697 avdd_ip.n26 avdd_ip.n25 0.9903
R2698 avdd_ip.n30 avdd_ip.n29 0.919312
R2699 avdd_ip.n33 avdd_ip.n32 0.887629
R2700 avdd_ip.n25 avdd_ip.n18 0.827286
R2701 avdd_ip.n34 avdd_ip.n30 0.793513
R2702 avdd_ip.n49 avdd_ip.n48 0.793513
R2703 avdd_ip.n12 avdd_ip.n10 0.793513
R2704 avdd_ip.n39 avdd_ip.n37 0.793049
R2705 avdd_ip.n63 avdd_ip.n62 0.530586
R2706 avdd_ip.n62 avdd_ip.n61 0.530586
R2707 avdd_ip.n58 avdd_ip.n57 0.530586
R2708 avdd_ip.n59 avdd_ip.n58 0.530586
R2709 avdd_ip.n17 avdd_ip 0.502794
R2710 avdd_ip.n44 avdd_ip.n42 0.448948
R2711 avdd_ip.n40 avdd_ip.n39 0.373511
R2712 avdd_ip.n48 avdd_ip.n0 0.373046
R2713 avdd_ip.n36 avdd_ip.n12 0.373046
R2714 avdd_ip.n35 avdd_ip.n34 0.373046
R2715 avdd_ip.n48 avdd_ip.n47 0.282318
R2716 avdd_ip.n39 avdd_ip.n38 0.282318
R2717 avdd_ip.n12 avdd_ip.n11 0.282318
R2718 avdd_ip.n34 avdd_ip.n33 0.282318
R2719 avdd_ip.n16 avdd_ip.n15 0.267392
R2720 avdd_ip.n25 avdd_ip.n24 0.255087
R2721 avdd_ip.n35 avdd_ip.n28 0.245735
R2722 avdd_ip.n55 avdd_ip.n7 0.174542
R2723 avdd_ip.n31 avdd_ip.n9 0.174542
R2724 avdd_ip.n92 avdd_ip.n91 0.166571
R2725 avdd_ip.n36 avdd_ip.n35 0.150396
R2726 avdd_ip.n40 avdd_ip.n0 0.150396
R2727 avdd_ip.n17 avdd_ip.t33 0.125045
R2728 avdd_ip.n21 avdd_ip.n18 0.123905
R2729 avdd_ip.n41 avdd_ip.n40 0.117461
R2730 avdd_ip.n24 avdd_ip.n23 0.111971
R2731 avdd_ip.n22 avdd_ip.n21 0.110265
R2732 avdd_ip.n41 avdd_ip.n36 0.108384
R2733 avdd_ip.n20 avdd_ip.n19 0.106696
R2734 avdd_ip.n23 avdd_ip.n22 0.106696
R2735 avdd_ip.n91 avdd_ip.n76 0.0839309
R2736 avdd_ip.n91 avdd_ip.n90 0.0812962
R2737 avdd_ip.n15 avdd_ip 0.0511757
R2738 avdd_ip.n19 avdd_ip.t30 0.0180781
R2739 avdd_ip.n23 avdd_ip.t32 0.0180781
R2740 avdd_ip.n22 avdd_ip.t29 0.0180781
R2741 avdd_ip.n20 avdd_ip.t31 0.0180781
R2742 avdd_ip.n24 avdd_ip.n19 0.0174228
R2743 avdd_ip.n28 avdd_ip.n27 0.0173478
R2744 avdd_ip.n21 avdd_ip.n20 0.0150053
R2745 avdd_ip.n27 avdd_ip.n8 0.0119388
R2746 avdd_ip.n42 avdd_ip.n41 0.0117727
R2747 avdd_ip avdd_ip.n0 0.0112624
R2748 avdd_ip avdd_ip.n16 0.0055
R2749 avdd_ip.n28 avdd_ip.n26 0.000627812
R2750 xout.n35 xout.t26 594.784
R2751 xout.n35 xout.t24 194.649
R2752 xout.t23 xout.n29 86.3125
R2753 xout.n30 xout.t23 86.3125
R2754 xout.t25 xout.n27 86.3125
R2755 xout.n31 xout.t25 86.3125
R2756 xout.n3 xout.t16 60.5632
R2757 xout.n4 xout.t14 60.5632
R2758 xout.n5 xout.t21 60.1061
R2759 xout.n6 xout.t22 60.1061
R2760 xout.n12 xout.t12 60.1061
R2761 xout.n12 xout.t11 60.1061
R2762 xout.n14 xout.t15 60.1061
R2763 xout.n14 xout.t13 60.1061
R2764 xout.n0 xout.t18 60.1061
R2765 xout.n0 xout.t20 60.1061
R2766 xout.n1 xout.t17 60.1061
R2767 xout.n1 xout.t19 60.1061
R2768 xout.n31 xout.n30 58.6245
R2769 xout.n29 xout.n27 58.6245
R2770 xout.n26 xout.t1 43.5339
R2771 xout.n34 xout.n33 21.3269
R2772 xout.n20 xout.n19 18.5533
R2773 xout.n24 xout.n17 18.553
R2774 xout.n23 xout.n22 18.4723
R2775 xout.n23 xout.n21 18.4564
R2776 xout.n20 xout.n18 18.4564
R2777 xout.n33 xout.n27 12.2455
R2778 xout.n32 xout.n31 11.1505
R2779 xout.n22 xout.t5 4.133
R2780 xout.n22 xout.t3 4.133
R2781 xout.n21 xout.t10 4.133
R2782 xout.n21 xout.t2 4.133
R2783 xout.n19 xout.t8 4.133
R2784 xout.n19 xout.t0 4.133
R2785 xout.n18 xout.t9 4.133
R2786 xout.n18 xout.t4 4.133
R2787 xout.n17 xout.t6 4.133
R2788 xout.n17 xout.t7 4.133
R2789 xout.n7 xout.n5 3.62822
R2790 xout.n7 xout.n6 3.62822
R2791 xout.n29 xout.n28 3.26098
R2792 xout.n30 xout.n28 2.3255
R2793 xout.n26 xout.n25 2.24362
R2794 xout.n35 xout.n34 2.18092
R2795 xout.n34 xout.n26 1.03102
R2796 xout.n32 xout.n28 0.546796
R2797 xout xout.n35 0.527063
R2798 xout.n15 xout.n13 0.511695
R2799 xout.n2 xout.n0 0.478991
R2800 xout.n33 xout.n32 0.470755
R2801 xout.n25 xout.n16 0.464586
R2802 xout.n5 xout.n3 0.44563
R2803 xout.n6 xout.n4 0.44563
R2804 xout.n2 xout.n1 0.344956
R2805 xout.n10 xout.n2 0.310704
R2806 xout.n15 xout.n14 0.282318
R2807 xout.n13 xout.n12 0.282318
R2808 xout.n16 xout.n11 0.273717
R2809 xout.n11 xout.n10 0.261913
R2810 xout.n8 xout.n4 0.247581
R2811 xout.n9 xout.n3 0.247391
R2812 xout.n8 xout.n7 0.233
R2813 xout.n16 xout.n15 0.126542
R2814 xout.n13 xout.n11 0.1255
R2815 xout.n25 xout.n24 0.0947164
R2816 xout.n24 xout.n20 0.0657574
R2817 xout.n10 xout.n9 0.0505
R2818 xout.n24 xout.n23 0.0480746
R2819 xout.n9 xout.n8 0.00068997
R2820 inv_in.n19 inv_in.t0 45.9706
R2821 inv_in.n18 inv_in.t3 6.48745
R2822 inv_in.n19 inv_in.t1 6.24255
R2823 inv_in inv_in.n17 2.2182
R2824 inv_in.n18 inv_in 0.342687
R2825 inv_in inv_in.n18 0.217687
R2826 inv_in.n5 inv_in.n4 0.110198
R2827 inv_in.n7 inv_in.n6 0.110101
R2828 inv_in.n10 inv_in.n9 0.110101
R2829 inv_in.n8 inv_in.n2 0.110101
R2830 inv_in.n16 inv_in.n15 0.109734
R2831 inv_in.n14 inv_in.n0 0.109734
R2832 inv_in.n13 inv_in.n12 0.109709
R2833 inv_in.n11 inv_in.n1 0.109709
R2834 inv_in.n9 inv_in.n7 0.109325
R2835 inv_in.n9 inv_in.n8 0.109325
R2836 inv_in.n12 inv_in.n11 0.109325
R2837 inv_in.n11 inv_in.n3 0.109325
R2838 inv_in.n15 inv_in.n14 0.1086
R2839 inv_in.n16 inv_in.n0 0.1086
R2840 inv_in.n4 inv_in.n3 0.10222
R2841 inv_in.n7 inv_in.n5 0.101755
R2842 inv_in inv_in.n19 0.09425
R2843 inv_in.n18 inv_in 0.063
R2844 inv_in.n0 inv_in.t11 0.00880157
R2845 inv_in.n7 inv_in.t9 0.00848368
R2846 inv_in.n9 inv_in.t10 0.00848368
R2847 inv_in.n8 inv_in.t2 0.00848368
R2848 inv_in.n5 inv_in.t12 0.00838586
R2849 inv_in.n4 inv_in.t14 0.0083125
R2850 inv_in.n6 inv_in.t13 0.0083125
R2851 inv_in.n2 inv_in.t6 0.0083125
R2852 inv_in.n10 inv_in.t4 0.0083125
R2853 inv_in.n1 inv_in.t5 0.0083125
R2854 inv_in.n13 inv_in.t8 0.0083125
R2855 inv_in.n17 inv_in.t7 0.0083125
R2856 inv_in.n6 inv_in.n3 0.00106244
R2857 inv_in.n12 inv_in.n2 0.00106244
R2858 inv_in.n11 inv_in.n10 0.00106244
R2859 inv_in.n17 inv_in.n16 0.000989074
R2860 inv_in.n15 inv_in.n1 0.000548907
R2861 inv_in.n14 inv_in.n13 0.000548907
R2862 inv_m1.t0 inv_m1.n8 651.431
R2863 inv_m1 inv_m1.n7 0.00675
R2864 inv_m1.n7 inv_m1.n8 0.0451429
R2865 inv_m1.n8 inv_m1.n6 0.0451429
R2866 inv_m1 inv_m1.n7 0.893357
R2867 inv_m1 inv_m1.n6 0.13425
R2868 inv_m1.n6 inv_m1.n0 0.60925
R2869 inv_m1.n0 inv_m1.n5 0.533
R2870 inv_m1 inv_m1.n5 1.063
R2871 inv_m1.n5 inv_m1.n4 0.0525833
R2872 inv_m1 inv_m1.n4 1.45258
R2873 inv_m1.n4 inv_m1.t1 229.101
R2874 inv_m1.n0 inv_m1.n3 5.613
R2875 inv_m1.n3 inv_m1.n2 24.8426
R2876 inv_m1.n2 inv_m1.t4 20.438
R2877 inv_m1.n2 inv_m1.t3 20.4375
R2878 inv_m1.n3 inv_m1.n1 24.7082
R2879 inv_m1.n1 inv_m1.t5 21.9207
R2880 inv_m1.n1 inv_m1.t2 21.9202
R2881 a_2132_n15590.t0 a_2132_n15590.t1 82.3309
R2882 a_18932_n15756.t0 a_18932_n15756.t1 83.5579
R2883 inv_m2 inv_m2.t0 651.431
R2884 inv_m2 inv_m2.t1 229.101
R2885 inv_m2 inv_m2.n1 24.0208
R2886 inv_m2 inv_m2.n0 23.8727
R2887 inv_m2.n0 inv_m2.t5 21.9784
R2888 inv_m2.n0 inv_m2.t2 21.8626
R2889 inv_m2.n1 inv_m2.t3 20.4885
R2890 inv_m2.n1 inv_m2.t4 20.387
R2891 dout_ip dout_ip.t0 651.431
R2892 dout_ip dout_ip.t1 651.431
R2893 dout_ip.n0 dout_ip.t10 288.204
R2894 dout_ip.n4 dout_ip.t6 264.103
R2895 dout_ip.n1 dout_ip.t7 264.103
R2896 dout_ip dout_ip.t4 230.433
R2897 dout_ip dout_ip.t3 229.15
R2898 dout_ip dout_ip.t2 229.101
R2899 dout_ip.n0 dout_ip.t8 195.017
R2900 dout_ip dout_ip.n4 159.236
R2901 dout_ip dout_ip.n1 159.236
R2902 dout_ip dout_ip.n0 153.153
R2903 dout_ip.n3 dout_ip 152
R2904 dout_ip dout_ip.n2 152
R2905 dout_ip.n3 dout_ip.t9 145.209
R2906 dout_ip.n2 dout_ip.t5 145.209
R2907 dout_ip.n6 dout_ip.n5 117.519
R2908 dout_ip.n5 dout_ip 68.1959
R2909 dout_ip.n4 dout_ip.n3 37.6741
R2910 dout_ip.n2 dout_ip.n1 37.6741
R2911 dout_ip dout_ip.n6 31.6505
R2912 dout_ip.n6 dout_ip 24.4485
R2913 dout_ip.n5 dout_ip 9.3005
R2914 a_20689_n2549.n3 a_20689_n2549.n2 647.119
R2915 a_20689_n2549.n1 a_20689_n2549.t4 350.253
R2916 a_20689_n2549.n2 a_20689_n2549.n0 260.339
R2917 a_20689_n2549.n2 a_20689_n2549.n1 246.119
R2918 a_20689_n2549.n1 a_20689_n2549.t5 189.588
R2919 a_20689_n2549.n3 a_20689_n2549.t3 89.1195
R2920 a_20689_n2549.n0 a_20689_n2549.t2 63.3338
R2921 a_20689_n2549.t0 a_20689_n2549.n3 41.0422
R2922 a_20689_n2549.n0 a_20689_n2549.t1 31.9797
R2923 a_20567_n2791.t0 a_20567_n2791.t1 198.571
R2924 a_20733_n2791.t0 a_20733_n2791.t1 60.0005
R2925 a_17576_n6897.n0 a_17576_n6897.t3 3.48032
R2926 a_17576_n6897.t0 a_17576_n6897.n0 27.3396
R2927 a_17576_n6897.t4 a_17576_n6897.n0 9.97518
R2928 a_17576_n6897.t0 a_17576_n6897.n1 8.84728
R2929 a_17576_n6897.n1 a_17576_n6897.t2 6.06443
R2930 a_17576_n6897.n1 a_17576_n6897.t1 2.20565
R2931 a_15000_n1881.n2 a_15000_n1881.n1 682.193
R2932 a_15000_n1881.n0 a_15000_n1881.t4 279.142
R2933 a_15000_n1881.n1 a_15000_n1881.t1 250.737
R2934 a_15000_n1881.n0 a_15000_n1881.t3 145.958
R2935 a_15000_n1881.n1 a_15000_n1881.n0 118.45
R2936 a_15000_n1881.t0 a_15000_n1881.n2 70.3576
R2937 a_15000_n1881.n2 a_15000_n1881.t2 65.6672
R2938 x7.x1.x2.CLK x7.x1.x2.CLK.t0 716.451
R2939 x7.x1.x2.CLK.t0 x7.x1.x2.CLK.n3 707.66
R2940 x7.x1.x2.CLK.n0 x7.x1.x2.CLK.t2 294.557
R2941 x7.x1.x2.CLK.n2 x7.x1.x2.CLK.t1 271.777
R2942 x7.x1.x2.CLK.n0 x7.x1.x2.CLK.t3 211.01
R2943 x7.x1.x2.CLK.n1 x7.x1.x2.CLK.n0 152
R2944 x7.x1.x2.CLK.n3 x7.x1.x2.CLK.n2 38.2982
R2945 x7.x1.x2.CLK.n2 x7.x1.x2.CLK.n1 33.0611
R2946 x7.x1.x2.CLK x7.x1.x2.CLK.n3 8.88521
R2947 x7.x1.x2.CLK.n1 x7.x1.x2.CLK 4.20621
R2948 a_16151_n1869.t0 a_16151_n1869.t1 198.571
R2949 a_16317_n1881.t0 a_16317_n1881.t1 60.0005
R2950 a_21775_n2791.t1 a_21775_n2791.n1 386.31
R2951 a_21775_n2791.n1 a_21775_n2791.t0 249.956
R2952 a_21775_n2791.n0 a_21775_n2791.t3 239.04
R2953 a_21775_n2791.n1 a_21775_n2791.n0 175.661
R2954 a_21775_n2791.n0 a_21775_n2791.t2 166.739
R2955 x7.x5.TE_B.n3 x7.x5.TE_B.t0 319.219
R2956 x7.x5.TE_B.n1 x7.x5.TE_B.t4 268.313
R2957 x7.x5.TE_B x7.x5.TE_B.t1 249.867
R2958 x7.x5.TE_B.n2 x7.x5.TE_B.t2 206.19
R2959 x7.x5.TE_B.n1 x7.x5.TE_B.t5 186.374
R2960 x7.x5.TE_B x7.x5.TE_B.n2 152
R2961 x7.x5.TE_B.n2 x7.x5.TE_B.n1 148.35
R2962 x7.x5.TE_B x7.x5.TE_B.t3 38.3302
R2963 x7.x5.TE_B x7.x5.TE_B.n0 32.2121
R2964 x7.x5.TE_B.n3 x7.x5.TE_B 21.8175
R2965 x7.x5.TE_B.n0 x7.x5.TE_B 11.0708
R2966 x7.x5.TE_B.n0 x7.x5.TE_B 8.03187
R2967 x7.x5.TE_B x7.x5.TE_B.n3 4.14393
R2968 a_14009_n2701.t0 a_14009_n2701.n0 753.673
R2969 a_14009_n2701.n0 a_14009_n2701.t2 354.81
R2970 a_14009_n2701.n0 a_14009_n2701.t1 303.562
R2971 standby_ip.t1 standby_ip.n4 368.26
R2972 standby_ip.n3 standby_ip.n4 1.85916
R2973 standby_ip.t15 standby_ip.n22 381.469
R2974 standby_ip.n25 standby_ip.t15 381.462
R2975 standby_ip.t6 standby_ip.n17 375.649
R2976 standby_ip.n32 standby_ip.t6 375.649
R2977 standby_ip.n19 standby_ip.t17 375.649
R2978 standby_ip.t17 standby_ip.n7 375.649
R2979 standby_ip.t18 standby_ip.n30 375.649
R2980 standby_ip.n31 standby_ip.t18 375.649
R2981 standby_ip.n11 standby_ip.t5 375.649
R2982 standby_ip.t5 standby_ip.n18 375.649
R2983 standby_ip.n29 standby_ip.t11 375.649
R2984 standby_ip.t11 standby_ip.n28 375.649
R2985 standby_ip.t12 standby_ip.n20 375.649
R2986 standby_ip.n21 standby_ip.t12 375.649
R2987 standby_ip.t8 standby_ip.n26 375.649
R2988 standby_ip.n27 standby_ip.t8 375.649
R2989 standby_ip.n24 standby_ip.t9 375.649
R2990 standby_ip.t9 standby_ip.n23 375.649
R2991 standby_ip.t13 standby_ip.n33 332.752
R2992 standby_ip.n34 standby_ip.t13 332.75
R2993 standby_ip.t7 standby_ip.n33 332.411
R2994 standby_ip.n34 standby_ip.t7 332.411
R2995 standby_ip.n15 standby_ip.t3 231.718
R2996 standby_ip standby_ip.t0 216.155
R2997 standby_ip standby_ip.n16 161.314
R2998 standby_ip.n15 standby_ip.t14 159.417
R2999 standby_ip.n16 standby_ip.n15 152
R3000 standby_ip.n2 standby_ip.t16 59.9857
R3001 standby_ip standby_ip.t2 59.3654
R3002 standby_ip standby_ip.n3 46.2227
R3003 standby_ip.n27 standby_ip.n23 29.7417
R3004 standby_ip.n27 standby_ip.n5 5.72268
R3005 standby_ip.n28 standby_ip.n21 29.7417
R3006 standby_ip.n6 standby_ip.n18 5.72268
R3007 standby_ip.n31 standby_ip.n18 29.7417
R3008 standby_ip.n8 standby_ip.n7 5.72268
R3009 standby_ip.n32 standby_ip.n7 29.7417
R3010 standby_ip.t4 standby_ip.n9 381.37
R3011 standby_ip.n26 standby_ip.n24 29.7417
R3012 standby_ip.n26 standby_ip.n10 5.72268
R3013 standby_ip.n29 standby_ip.n20 29.7417
R3014 standby_ip.n12 standby_ip.n11 5.72268
R3015 standby_ip.n30 standby_ip.n11 29.7417
R3016 standby_ip.n13 standby_ip.n19 5.72268
R3017 standby_ip.n19 standby_ip.n17 29.7417
R3018 standby_ip.t4 standby_ip.n14 381.37
R3019 standby_ip.n0 standby_ip 13.0593
R3020 standby_ip standby_ip.t10 12.6603
R3021 standby_ip.n1 standby_ip.n5 1.79016
R3022 standby_ip.n5 standby_ip.n21 5.72268
R3023 standby_ip.n28 standby_ip.n6 5.72268
R3024 standby_ip.n6 standby_ip.n1 1.79016
R3025 standby_ip.n8 standby_ip.n31 5.72268
R3026 standby_ip.n1 standby_ip.n8 1.79016
R3027 standby_ip.n32 standby_ip.n9 5.72268
R3028 standby_ip.n20 standby_ip.n10 5.72268
R3029 standby_ip.n12 standby_ip.n29 5.72268
R3030 standby_ip.n0 standby_ip.n12 1.79016
R3031 standby_ip.n30 standby_ip.n13 5.72268
R3032 standby_ip.n0 standby_ip.n13 1.79016
R3033 standby_ip.n17 standby_ip.n14 5.72268
R3034 standby_ip.n0 standby_ip.n14 1.79016
R3035 standby_ip standby_ip.n36 9.27339
R3036 standby_ip standby_ip.n0 7.693
R3037 standby_ip.n25 standby_ip.n24 5.70112
R3038 standby_ip.n23 standby_ip.n22 5.6994
R3039 standby_ip.n35 standby_ip.n33 5.53161
R3040 standby_ip.n36 standby_ip.n3 5.46183
R3041 standby_ip.n35 standby_ip.n34 4.67076
R3042 standby_ip.n4 standby_ip 1.88798
R3043 standby_ip.n2 standby_ip.n35 3.51723
R3044 standby_ip.n10 standby_ip.n0 3.39911
R3045 standby_ip.n9 standby_ip.n1 3.17266
R3046 standby_ip.n3 standby_ip 2.98717
R3047 standby_ip.n16 standby_ip 2.74336
R3048 standby_ip.n0 standby_ip.n1 2.40496
R3049 standby_ip.n1 standby_ip.n22 2.01822
R3050 standby_ip.n0 standby_ip.n25 2.00133
R3051 standby_ip.n36 standby_ip 1.8605
R3052 standby_ip standby_ip.n2 1.82266
R3053 a_2971_n1521.t1 a_2971_n1521.n1 405.735
R3054 a_2971_n1521.n1 a_2971_n1521.t0 294.611
R3055 a_2971_n1521.n0 a_2971_n1521.t3 254.389
R3056 a_2971_n1521.n0 a_2971_n1521.t2 211.01
R3057 a_2971_n1521.n1 a_2971_n1521.n0 152
R3058 a_14035_n1997.t0 a_14035_n1997.t1 38.7697
R3059 a_2132_n17582.t0 a_2132_n17582.t1 83.9053
R3060 a_18932_n17416.t0 a_18932_n17416.t1 83.5579
R3061 avss.n20 avss.n19 18715.6
R3062 avss.n38 avss.n37 15510.3
R3063 avss.n75 avss.n20 12243.6
R3064 avss.n39 avss.n33 3599.36
R3065 avss.n40 avss.n33 3599.36
R3066 avss.n40 avss.n35 3599.36
R3067 avss.n39 avss.n35 3599.36
R3068 avss.n66 avss.n25 2489.59
R3069 avss.n66 avss.n26 2489.59
R3070 avss.n68 avss.n26 2489.59
R3071 avss.n68 avss.n25 2489.59
R3072 avss.n28 avss.n21 2489.59
R3073 avss.n28 avss.n22 2489.59
R3074 avss.n73 avss.n22 2489.59
R3075 avss.n73 avss.n21 2489.59
R3076 avss.n77 avss.n13 2489.59
R3077 avss.n77 avss.n14 2489.59
R3078 avss.n16 avss.n14 2489.59
R3079 avss.n16 avss.n13 2489.59
R3080 avss.n87 avss.n6 2489.59
R3081 avss.n89 avss.n6 2489.59
R3082 avss.n89 avss.n5 2489.59
R3083 avss.n87 avss.n5 2489.59
R3084 avss.n36 avss.n20 2350.09
R3085 avss.n76 avss.n75 928.033
R3086 avss.n75 avss.n74 928.033
R3087 avss.n19 avss.t24 631.537
R3088 avss.n15 avss.t22 631.537
R3089 avss.t10 avss.n17 631.537
R3090 avss.n76 avss.t12 631.537
R3091 avss.n74 avss.t16 631.537
R3092 avss.n29 avss.t18 631.537
R3093 avss.t0 avss.n30 631.537
R3094 avss.n37 avss.t2 631.537
R3095 avss.n42 avss.n32 499.257
R3096 avss.n42 avss.n41 499.257
R3097 avss.n34 avss.n32 416
R3098 avss.n41 avss.n34 416
R3099 avss.t20 avss.n36 413.959
R3100 avss.t6 avss.n38 390.637
R3101 avss.n17 avss.n15 361.726
R3102 avss.n30 avss.n29 361.726
R3103 avss.t14 avss.t20 307.067
R3104 avss.t8 avss.t14 307.067
R3105 avss.t8 avss.t4 307.067
R3106 avss.t4 avss.t6 307.067
R3107 avss.n65 avss.n64 289.13
R3108 avss.n86 avss.n3 289.13
R3109 avss.n91 avss.n90 288.753
R3110 avss.n69 avss.n24 288.753
R3111 avss.n88 avss.t24 234.232
R3112 avss.n88 avss.t22 234.232
R3113 avss.n18 avss.t10 234.232
R3114 avss.t12 avss.n18 234.232
R3115 avss.n27 avss.t16 234.232
R3116 avss.t18 avss.n27 234.232
R3117 avss.n67 avss.t0 234.232
R3118 avss.n67 avss.t2 234.232
R3119 avss.n31 avss.n10 152.73
R3120 avss.n72 avss.n71 152.73
R3121 avss.n79 avss.n7 152.73
R3122 avss.n78 avss.n12 152.73
R3123 avss.n90 avss.n4 103.529
R3124 avss.n63 avss.n31 103.529
R3125 avss.n71 avss.n70 103.529
R3126 avss.n65 avss.n63 103.529
R3127 avss.n70 avss.n69 103.529
R3128 avss.n85 avss.n7 103.529
R3129 avss.n12 avss.n4 103.529
R3130 avss.n86 avss.n85 103.529
R3131 avss.n87 avss.n86 97.5005
R3132 avss.n88 avss.n87 97.5005
R3133 avss.n90 avss.n89 97.5005
R3134 avss.n89 avss.n88 97.5005
R3135 avss.n13 avss.n7 97.5005
R3136 avss.n18 avss.n13 97.5005
R3137 avss.n14 avss.n12 97.5005
R3138 avss.n18 avss.n14 97.5005
R3139 avss.n31 avss.n21 97.5005
R3140 avss.n27 avss.n21 97.5005
R3141 avss.n71 avss.n22 97.5005
R3142 avss.n27 avss.n22 97.5005
R3143 avss.n69 avss.n68 97.5005
R3144 avss.n68 avss.n67 97.5005
R3145 avss.n66 avss.n65 97.5005
R3146 avss.n67 avss.n66 97.5005
R3147 avss.n38 avss.n33 62.3221
R3148 avss.n5 avss.n3 48.7505
R3149 avss.n19 avss.n5 48.7505
R3150 avss.n8 avss.n6 48.7505
R3151 avss.n15 avss.n6 48.7505
R3152 avss.n16 avss.n8 48.7505
R3153 avss.n17 avss.n16 48.7505
R3154 avss.n78 avss.n77 48.7505
R3155 avss.n77 avss.n76 48.7505
R3156 avss.n73 avss.n72 48.7505
R3157 avss.n74 avss.n73 48.7505
R3158 avss.n28 avss.n23 48.7505
R3159 avss.n29 avss.n28 48.7505
R3160 avss.n25 avss.n23 48.7505
R3161 avss.n30 avss.n25 48.7505
R3162 avss.n64 avss.n26 48.7505
R3163 avss.n37 avss.n26 48.7505
R3164 avss.n39 avss.n32 45.0005
R3165 avss.t8 avss.n39 45.0005
R3166 avss.n41 avss.n40 45.0005
R3167 avss.n40 avss.t8 45.0005
R3168 avss.n63 avss.n62 40.3697
R3169 avss.n70 avss.n23 40.3697
R3170 avss.n85 avss.n84 40.3697
R3171 avss.n8 avss.n4 40.3697
R3172 avss.n93 avss.n1 39.7977
R3173 avss.n35 avss.n34 39.0005
R3174 avss.n36 avss.n35 39.0005
R3175 avss.n42 avss.n33 39.0005
R3176 avss.n93 avss 33.7505
R3177 avss.n83 avss.t11 29.9199
R3178 avss.n61 avss.t1 29.9199
R3179 avss.n61 avss.t19 29.9199
R3180 avss.n83 avss.t23 29.9199
R3181 avss.n2 avss.t25 29.798
R3182 avss.n56 avss.t3 29.798
R3183 avss.n11 avss.t13 29.798
R3184 avss.n11 avss.t17 29.798
R3185 avss.n42 avss.t7 20.9512
R3186 avss.n45 avss.n44 18.7295
R3187 avss.n45 avss.n43 18.5391
R3188 avss.n43 avss.t9 4.133
R3189 avss.n43 avss.t5 4.133
R3190 avss.n44 avss.t21 4.133
R3191 avss.n44 avss.t15 4.133
R3192 avss.n46 avss.n42 1.61679
R3193 avss.n54 avss 1.33946
R3194 avss.n57 avss.n24 1.21803
R3195 avss.n92 avss.n91 1.21803
R3196 avss.n53 avss.n46 0.8655
R3197 avss.n62 avss.n61 0.664786
R3198 avss.n80 avss.n10 0.664786
R3199 avss.n80 avss.n79 0.664786
R3200 avss.n84 avss.n83 0.664786
R3201 avss.n54 avss.n53 0.53175
R3202 avss.n55 avss.n9 0.434977
R3203 avss.n94 avss.n0 0.433066
R3204 avss.n60 avss.n58 0.433066
R3205 avss.n60 avss.n59 0.433066
R3206 avss.n59 avss.n0 0.433066
R3207 avss.n64 avss.n24 0.376971
R3208 avss.n91 avss.n3 0.376971
R3209 avss.n83 avss.n0 0.299413
R3210 avss.n61 avss.n60 0.299413
R3211 avss.n61 avss.n9 0.247783
R3212 avss.n83 avss.n82 0.247783
R3213 avss.n58 avss.n57 0.231236
R3214 avss.n82 avss 0.215995
R3215 avss.n81 avss.n9 0.201672
R3216 avss.n82 avss.n81 0.201672
R3217 avss.n2 avss.n1 0.2005
R3218 avss.n94 avss.n93 0.2005
R3219 avss.n46 avss.n45 0.1855
R3220 avss.n48 avss.n47 0.122162
R3221 avss.n81 avss.n80 0.120904
R3222 avss.n49 avss.n48 0.105544
R3223 avss.n50 avss.n49 0.101695
R3224 avss.n72 avss.n10 0.1005
R3225 avss.n79 avss.n78 0.1005
R3226 avss.n59 avss.n11 0.0997647
R3227 avss.n52 avss.n47 0.0989292
R3228 avss.n55 avss.n54 0.096886
R3229 avss.n53 avss.n52 0.0847138
R3230 avss.n62 avss.n23 0.0825513
R3231 avss.n84 avss.n8 0.0825513
R3232 avss.n50 avss.n47 0.0586846
R3233 avss.n56 avss.n55 0.0480171
R3234 avss avss.n1 0.0333776
R3235 avss avss.n94 0.0332586
R3236 avss.n58 avss 0.0330342
R3237 avss.n93 avss.n92 0.0328276
R3238 avss.n52 avss.n51 0.0277801
R3239 avss.n49 avss.t28 0.0083125
R3240 avss.n48 avss.t29 0.0083125
R3241 avss.n47 avss.t26 0.0083125
R3242 avss.n51 avss.t27 0.0083125
R3243 avss.n92 avss.n2 0.000931034
R3244 avss.n57 avss.n56 0.000928082
R3245 avss.n80 avss.n11 0.000683824
R3246 avss.n51 avss.n50 0.000622332
R3247 avdd.n92 avdd.n91 15787.9
R3248 avdd.n93 avdd.n92 15787.9
R3249 avdd.n93 avdd.n28 15787.9
R3250 avdd.n91 avdd.n28 15787.9
R3251 avdd.n90 avdd.n27 8103.24
R3252 avdd.n94 avdd.n27 8103.24
R3253 avdd.n94 avdd.n26 8103.24
R3254 avdd.n90 avdd.n26 8103.24
R3255 avdd.n98 avdd.n6 2166
R3256 avdd.n97 avdd.n6 2166
R3257 avdd.n98 avdd.n7 2166
R3258 avdd.n97 avdd.n7 2166
R3259 avdd.n66 avdd.n25 1699.15
R3260 avdd.n78 avdd.n77 1643.17
R3261 avdd.n77 avdd.n76 1643.17
R3262 avdd.n74 avdd.n69 1643.17
R3263 avdd.n80 avdd.n69 1643.17
R3264 avdd.n52 avdd.n37 1643.17
R3265 avdd.n60 avdd.n37 1643.17
R3266 avdd.n55 avdd.n54 1643.17
R3267 avdd.n58 avdd.n55 1643.17
R3268 avdd.n89 avdd.n29 1539.31
R3269 avdd.n89 avdd.n88 1532.98
R3270 avdd.n71 avdd.n70 1106.59
R3271 avdd.n70 avdd.n68 1106.59
R3272 avdd.n40 avdd.n39 1106.59
R3273 avdd.n39 avdd.n36 1106.59
R3274 avdd.n78 avdd.n68 536.587
R3275 avdd.n76 avdd.n71 536.587
R3276 avdd.n74 avdd.n71 536.587
R3277 avdd.n80 avdd.n68 536.587
R3278 avdd.n52 avdd.n40 536.587
R3279 avdd.n54 avdd.n40 536.587
R3280 avdd.n58 avdd.n36 536.587
R3281 avdd.n60 avdd.n36 536.587
R3282 avdd.n75 avdd.t4 382.582
R3283 avdd.n79 avdd.t4 382.582
R3284 avdd.n53 avdd.t0 382.582
R3285 avdd.n59 avdd.t0 382.582
R3286 avdd.n73 avdd.n30 319.248
R3287 avdd.n57 avdd.n56 319.248
R3288 avdd.n88 avdd.n31 287.265
R3289 avdd.n38 avdd.n29 287.265
R3290 avdd.n88 avdd.n30 276.295
R3291 avdd.n56 avdd.n29 276.295
R3292 avdd.n25 avdd.n4 263.788
R3293 avdd.n100 avdd.n4 253.528
R3294 avdd.n86 avdd.t19 227.377
R3295 avdd.n1 avdd.t5 227.377
R3296 avdd.n34 avdd.t1 227.377
R3297 avdd.n43 avdd.t12 227.377
R3298 avdd.n66 avdd.n3 205.554
R3299 avdd.n72 avdd.n31 189.742
R3300 avdd.n38 avdd.n35 189.742
R3301 avdd.n101 avdd.n3 186.73
R3302 avdd.t2 avdd.n6 157.492
R3303 avdd.t6 avdd.n7 157.492
R3304 avdd.n73 avdd.n72 108.569
R3305 avdd.n57 avdd.n35 108.569
R3306 avdd.t17 avdd.t2 107.677
R3307 avdd.t15 avdd.t17 107.677
R3308 avdd.t15 avdd.t13 107.677
R3309 avdd.t13 avdd.t6 107.677
R3310 avdd.n62 avdd.n5 63.4672
R3311 avdd.n23 avdd.t3 60.1061
R3312 avdd.n21 avdd.n20 54.9038
R3313 avdd.n21 avdd.n19 54.9038
R3314 avdd.n72 avdd.n2 32.2138
R3315 avdd.n61 avdd.n35 32.2138
R3316 avdd.n101 avdd.n100 31.7005
R3317 avdd.n102 avdd.n101 30.3938
R3318 avdd.n76 avdd.n73 26.4291
R3319 avdd.n76 avdd.n75 26.4291
R3320 avdd.n74 avdd.n2 26.4291
R3321 avdd.n75 avdd.n74 26.4291
R3322 avdd.n78 avdd.n32 26.4291
R3323 avdd.n79 avdd.n78 26.4291
R3324 avdd.n81 avdd.n80 26.4291
R3325 avdd.n80 avdd.n79 26.4291
R3326 avdd.n58 avdd.n57 26.4291
R3327 avdd.n59 avdd.n58 26.4291
R3328 avdd.n61 avdd.n60 26.4291
R3329 avdd.n60 avdd.n59 26.4291
R3330 avdd.n54 avdd.n41 26.4291
R3331 avdd.n54 avdd.n53 26.4291
R3332 avdd.n52 avdd.n51 26.4291
R3333 avdd.n53 avdd.n52 26.4291
R3334 avdd.n96 avdd.n24 15.7582
R3335 avdd.n97 avdd.n96 14.2313
R3336 avdd.t15 avdd.n97 14.2313
R3337 avdd.n99 avdd.n98 14.2313
R3338 avdd.n98 avdd.t15 14.2313
R3339 avdd.n77 avdd.n30 13.2148
R3340 avdd.n77 avdd.t4 13.2148
R3341 avdd.n70 avdd.n31 13.2148
R3342 avdd.n70 avdd.t4 13.2148
R3343 avdd.n69 avdd.n3 13.2148
R3344 avdd.t4 avdd.n69 13.2148
R3345 avdd.n39 avdd.n38 13.2148
R3346 avdd.n39 avdd.t0 13.2148
R3347 avdd.n56 avdd.n55 13.2148
R3348 avdd.n55 avdd.t0 13.2148
R3349 avdd.n49 avdd.n37 13.2148
R3350 avdd.t0 avdd.n37 13.2148
R3351 avdd.n7 avdd.n4 12.3338
R3352 avdd.n47 avdd.n6 12.3338
R3353 avdd.n100 avdd.n99 8.13132
R3354 avdd.n95 avdd.n25 7.55272
R3355 avdd.n82 avdd.n32 7.35838
R3356 avdd.n46 avdd.n41 7.25772
R3357 avdd.n20 avdd.t18 6.92425
R3358 avdd.n20 avdd.t16 6.92425
R3359 avdd.n19 avdd.t14 6.92425
R3360 avdd.n19 avdd.t7 6.92425
R3361 avdd.n48 avdd.n47 6.8963
R3362 avdd.n99 avdd.n5 6.16704
R3363 avdd.n67 avdd.n66 3.62858
R3364 avdd.n50 avdd.n49 3.40824
R3365 avdd.n82 avdd.n81 2.88262
R3366 avdd.n90 avdd.n89 2.84665
R3367 avdd.n91 avdd.n90 2.84665
R3368 avdd.n95 avdd.n94 2.84665
R3369 avdd.n94 avdd.n93 2.84665
R3370 avdd.n51 avdd.n46 2.79686
R3371 avdd.n48 avdd.n5 2.51338
R3372 avdd.n49 avdd.n48 2.33947
R3373 avdd.n67 avdd.n27 2.28445
R3374 avdd.n92 avdd.n27 2.28445
R3375 avdd.n50 avdd.n26 2.28445
R3376 avdd.n28 avdd.n26 2.28445
R3377 avdd.n84 avdd 1.89829
R3378 avdd.n23 avdd.n22 1.87575
R3379 avdd.n102 avdd.n2 1.70717
R3380 avdd.n62 avdd.n61 1.70717
R3381 avdd.n81 avdd.n67 1.49242
R3382 avdd.n51 avdd.n50 1.46526
R3383 avdd.n85 avdd.n1 1.11161
R3384 avdd.n96 avdd.n95 1.03039
R3385 avdd.n65 avdd.n33 0.909856
R3386 avdd.n87 avdd.n65 0.871595
R3387 avdd.n42 avdd.n29 0.517167
R3388 avdd.n63 avdd.n62 0.517167
R3389 avdd.n103 avdd.n102 0.517167
R3390 avdd.n88 avdd.n87 0.517167
R3391 avdd.n83 avdd.n1 0.457832
R3392 avdd.n88 avdd.n32 0.305666
R3393 avdd.n41 avdd.n29 0.30011
R3394 avdd.n44 avdd.n34 0.277965
R3395 avdd.n44 avdd.n43 0.242141
R3396 avdd.n13 avdd.n12 0.221624
R3397 avdd.n45 avdd.n44 0.191202
R3398 avdd.n15 avdd.n8 0.171
R3399 avdd.n64 avdd 0.165618
R3400 avdd.n18 avdd.n8 0.158572
R3401 avdd.n45 avdd.n33 0.155105
R3402 avdd.n22 avdd.n18 0.129984
R3403 avdd.n65 avdd.n64 0.124867
R3404 avdd.n24 avdd.n23 0.0960224
R3405 avdd.n18 avdd.n17 0.0860931
R3406 avdd.n16 avdd.n15 0.0718577
R3407 avdd.n15 avdd.n14 0.0677409
R3408 avdd.n46 avdd.n45 0.058264
R3409 avdd.n83 avdd.n82 0.058264
R3410 avdd.n86 avdd.n85 0.0482015
R3411 avdd avdd.n63 0.0421667
R3412 avdd avdd.n0 0.035342
R3413 avdd.n12 avdd.n0 0.0293462
R3414 avdd.n22 avdd.n21 0.0285269
R3415 avdd.n17 avdd.n16 0.0255438
R3416 avdd.n14 avdd.n13 0.0253723
R3417 avdd.n12 avdd.n8 0.0246031
R3418 avdd.n85 avdd.n84 0.0240664
R3419 avdd.n11 avdd.t10 0.0122401
R3420 avdd avdd.n103 0.0122337
R3421 avdd.n17 avdd.t8 0.0122173
R3422 avdd.n10 avdd.t11 0.0113908
R3423 avdd.n9 avdd.t9 0.011362
R3424 avdd.n63 avdd.n34 0.0105575
R3425 avdd.n103 avdd.n1 0.0105575
R3426 avdd.n17 avdd.n9 0.00991802
R3427 avdd.n11 avdd.n10 0.00930403
R3428 avdd.n47 avdd.n24 0.00806949
R3429 avdd.n64 avdd 0.00600766
R3430 avdd.n43 avdd.n42 0.00573256
R3431 avdd.n42 avdd.n33 0.00515116
R3432 avdd.n87 avdd.n86 0.00333375
R3433 avdd.n14 avdd.n9 0.00220261
R3434 avdd.n16 avdd.n10 0.00176706
R3435 avdd.n84 avdd.n83 0.00111075
R3436 avdd.n64 avdd.n0 0.00109866
R3437 avdd.n13 avdd.n11 0.000671533
R3438 a_10620_n9666.t0 a_10620_n9666.t1 83.9243
R3439 a_20567_n1869.t0 a_20567_n1869.t1 198.571
R3440 a_20733_n1881.t0 a_20733_n1881.t1 60.0005
R3441 a_15539_n2791.n1 a_15539_n2791.t6 530.01
R3442 a_15539_n2791.t0 a_15539_n2791.n5 421.021
R3443 a_15539_n2791.n0 a_15539_n2791.t5 337.142
R3444 a_15539_n2791.n3 a_15539_n2791.t1 280.223
R3445 a_15539_n2791.n4 a_15539_n2791.t2 263.173
R3446 a_15539_n2791.n4 a_15539_n2791.t4 227.826
R3447 a_15539_n2791.n0 a_15539_n2791.t7 199.762
R3448 a_15539_n2791.n2 a_15539_n2791.n1 170.81
R3449 a_15539_n2791.n2 a_15539_n2791.n0 167.321
R3450 a_15539_n2791.n5 a_15539_n2791.n4 152
R3451 a_15539_n2791.n1 a_15539_n2791.t3 141.923
R3452 a_15539_n2791.n3 a_15539_n2791.n2 10.8376
R3453 a_15539_n2791.n5 a_15539_n2791.n3 2.50485
R3454 a_15705_n2791.t0 a_15705_n2791.n3 370.026
R3455 a_15705_n2791.n0 a_15705_n2791.t5 351.356
R3456 a_15705_n2791.n1 a_15705_n2791.t3 334.717
R3457 a_15705_n2791.n3 a_15705_n2791.t1 325.971
R3458 a_15705_n2791.n1 a_15705_n2791.t4 309.935
R3459 a_15705_n2791.n0 a_15705_n2791.t2 305.683
R3460 a_15705_n2791.n2 a_15705_n2791.n0 16.879
R3461 a_15705_n2791.n3 a_15705_n2791.n2 10.8867
R3462 a_15705_n2791.n2 a_15705_n2791.n1 9.3005
R3463 a_16782_n2425.t0 a_16782_n2425.t1 126.644
R3464 standby.n1 standby.t0 260.322
R3465 standby.n0 standby.t1 194.635
R3466 standby.n1 standby.t2 175.169
R3467 standby.n2 standby.n1 152
R3468 standby.n2 standby.n0 69.674
R3469 standby standby.n2 1.55726
R3470 standby.n0 standby 0.748625
R3471 a_4857_n1521.t0 a_4857_n1521.n1 405.735
R3472 a_4857_n1521.n1 a_4857_n1521.t1 294.611
R3473 a_4857_n1521.n0 a_4857_n1521.t2 254.389
R3474 a_4857_n1521.n0 a_4857_n1521.t3 211.01
R3475 a_4857_n1521.n1 a_4857_n1521.n0 152
R3476 ena_b_33.n5 ena_b_33.t8 402.978
R3477 ena_b_33.n6 ena_b_33.t8 402.978
R3478 ena_b_33.t4 ena_b_33.n2 402.978
R3479 ena_b_33.n3 ena_b_33.t4 402.978
R3480 ena_b_33.t3 ena_b_33.n5 375.649
R3481 ena_b_33.n6 ena_b_33.t3 375.649
R3482 ena_b_33.n4 ena_b_33.t6 375.649
R3483 ena_b_33.n7 ena_b_33.t6 375.649
R3484 ena_b_33.n3 ena_b_33.t7 375.649
R3485 ena_b_33.t7 ena_b_33.n2 375.649
R3486 ena_b_33.n1 ena_b_33.t2 227.887
R3487 ena_b_33.n7 ena_b_33.n2 27.3302
R3488 ena_b_33.n7 ena_b_33.n6 27.3302
R3489 ena_b_33.n4 ena_b_33.n3 27.3302
R3490 ena_b_33.n5 ena_b_33.n4 27.3302
R3491 ena_b_33.n1 ena_b_33.n8 25.0905
R3492 ena_b_33.n1 ena_b_33.t5 12.777
R3493 ena_b_33.n8 ena_b_33.t0 5.5105
R3494 ena_b_33.n8 ena_b_33.t1 5.5105
R3495 ena_b_33.n4 ena_b_33 4.19717
R3496 ena_b_33.n0 ena_b_33.n7 2.93675
R3497 ena_b_33.n1 ena_b_33.n0 1.06508
R3498 ena_b_33.n0 ena_b_33 0.867167
R3499 a_19955_n2791.n1 a_19955_n2791.t4 530.01
R3500 a_19955_n2791.t1 a_19955_n2791.n5 421.021
R3501 a_19955_n2791.n0 a_19955_n2791.t3 337.142
R3502 a_19955_n2791.n3 a_19955_n2791.t0 280.223
R3503 a_19955_n2791.n4 a_19955_n2791.t6 263.173
R3504 a_19955_n2791.n4 a_19955_n2791.t2 227.826
R3505 a_19955_n2791.n0 a_19955_n2791.t5 199.762
R3506 a_19955_n2791.n2 a_19955_n2791.n1 170.81
R3507 a_19955_n2791.n2 a_19955_n2791.n0 167.321
R3508 a_19955_n2791.n5 a_19955_n2791.n4 152
R3509 a_19955_n2791.n1 a_19955_n2791.t7 141.923
R3510 a_19955_n2791.n3 a_19955_n2791.n2 10.8376
R3511 a_19955_n2791.n5 a_19955_n2791.n3 2.50485
R3512 a_20121_n2791.t0 a_20121_n2791.n3 370.026
R3513 a_20121_n2791.n0 a_20121_n2791.t4 351.356
R3514 a_20121_n2791.n1 a_20121_n2791.t3 334.717
R3515 a_20121_n2791.n3 a_20121_n2791.t1 325.971
R3516 a_20121_n2791.n1 a_20121_n2791.t2 309.935
R3517 a_20121_n2791.n0 a_20121_n2791.t5 305.683
R3518 a_20121_n2791.n2 a_20121_n2791.n0 16.879
R3519 a_20121_n2791.n3 a_20121_n2791.n2 10.8867
R3520 a_20121_n2791.n2 a_20121_n2791.n1 9.3005
R3521 a_19567_n2247.t0 a_19567_n2247.n1 386.31
R3522 a_19567_n2247.n1 a_19567_n2247.t1 249.956
R3523 a_19567_n2247.n0 a_19567_n2247.t3 239.04
R3524 a_19567_n2247.n1 a_19567_n2247.n0 175.661
R3525 a_19567_n2247.n0 a_19567_n2247.t2 166.739
R3526 ena.n0 ena.t2 260.322
R3527 ena.n2 ena.t0 194.63
R3528 ena.n0 ena.t1 175.169
R3529 ena.n1 ena.n0 152
R3530 ena.n3 ena.n2 51.6747
R3531 ena ena.n3 4.94983
R3532 ena.n3 ena.n1 3.45996
R3533 ena.n1 ena 1.55726
R3534 ena.n2 ena 0.746125
R3535 a_19003_n2817.n6 a_19003_n2817.n5 746.659
R3536 a_19003_n2817.n0 a_19003_n2817.t5 389.183
R3537 a_19003_n2817.n2 a_19003_n2817.t3 256.988
R3538 a_19003_n2817.n1 a_19003_n2817.n0 251.167
R3539 a_19003_n2817.n1 a_19003_n2817.t1 223.571
R3540 a_19003_n2817.n4 a_19003_n2817.t8 212.081
R3541 a_19003_n2817.n5 a_19003_n2817.n4 181.942
R3542 a_19003_n2817.n0 a_19003_n2817.t4 174.891
R3543 a_19003_n2817.n2 a_19003_n2817.t6 163.803
R3544 a_19003_n2817.n3 a_19003_n2817.t7 139.78
R3545 a_19003_n2817.n3 a_19003_n2817.n2 129.264
R3546 a_19003_n2817.t0 a_19003_n2817.n6 63.3219
R3547 a_19003_n2817.n6 a_19003_n2817.t2 63.3219
R3548 a_19003_n2817.n5 a_19003_n2817.n1 24.6993
R3549 a_19003_n2817.n4 a_19003_n2817.n3 22.6399
R3550 a_19567_n2791.t0 a_19567_n2791.n1 386.31
R3551 a_19567_n2791.n1 a_19567_n2791.t1 249.956
R3552 a_19567_n2791.n0 a_19567_n2791.t3 239.04
R3553 a_19567_n2791.n1 a_19567_n2791.n0 175.661
R3554 a_19567_n2791.n0 a_19567_n2791.t2 166.739
R3555 vg1.t1 vg1.n1 85.228
R3556 vg1.n0 vg1.t3 61.06
R3557 vg1.n2 vg1.t5 54.828
R3558 vg1.n2 vg1.t1 54.828
R3559 vg1.n9 vg1.t0 41.5052
R3560 vg1.n4 vg1.n2 32.951
R3561 vg1.n3 vg1.n1 30.9745
R3562 vg1.n3 vg1.t2 20.9512
R3563 vg1.n10 vg1.n9 3.63479
R3564 vg1.n11 vg1.n1 2.43287
R3565 vg1.n12 vg1.n0 0.471594
R3566 vg1.n9 vg1.n8 0.390524
R3567 vg1.n4 vg1.n3 0.221756
R3568 vg1.n12 vg1.n11 0.146594
R3569 vg1.n11 vg1.n10 0.144647
R3570 vg1 vg1.n12 0.133236
R3571 vg1.n5 vg1.t9 0.0767969
R3572 vg1.n6 vg1.n5 0.0752537
R3573 vg1.n7 vg1.n6 0.0752537
R3574 vg1.n8 vg1.t8 0.0717511
R3575 vg1.n0 vg1 0.0387813
R3576 vg1.n10 vg1.n4 0.0123896
R3577 vg1.n8 vg1.n7 0.00554581
R3578 vg1.n5 vg1.t4 0.00204321
R3579 vg1.n6 vg1.t7 0.00204321
R3580 vg1.n7 vg1.t6 0.00204321
R3581 a_21145_n1869.n0 a_21145_n1869.t0 68.3338
R3582 a_21145_n1869.n0 a_21145_n1869.t1 26.3935
R3583 a_21145_n1869.n1 a_21145_n1869.n0 14.4005
R3584 a_21211_n2817.n4 a_21211_n2817.n0 746.659
R3585 a_21211_n2817.n5 a_21211_n2817.t8 389.183
R3586 a_21211_n2817.n1 a_21211_n2817.t6 256.988
R3587 a_21211_n2817.n6 a_21211_n2817.n5 251.167
R3588 a_21211_n2817.t0 a_21211_n2817.n6 223.571
R3589 a_21211_n2817.n3 a_21211_n2817.t5 212.081
R3590 a_21211_n2817.n4 a_21211_n2817.n3 181.942
R3591 a_21211_n2817.n5 a_21211_n2817.t7 174.891
R3592 a_21211_n2817.n1 a_21211_n2817.t3 163.803
R3593 a_21211_n2817.n2 a_21211_n2817.t4 139.78
R3594 a_21211_n2817.n2 a_21211_n2817.n1 129.264
R3595 a_21211_n2817.n0 a_21211_n2817.t1 63.3219
R3596 a_21211_n2817.n0 a_21211_n2817.t2 63.3219
R3597 a_21211_n2817.n6 a_21211_n2817.n4 24.6993
R3598 a_21211_n2817.n3 a_21211_n2817.n2 22.6399
R3599 xin.n38 xin.t8 594.832
R3600 xin.t18 xin.n5 380.808
R3601 xin.n6 xin.t18 380.808
R3602 xin.n6 xin.t15 380.611
R3603 xin.t15 xin.n5 380.611
R3604 xin.t13 xin.n7 380.611
R3605 xin.n8 xin.t13 380.611
R3606 xin.t19 xin.n4 380.611
R3607 xin.n9 xin.t19 380.611
R3608 xin.n11 xin.t16 380.611
R3609 xin.t16 xin.n10 380.611
R3610 xin.n12 xin.t11 380.611
R3611 xin.t11 xin.n3 380.611
R3612 xin.t10 xin.n13 380.611
R3613 xin.n14 xin.t10 380.611
R3614 xin.t17 xin.n2 380.611
R3615 xin.n15 xin.t17 380.611
R3616 xin.n17 xin.t14 380.611
R3617 xin.t14 xin.n16 380.611
R3618 xin.n18 xin.t12 380.611
R3619 xin.t12 xin.n1 380.611
R3620 xin.t9 xin.n19 380.611
R3621 xin.n20 xin.t9 380.611
R3622 xin.n21 xin.t6 380.611
R3623 xin.t6 xin.n0 380.611
R3624 xin.n38 xin.t21 194.639
R3625 xin.n27 xin.t7 86.3125
R3626 xin.t7 xin.n23 86.3125
R3627 xin.t20 xin.n25 86.3125
R3628 xin.n26 xin.t20 86.3125
R3629 xin.n25 xin.n23 58.6245
R3630 xin.n27 xin.n26 58.6245
R3631 xin.n32 xin.t0 45.927
R3632 xin.n30 xin.n29 20.1298
R3633 xin.n29 xin.n23 12.2455
R3634 xin.n28 xin.n27 11.1505
R3635 xin.n37 xin.n36 4.04311
R3636 xin.n36 xin.n31 3.51336
R3637 xin.n32 xin.n31 3.51061
R3638 xin.n25 xin.n24 3.26098
R3639 xin.n26 xin.n24 2.3255
R3640 xin.n30 xin.n22 1.95915
R3641 xin.n37 xin.n30 1.1106
R3642 xin.n22 xin.n21 0.8105
R3643 xin.n22 xin.n0 0.7905
R3644 xin.n28 xin.n24 0.546796
R3645 xin xin.n38 0.502062
R3646 xin.n38 xin.n37 0.4755
R3647 xin.n29 xin.n28 0.4698
R3648 xin.n8 xin.n5 0.198
R3649 xin.n9 xin.n8 0.198
R3650 xin.n10 xin.n9 0.198
R3651 xin.n10 xin.n3 0.198
R3652 xin.n14 xin.n3 0.198
R3653 xin.n15 xin.n14 0.198
R3654 xin.n16 xin.n15 0.198
R3655 xin.n16 xin.n1 0.198
R3656 xin.n20 xin.n1 0.198
R3657 xin.n21 xin.n20 0.198
R3658 xin.n7 xin.n6 0.198
R3659 xin.n7 xin.n4 0.198
R3660 xin.n11 xin.n4 0.198
R3661 xin.n12 xin.n11 0.198
R3662 xin.n13 xin.n12 0.198
R3663 xin.n13 xin.n2 0.198
R3664 xin.n17 xin.n2 0.198
R3665 xin.n18 xin.n17 0.198
R3666 xin.n19 xin.n18 0.198
R3667 xin.n19 xin.n0 0.198
R3668 xin.t4 xin.t2 0.0760058
R3669 xin.n33 xin.n32 0.0410952
R3670 xin.n34 xin.n31 0.0410952
R3671 xin.n36 xin.n35 0.0410952
R3672 xin.n34 xin.t5 0.0264927
R3673 xin.n33 xin.t1 0.0264885
R3674 xin.n35 xin.t4 0.0264703
R3675 xin.n35 xin.t3 0.0264296
R3676 xin.t3 xin.n34 0.0264114
R3677 xin.t5 xin.n33 0.0264072
R3678 a_19182_n2791.t0 a_19182_n2791.t1 87.1434
R3679 a_2132_n17250.t0 a_2132_n17250.t1 82.3314
R3680 a_24220_n9500.t0 a_24220_n9500.t1 83.56
R3681 a_17913_n2241.t0 a_17913_n2241.n3 370.026
R3682 a_17913_n2241.n0 a_17913_n2241.t3 351.356
R3683 a_17913_n2241.n1 a_17913_n2241.t2 334.717
R3684 a_17913_n2241.n3 a_17913_n2241.t1 325.971
R3685 a_17913_n2241.n1 a_17913_n2241.t4 309.935
R3686 a_17913_n2241.n0 a_17913_n2241.t5 305.683
R3687 a_17913_n2241.n2 a_17913_n2241.n0 16.879
R3688 a_17913_n2241.n3 a_17913_n2241.n2 10.8867
R3689 a_17913_n2241.n2 a_17913_n2241.n1 9.3005
R3690 a_18263_n1869.n3 a_18263_n1869.n2 674.338
R3691 a_18263_n1869.n1 a_18263_n1869.t4 332.58
R3692 a_18263_n1869.n2 a_18263_n1869.n0 284.012
R3693 a_18263_n1869.n2 a_18263_n1869.n1 253.648
R3694 a_18263_n1869.n1 a_18263_n1869.t5 168.701
R3695 a_18263_n1869.n3 a_18263_n1869.t3 96.1553
R3696 a_18263_n1869.t1 a_18263_n1869.n3 65.6672
R3697 a_18263_n1869.n0 a_18263_n1869.t0 65.0005
R3698 a_18263_n1869.n0 a_18263_n1869.t2 45.0005
R3699 a_18359_n1869.t1 a_18359_n1869.t0 198.571
R3700 vg2.n9 vg2.t9 87.8852
R3701 vg2.n2 vg2.t5 87.8852
R3702 vg2.n12 vg2.t6 85.228
R3703 vg2.n5 vg2.t7 85.228
R3704 vg2.n15 vg2.t8 67.0783
R3705 vg2.n11 vg2.t9 54.828
R3706 vg2.t6 vg2.n11 54.828
R3707 vg2.n4 vg2.t5 54.828
R3708 vg2.t7 vg2.n4 54.828
R3709 vg2.n16 vg2.t0 41.0854
R3710 vg2.n11 vg2.n10 30.4005
R3711 vg2.n4 vg2.n3 30.4005
R3712 vg2.n10 vg2.n8 29.1205
R3713 vg2.n12 vg2.n8 29.1205
R3714 vg2.n3 vg2.n1 29.1205
R3715 vg2.n5 vg2.n1 29.1205
R3716 vg2.n13 vg2.n12 2.3255
R3717 vg2.n6 vg2.n5 2.3255
R3718 vg2.n10 vg2.n9 2.13477
R3719 vg2.n3 vg2.n2 2.13477
R3720 vg2.n17 vg2.n16 0.861168
R3721 vg2.n16 vg2.n15 0.714316
R3722 vg2.n8 vg2.n7 0.423227
R3723 vg2.n1 vg2.n0 0.423227
R3724 vg2.n17 vg2.n14 0.371594
R3725 vg2.n18 vg2.n17 0.371594
R3726 vg2.n9 vg2.n7 0.308459
R3727 vg2.n2 vg2.n0 0.308459
R3728 vg2.n13 vg2.n7 0.284875
R3729 vg2.n6 vg2.n0 0.284875
R3730 vg2.n15 vg2.t3 0.170134
R3731 vg2 vg2.n18 0.15675
R3732 vg2.n14 vg2.n13 0.103625
R3733 vg2.n18 vg2.n6 0.103625
R3734 vg2.t1 vg2.t2 0.0652716
R3735 vg2.t4 vg2.t1 0.0652716
R3736 vg2.t3 vg2.t4 0.0652716
R3737 vg2.n14 vg2 0.0505
R3738 vg2.n18 vg2 0.0505
R3739 vrb.n2 vrb.t0 43.1048
R3740 vrb.n0 vrb.t4 22.3777
R3741 vrb.n1 vrb.t1 22.1989
R3742 vrb.n1 vrb.t3 21.3671
R3743 vrb.n0 vrb.t2 21.3663
R3744 vrb.n3 vrb.n2 1.11856
R3745 vrb.n3 vrb.n0 0.759192
R3746 vrb.n2 vrb.n1 0.758408
R3747 vrb vrb.n3 0.0491111
R3748 ena_33.n4 ena_33.t3 398.64
R3749 ena_33.t3 ena_33.n2 398.64
R3750 ena_33.t5 ena_33.n1 398.64
R3751 ena_33.n3 ena_33.t5 398.64
R3752 ena_33.n4 ena_33.t6 371.31
R3753 ena_33.t6 ena_33.n2 371.31
R3754 ena_33.t7 ena_33.n5 371.31
R3755 ena_33.n6 ena_33.t7 371.31
R3756 ena_33.n3 ena_33.t8 371.31
R3757 ena_33.t8 ena_33.n1 371.31
R3758 ena_33.n0 ena_33.t2 227.886
R3759 ena_33.n6 ena_33.n2 27.3302
R3760 ena_33.n5 ena_33.n3 27.3302
R3761 ena_33.n5 ena_33.n4 27.3302
R3762 ena_33.n7 ena_33.n1 25.7735
R3763 ena_33.n0 ena_33.n9 25.0903
R3764 ena_33.n0 ena_33.t4 12.7763
R3765 ena_33.n9 ena_33.t0 5.5105
R3766 ena_33.n9 ena_33.t1 5.5105
R3767 ena_33.n5 ena_33 4.19404
R3768 ena_33.n8 ena_33.n7 2.91956
R3769 ena_33.n7 ena_33.n6 1.55726
R3770 ena_33 ena_33.n8 0.88175
R3771 ena_33.n8 ena_33 0.848417
R3772 ena_33 ena_33.n0 0.794875
R3773 a_18359_n2791.t1 a_18359_n2791.t0 198.571
R3774 a_18525_n2791.t0 a_18525_n2791.t1 60.0005
R3775 a_2130_n20844.t0 a_2130_n20844.t1 82.0028
R3776 a_24530_n21010.t0 a_24530_n21010.t1 81.9478
R3777 a_15083_n2791.t0 a_15083_n2791.t1 60.0005
R3778 a_18932_n15424.t0 a_18932_n15424.t1 83.5579
R3779 a_14285_n2281.n1 a_14285_n2281.n0 953.039
R3780 a_14285_n2281.t0 a_14285_n2281.n1 33.4905
R3781 a_14285_n2281.n1 a_14285_n2281.t3 31.5205
R3782 a_14285_n2281.n0 a_14285_n2281.t2 26.5955
R3783 a_14285_n2281.n0 a_14285_n2281.t1 26.5955
R3784 a_14285_n2079.n0 a_14285_n2079.t1 1201.3
R3785 a_14285_n2079.t0 a_14285_n2079.n0 26.5955
R3786 a_14285_n2079.n0 a_14285_n2079.t2 26.5955
R3787 a_18828_n1869.n3 a_18828_n1869.n2 636.953
R3788 a_18828_n1869.n1 a_18828_n1869.t4 366.856
R3789 a_18828_n1869.n2 a_18828_n1869.n0 300.2
R3790 a_18828_n1869.n2 a_18828_n1869.n1 225.036
R3791 a_18828_n1869.n1 a_18828_n1869.t5 174.056
R3792 a_18828_n1869.n0 a_18828_n1869.t1 70.0005
R3793 a_18828_n1869.n3 a_18828_n1869.t2 68.0124
R3794 a_18828_n1869.t0 a_18828_n1869.n3 63.3219
R3795 a_18828_n1869.n0 a_18828_n1869.t3 61.6672
R3796 a_19182_n1881.t0 a_19182_n1881.t1 87.1434
R3797 a_19003_n1943.n6 a_19003_n1943.n5 746.659
R3798 a_19003_n1943.n0 a_19003_n1943.t8 389.183
R3799 a_19003_n1943.n2 a_19003_n1943.t5 256.988
R3800 a_19003_n1943.n1 a_19003_n1943.n0 251.167
R3801 a_19003_n1943.n1 a_19003_n1943.t1 223.571
R3802 a_19003_n1943.n4 a_19003_n1943.t7 212.081
R3803 a_19003_n1943.n5 a_19003_n1943.n4 181.942
R3804 a_19003_n1943.n0 a_19003_n1943.t3 174.891
R3805 a_19003_n1943.n2 a_19003_n1943.t6 163.803
R3806 a_19003_n1943.n3 a_19003_n1943.t4 139.78
R3807 a_19003_n1943.n3 a_19003_n1943.n2 129.264
R3808 a_19003_n1943.t0 a_19003_n1943.n6 63.3219
R3809 a_19003_n1943.n6 a_19003_n1943.t2 63.3219
R3810 a_19003_n1943.n5 a_19003_n1943.n1 24.6993
R3811 a_19003_n1943.n4 a_19003_n1943.n3 22.6399
R3812 vn.n0 vn.t9 59.0048
R3813 vn.n3 vn.t5 125.335
R3814 vn.n3 vn.n6 96.4272
R3815 vn.n4 vn.n2 96.4272
R3816 vn.n1 vn.n0 0.750908
R3817 vn.n3 vn.t3 85.228
R3818 vn.t3 vn.n2 85.228
R3819 vn.n4 vn.t8 85.228
R3820 vn.n6 vn.t8 85.228
R3821 vn vn.t1 60.9515
R3822 vn vn.n5 53.6683
R3823 vn.n2 vn 2.35462
R3824 vn vn.t7 22.0141
R3825 vn vn.n3 2.50212
R3826 vn vn.n7 16.8187
R3827 vn.n5 vn.t2 6.92425
R3828 vn.n5 vn.t0 6.92425
R3829 vn.n7 vn.t4 4.3505
R3830 vn.n7 vn.t6 4.3505
R3831 vn.t5 vn 87.6035
R3832 vn.n1 vn 2.77387
R3833 vn.n6 vn.n0 1.55632
R3834 vn.n1 vn.n4 2.20282
R3835 a_10620_n7674.t0 a_10620_n7674.t1 82.5973
R3836 a_24220_n7840.t0 a_24220_n7840.t1 83.56
R3837 x7.x2.x3.CLK.n3 x7.x2.x3.CLK.t0 372.361
R3838 x7.x2.x3.CLK.n2 x7.x2.x3.CLK.t5 333.651
R3839 x7.x2.x3.CLK.n2 x7.x2.x3.CLK.t2 297.233
R3840 x7.x2.x3.CLK.n1 x7.x2.x3.CLK.t3 294.557
R3841 x7.x2.x3.CLK.n4 x7.x2.x3.CLK.t1 231.921
R3842 x7.x2.x3.CLK.n1 x7.x2.x3.CLK.t4 211.01
R3843 x7.x2.x3.CLK x7.x2.x3.CLK.n2 195.701
R3844 x7.x2.x3.CLK.n0 x7.x2.x3.CLK.n1 152
R3845 x7.x2.x3.CLK.n4 x7.x2.x3.CLK.n0 40.9605
R3846 x7.x2.x3.CLK.n3 x7.x2.x3.CLK 25.2739
R3847 x7.x2.x3.CLK.n4 x7.x2.x3.CLK.n3 18.1966
R3848 x7.x2.x3.CLK.n0 x7.x2.x3.CLK 10.4234
R3849 x7.x2.x3.CLK x7.x2.x3.CLK.n4 2.5605
R3850 x7.x2.x3.CLK.n0 x7.x2.x3.CLK 2.01193
R3851 a_15960_n2791.n1 a_15960_n2791.n0 926.024
R3852 a_15960_n2791.t0 a_15960_n2791.n1 82.0838
R3853 a_15960_n2791.n0 a_15960_n2791.t1 63.3338
R3854 a_15960_n2791.n1 a_15960_n2791.t2 63.3219
R3855 a_15960_n2791.n0 a_15960_n2791.t3 29.7268
R3856 a_2130_n19516.t0 a_2130_n19516.t1 82.0028
R3857 a_24530_n19682.t0 a_24530_n19682.t1 81.9478
R3858 a_20579_n2247.n0 a_20579_n2247.t2 1327.82
R3859 a_20579_n2247.n0 a_20579_n2247.t1 194.655
R3860 a_20579_n2247.t0 a_20579_n2247.n0 63.3219
R3861 a_15083_n1881.t0 a_15083_n1881.t1 60.0005
R3862 a_18481_n2273.n3 a_18481_n2273.n2 647.119
R3863 a_18481_n2273.n1 a_18481_n2273.t4 350.253
R3864 a_18481_n2273.n2 a_18481_n2273.n0 260.339
R3865 a_18481_n2273.n2 a_18481_n2273.n1 246.119
R3866 a_18481_n2273.n1 a_18481_n2273.t5 189.588
R3867 a_18481_n2273.n3 a_18481_n2273.t3 89.1195
R3868 a_18481_n2273.n0 a_18481_n2273.t0 63.3338
R3869 a_18481_n2273.t1 a_18481_n2273.n3 41.0422
R3870 a_18481_n2273.n0 a_18481_n2273.t2 31.9797
R3871 a_18525_n1881.t0 a_18525_n1881.t1 60.0005
R3872 x7.x2.x4.CLK.n3 x7.x2.x4.CLK.t0 372.361
R3873 x7.x2.x4.CLK.n2 x7.x2.x4.CLK.t5 333.651
R3874 x7.x2.x4.CLK.n2 x7.x2.x4.CLK.t2 297.233
R3875 x7.x2.x4.CLK.n1 x7.x2.x4.CLK.t3 294.557
R3876 x7.x2.x4.CLK.n4 x7.x2.x4.CLK.t1 231.921
R3877 x7.x2.x4.CLK.n1 x7.x2.x4.CLK.t4 211.01
R3878 x7.x2.x4.CLK x7.x2.x4.CLK.n2 195.701
R3879 x7.x2.x4.CLK.n0 x7.x2.x4.CLK.n1 152
R3880 x7.x2.x4.CLK.n4 x7.x2.x4.CLK.n0 40.9605
R3881 x7.x2.x4.CLK.n3 x7.x2.x4.CLK 25.2781
R3882 x7.x2.x4.CLK.n4 x7.x2.x4.CLK.n3 18.1966
R3883 x7.x2.x4.CLK.n0 x7.x2.x4.CLK 10.4234
R3884 x7.x2.x4.CLK x7.x2.x4.CLK.n4 2.5605
R3885 x7.x2.x4.CLK.n0 x7.x2.x4.CLK 2.01193
R3886 a_18168_n2791.n1 a_18168_n2791.n0 926.024
R3887 a_18168_n2791.t0 a_18168_n2791.n1 82.0838
R3888 a_18168_n2791.n0 a_18168_n2791.t3 63.3338
R3889 a_18168_n2791.n1 a_18168_n2791.t1 63.3219
R3890 a_18168_n2791.n0 a_18168_n2791.t2 29.7268
R3891 a_16055_n2791.n3 a_16055_n2791.n2 674.338
R3892 a_16055_n2791.n1 a_16055_n2791.t4 332.58
R3893 a_16055_n2791.n2 a_16055_n2791.n0 284.012
R3894 a_16055_n2791.n2 a_16055_n2791.n1 253.648
R3895 a_16055_n2791.n1 a_16055_n2791.t5 168.701
R3896 a_16055_n2791.n3 a_16055_n2791.t3 96.1553
R3897 a_16055_n2791.t0 a_16055_n2791.n3 65.6672
R3898 a_16055_n2791.n0 a_16055_n2791.t2 65.0005
R3899 a_16055_n2791.n0 a_16055_n2791.t1 45.0005
R3900 x7.x1.x4.Q x7.x1.x4.Q.t0 240.05
R3901 x7.x1.x4.Q x7.x1.x4.Q.t1 155.386
R3902 a_14009_n2404.t0 a_14009_n2404.n3 669.389
R3903 a_14009_n2404.n0 a_14009_n2404.t1 326.493
R3904 a_14009_n2404.n0 a_14009_n2404.t2 249.615
R3905 a_14009_n2404.n1 a_14009_n2404.t3 249.615
R3906 a_14009_n2404.n2 a_14009_n2404.t4 241.536
R3907 a_14009_n2404.n2 a_14009_n2404.t5 169.237
R3908 a_14009_n2404.n3 a_14009_n2404.n2 152
R3909 a_14009_n2404.n3 a_14009_n2404.n1 108.529
R3910 a_14009_n2404.n1 a_14009_n2404.n0 26.6245
R3911 a_24530_n20678.t0 a_24530_n20678.t1 81.9478
R3912 a_15539_n2241.n1 a_15539_n2241.t5 530.01
R3913 a_15539_n2241.t0 a_15539_n2241.n5 421.021
R3914 a_15539_n2241.n0 a_15539_n2241.t3 337.142
R3915 a_15539_n2241.n3 a_15539_n2241.t1 280.223
R3916 a_15539_n2241.n4 a_15539_n2241.t4 263.173
R3917 a_15539_n2241.n4 a_15539_n2241.t6 227.826
R3918 a_15539_n2241.n0 a_15539_n2241.t2 199.762
R3919 a_15539_n2241.n2 a_15539_n2241.n1 170.81
R3920 a_15539_n2241.n2 a_15539_n2241.n0 167.321
R3921 a_15539_n2241.n5 a_15539_n2241.n4 152
R3922 a_15539_n2241.n1 a_15539_n2241.t7 141.923
R3923 a_15539_n2241.n3 a_15539_n2241.n2 10.8376
R3924 a_15539_n2241.n5 a_15539_n2241.n3 2.50485
R3925 a_16729_n1869.n0 a_16729_n1869.t1 68.3338
R3926 a_16729_n1869.n0 a_16729_n1869.t0 26.3935
R3927 a_16729_n1869.n1 a_16729_n1869.n0 14.4005
R3928 a_16055_n1869.n3 a_16055_n1869.n2 674.338
R3929 a_16055_n1869.n1 a_16055_n1869.t4 332.58
R3930 a_16055_n1869.n2 a_16055_n1869.n0 284.012
R3931 a_16055_n1869.n2 a_16055_n1869.n1 253.648
R3932 a_16055_n1869.n1 a_16055_n1869.t5 168.701
R3933 a_16055_n1869.t0 a_16055_n1869.n3 96.1553
R3934 a_16055_n1869.n3 a_16055_n1869.t2 65.6672
R3935 a_16055_n1869.n0 a_16055_n1869.t1 65.0005
R3936 a_16055_n1869.n0 a_16055_n1869.t3 45.0005
R3937 a_2132_n15258.t0 a_2132_n15258.t1 83.9223
R3938 a_18990_n2425.t0 a_18990_n2425.t1 126.644
R3939 a_24530_n19350.t0 a_24530_n19350.t1 81.9478
R3940 a_16163_n2247.n0 a_16163_n2247.t2 1327.82
R3941 a_16163_n2247.t0 a_16163_n2247.n0 194.655
R3942 a_16163_n2247.n0 a_16163_n2247.t1 63.3219
R3943 a_2132_n16918.t0 a_2132_n16918.t1 82.3314
R3944 a_18932_n17084.t0 a_18932_n17084.t1 83.5579
R3945 a_10620_n9334.t0 a_10620_n9334.t1 83.9243
R3946 a_3134_n13324.t0 a_3134_n13324.t1 83.9223
R3947 x7.x1.x2.Q x7.x1.x2.Q.t0 240.05
R3948 x7.x1.x2.Q x7.x1.x2.Q.t1 155.386
R3949 a_18932_n17748.t0 a_18932_n17748.t1 83.5579
R3950 a_18937_n2791.t0 a_18937_n2791.t1 94.7268
R3951 a_17359_n2247.t0 a_17359_n2247.n1 386.31
R3952 a_17359_n2247.n1 a_17359_n2247.t1 249.956
R3953 a_17359_n2247.n0 a_17359_n2247.t2 239.04
R3954 a_17359_n2247.n1 a_17359_n2247.n0 175.661
R3955 a_17359_n2247.n0 a_17359_n2247.t3 166.739
R3956 a_24530_n22338.t0 a_24530_n22338.t1 81.9492
R3957 dout_filt.n1 dout_filt.t0 687.288
R3958 dout_filt dout_filt.t2 229.845
R3959 dout_filt.n2 dout_filt.t1 223.571
R3960 dout_filt.n2 dout_filt.n1 139.672
R3961 dout_filt.n0 dout_filt.t4 97.4114
R3962 dout_filt.n0 dout_filt.t3 56.9639
R3963 dout_filt dout_filt.n2 4.70638
R3964 dout_filt dout_filt.n1 4.70638
R3965 dout_filt dout_filt.n0 2.24782
R3966 x4.out_b.n0 x4.out_b.t0 227.887
R3967 x4.out_b.n0 x4.out_b.n1 25.0905
R3968 x4.out_b.n0 x4.out_b.t3 12.777
R3969 x4.out_b.n1 x4.out_b.t1 5.5105
R3970 x4.out_b.n1 x4.out_b.t2 5.5105
R3971 x4.out_b x4.out_b.n0 0.83175
R3972 a_15960_n1881.n1 a_15960_n1881.n0 926.024
R3973 a_15960_n1881.n0 a_15960_n1881.t2 82.0838
R3974 a_15960_n1881.n1 a_15960_n1881.t0 63.3338
R3975 a_15960_n1881.n0 a_15960_n1881.t3 63.3219
R3976 a_15960_n1881.t1 a_15960_n1881.n1 29.7268
R3977 a_20471_n2791.n3 a_20471_n2791.n2 674.338
R3978 a_20471_n2791.n1 a_20471_n2791.t5 332.58
R3979 a_20471_n2791.n2 a_20471_n2791.n0 284.012
R3980 a_20471_n2791.n2 a_20471_n2791.n1 253.648
R3981 a_20471_n2791.n1 a_20471_n2791.t4 168.701
R3982 a_20471_n2791.n3 a_20471_n2791.t2 96.1553
R3983 a_20471_n2791.t0 a_20471_n2791.n3 65.6672
R3984 a_20471_n2791.n0 a_20471_n2791.t3 65.0005
R3985 a_20471_n2791.n0 a_20471_n2791.t1 45.0005
R3986 a_24220_n9168.t0 a_24220_n9168.t1 83.56
R3987 a_21036_n2791.n3 a_21036_n2791.n2 636.953
R3988 a_21036_n2791.n1 a_21036_n2791.t5 366.856
R3989 a_21036_n2791.n2 a_21036_n2791.n0 300.2
R3990 a_21036_n2791.n2 a_21036_n2791.n1 225.036
R3991 a_21036_n2791.n1 a_21036_n2791.t4 174.056
R3992 a_21036_n2791.n0 a_21036_n2791.t0 70.0005
R3993 a_21036_n2791.n3 a_21036_n2791.t2 68.0124
R3994 a_21036_n2791.t1 a_21036_n2791.n3 63.3219
R3995 a_21036_n2791.n0 a_21036_n2791.t3 61.6672
R3996 a_18937_n1869.n0 a_18937_n1869.t1 68.3338
R3997 a_18937_n1869.n0 a_18937_n1869.t0 26.3935
R3998 a_18937_n1869.n1 a_18937_n1869.n0 14.4005
R3999 a_17747_n2791.n1 a_17747_n2791.t7 530.01
R4000 a_17747_n2791.t0 a_17747_n2791.n5 421.021
R4001 a_17747_n2791.n0 a_17747_n2791.t6 337.142
R4002 a_17747_n2791.n3 a_17747_n2791.t1 280.223
R4003 a_17747_n2791.n4 a_17747_n2791.t3 263.173
R4004 a_17747_n2791.n4 a_17747_n2791.t5 227.826
R4005 a_17747_n2791.n0 a_17747_n2791.t2 199.762
R4006 a_17747_n2791.n2 a_17747_n2791.n1 170.81
R4007 a_17747_n2791.n2 a_17747_n2791.n0 167.321
R4008 a_17747_n2791.n5 a_17747_n2791.n4 152
R4009 a_17747_n2791.n1 a_17747_n2791.t4 141.923
R4010 a_17747_n2791.n3 a_17747_n2791.n2 10.8376
R4011 a_17747_n2791.n5 a_17747_n2791.n3 2.50485
R4012 a_17359_n2791.t0 a_17359_n2791.n1 386.31
R4013 a_17359_n2791.n1 a_17359_n2791.t1 249.956
R4014 a_17359_n2791.n0 a_17359_n2791.t3 239.04
R4015 a_17359_n2791.n1 a_17359_n2791.n0 175.661
R4016 a_17359_n2791.n0 a_17359_n2791.t2 166.739
R4017 a_2130_n20512.t0 a_2130_n20512.t1 82.0028
R4018 a_18263_n2791.n3 a_18263_n2791.n2 674.338
R4019 a_18263_n2791.n1 a_18263_n2791.t4 332.58
R4020 a_18263_n2791.n2 a_18263_n2791.n0 284.012
R4021 a_18263_n2791.n2 a_18263_n2791.n1 253.648
R4022 a_18263_n2791.n1 a_18263_n2791.t5 168.701
R4023 a_18263_n2791.n3 a_18263_n2791.t3 96.1553
R4024 a_18263_n2791.t0 a_18263_n2791.n3 65.6672
R4025 a_18263_n2791.n0 a_18263_n2791.t2 65.0005
R4026 a_18263_n2791.n0 a_18263_n2791.t1 45.0005
R4027 a_2132_n14926.t0 a_2132_n14926.t1 83.9223
R4028 a_18932_n15092.t0 a_18932_n15092.t1 83.5579
R4029 a_14357_n2743.t0 a_14357_n2743.t1 64.6411
R4030 dout.n0 dout.t1 120.561
R4031 dout.n0 dout.t0 61.4115
R4032 dout dout.n0 3.88384
R4033 a_20376_n1881.n1 a_20376_n1881.n0 926.024
R4034 a_20376_n1881.t1 a_20376_n1881.n1 82.0838
R4035 a_20376_n1881.n0 a_20376_n1881.t0 63.3338
R4036 a_20376_n1881.n1 a_20376_n1881.t2 63.3219
R4037 a_20376_n1881.n0 a_20376_n1881.t3 29.7268
R4038 a_20471_n1869.n3 a_20471_n1869.n2 674.338
R4039 a_20471_n1869.n1 a_20471_n1869.t5 332.58
R4040 a_20471_n1869.n2 a_20471_n1869.n0 284.012
R4041 a_20471_n1869.n2 a_20471_n1869.n1 253.648
R4042 a_20471_n1869.n1 a_20471_n1869.t4 168.701
R4043 a_20471_n1869.t1 a_20471_n1869.n3 96.1553
R4044 a_20471_n1869.n3 a_20471_n1869.t2 65.6672
R4045 a_20471_n1869.n0 a_20471_n1869.t0 65.0005
R4046 a_20471_n1869.n0 a_20471_n1869.t3 45.0005
R4047 x7.x1.x3.CLK.n3 x7.x1.x3.CLK.t0 372.361
R4048 x7.x1.x3.CLK.n2 x7.x1.x3.CLK.t4 333.651
R4049 x7.x1.x3.CLK.n2 x7.x1.x3.CLK.t5 297.233
R4050 x7.x1.x3.CLK.n0 x7.x1.x3.CLK.t2 294.557
R4051 x7.x1.x3.CLK.n4 x7.x1.x3.CLK.t1 231.921
R4052 x7.x1.x3.CLK.n0 x7.x1.x3.CLK.t3 211.01
R4053 x7.x1.x3.CLK x7.x1.x3.CLK.n2 195.701
R4054 x7.x1.x3.CLK.n1 x7.x1.x3.CLK.n0 152
R4055 x7.x1.x3.CLK.n4 x7.x1.x3.CLK.n1 41.5091
R4056 x7.x1.x3.CLK.n3 x7.x1.x3.CLK 25.2739
R4057 x7.x1.x3.CLK.n4 x7.x1.x3.CLK.n3 18.1966
R4058 x7.x1.x3.CLK.n1 x7.x1.x3.CLK 4.20621
R4059 x7.x1.x3.CLK x7.x1.x3.CLK.n4 2.5605
R4060 x7.x2.x2.Q x7.x2.x2.Q.t0 246.839
R4061 x7.x2.x2.Q x7.x2.x2.Q.t1 148.597
R4062 a_14035_n2743.t0 a_14035_n2743.t1 60.0005
R4063 a_24530_n20346.t0 a_24530_n20346.t1 81.9478
R4064 a_18932_n14760.t0 a_18932_n14760.t1 83.5579
R4065 x7.x1.x3.Q x7.x1.x3.Q.t0 240.05
R4066 x7.x1.x3.Q x7.x1.x3.Q.t1 155.386
R4067 a_2130_n19184.t0 a_2130_n19184.t1 82.0028
R4068 a_24530_n19018.t0 a_24530_n19018.t1 81.9478
R4069 a_10620_n9002.t0 a_10620_n9002.t1 83.9243
R4070 a_14035_n2281.t0 a_14035_n2281.t1 60.9236
R4071 a_24220_n8836.t0 a_24220_n8836.t1 83.56
R4072 a_2130_n20180.t0 a_2130_n20180.t1 82.0028
R4073 a_2130_n22172.t0 a_2130_n22172.t1 82.0028
R4074 a_24530_n22006.t0 a_24530_n22006.t1 81.9492
R4075 a_2130_n21840.t0 a_2130_n21840.t1 82.0028
R4076 a_2132_n16586.t0 a_2132_n16586.t1 83.9223
R4077 a_18932_n16420.t0 a_18932_n16420.t1 83.5579
R4078 a_10620_n8670.t0 a_10620_n8670.t1 83.9243
R4079 a_22601_n15524.t0 a_22601_n15524.t1 120.212
R4080 a_20579_n2425.n0 a_20579_n2425.t2 1327.82
R4081 a_20579_n2425.n0 a_20579_n2425.t1 194.655
R4082 a_20579_n2425.t0 a_20579_n2425.n0 63.3219
R4083 a_21198_n2247.t0 a_21198_n2247.t1 126.644
R4084 a_17747_n2241.n1 a_17747_n2241.t4 530.01
R4085 a_17747_n2241.t0 a_17747_n2241.n5 421.021
R4086 a_17747_n2241.n0 a_17747_n2241.t2 337.142
R4087 a_17747_n2241.n3 a_17747_n2241.t1 280.223
R4088 a_17747_n2241.n4 a_17747_n2241.t3 263.173
R4089 a_17747_n2241.n4 a_17747_n2241.t6 227.826
R4090 a_17747_n2241.n0 a_17747_n2241.t5 199.762
R4091 a_17747_n2241.n2 a_17747_n2241.n1 170.81
R4092 a_17747_n2241.n2 a_17747_n2241.n0 167.321
R4093 a_17747_n2241.n5 a_17747_n2241.n4 152
R4094 a_17747_n2241.n1 a_17747_n2241.t7 141.923
R4095 a_17747_n2241.n3 a_17747_n2241.n2 10.8376
R4096 a_17747_n2241.n5 a_17747_n2241.n3 2.50485
R4097 a_2132_n14594.t0 a_2132_n14594.t1 82.3314
R4098 a_18932_n14428.t0 a_18932_n14428.t1 83.5579
R4099 a_16163_n2425.n0 a_16163_n2425.t2 1327.82
R4100 a_16163_n2425.t0 a_16163_n2425.n0 194.655
R4101 a_16163_n2425.n0 a_16163_n2425.t1 63.3219
R4102 a_18371_n2247.n0 a_18371_n2247.t1 1327.82
R4103 a_18371_n2247.n0 a_18371_n2247.t2 194.655
R4104 a_18371_n2247.t0 a_18371_n2247.n0 63.3219
R4105 a_24220_n8504.t0 a_24220_n8504.t1 83.56
R4106 x7.x2.x4.Q x7.x2.x4.Q.t0 246.839
R4107 x7.x2.x4.Q x7.x2.x4.Q.t1 148.597
R4108 a_18932_n16752.t0 a_18932_n16752.t1 83.5579
R4109 a_2130_n21508.t0 a_2130_n21508.t1 82.0028
R4110 a_24530_n21674.t0 a_24530_n21674.t1 81.9478
R4111 a_21390_n2791.t0 a_21390_n2791.t1 87.1434
R4112 a_2130_n18852.t0 a_2130_n18852.t1 82.0028
R4113 a_21390_n1881.t0 a_21390_n1881.t1 87.1434
R4114 a_8268_n12482.t0 a_8268_n12482.t1 199.762
R4115 a_21145_n2791.t0 a_21145_n2791.t1 94.7268
R4116 a_16782_n2247.t0 a_16782_n2247.t1 126.644
R4117 x7.x2.x3.Q x7.x2.x3.Q.t0 246.839
R4118 x7.x2.x3.Q x7.x2.x3.Q.t1 148.597
R4119 a_10620_n8006.t0 a_10620_n8006.t1 83.9243
R4120 a_2132_n16254.t0 a_2132_n16254.t1 83.9053
R4121 a_16729_n2791.t0 a_16729_n2791.t1 94.7268
R4122 a_2132_n17914.t0 a_2132_n17914.t1 83.9223
R4123 a_21198_n2425.t0 a_21198_n2425.t1 126.644
R4124 a_18932_n16088.t0 a_18932_n16088.t1 83.5579
R4125 a_18371_n2425.n0 a_18371_n2425.t2 1327.82
R4126 a_18371_n2425.n0 a_18371_n2425.t1 194.655
R4127 a_18371_n2425.t0 a_18371_n2425.n0 63.3219
R4128 a_18990_n2247.t0 a_18990_n2247.t1 126.644
R4129 a_2132_n14262.t0 a_2132_n14262.t1 83.9053
R4130 a_2132_n15922.t0 a_2132_n15922.t1 83.9223
C0 dvdd x7.x2.x4.CLK 1.2179f
C1 x7.x1.x4.CLK dvss_ip 0.069883f
C2 dvss_ip dout_ip 6.7836f
C3 dvdd x7.x3.B2 6.00136f
C4 ena_ip x7.x1.x2.CLK 0.073063f
C5 vg1 xout 0.637153f
C6 x4.in_b standby_ip 1.51792f
C7 ena_ip x7.x1.x3.CLK 0.347396f
C8 vg1 vg2 1.37396f
C9 ena_ip x7.x1.x2.Q 0.035311f
C10 vn dout_ip 0.038056f
C11 dvss_ip vg1 6.71865f
C12 x7.x5.TE_B dout_filt 0.716005f
C13 dvdd x7.x1.x2.CLK 0.406962f
C14 standby_33 x4.in_b 1.05054f
C15 avdd standby_ip 0.688025f
C16 x7.x2.x3.CLK x7.x2.x2.Q 0.040893f
C17 dvdd x7.x1.x3.CLK 1.22948f
C18 x7.x2.x3.Q x4.in_b 0.035311f
C19 ibias standby_ip 0.288754f
C20 dvdd x7.x1.x2.Q 0.116301f
C21 x4.in_b dout_ip 0.326219f
C22 avdd standby_33 8.99931f
C23 inv_m1 inv_m2 0.947856f
C24 ena_ip standby_ip 4.64341f
C25 inv_in tail 0.57662f
C26 dvss_ip dout_filt 7.44028f
C27 ibias standby_33 1.11373f
C28 x7.x2.x3.CLK x7.x3.A2 0.111333f
C29 inv_in standby_33 0.08455f
C30 dvdd standby_ip 10.3838f
C31 avdd_ip vg1 1.83228f
C32 x7.x1.x4.CLK ena_ip 0.347451f
C33 ena_ip dout_ip 0.203453f
C34 inv_in dout_ip 0.074891f
C35 x7.x2.x4.Q x7.x3.A2 0.061065f
C36 dvdd standby_33 0.092517f
C37 avdd ena 0.026836f
C38 avss standby_ip 1.86785f
C39 x4.in_b dout_filt 0.02156f
C40 x7.x1.x4.CLK dvdd 1.22125f
C41 ena_33 ena_b_33 1.23205f
C42 dvdd x7.x2.x3.Q 0.112734f
C43 x7.x3.B2 x7.x1.x2.CLK 0.044383f
C44 dvdd dout_ip 1.37976f
C45 ena_ip ena 0.081602f
C46 x4.out_b ena_b_33 0.019576f
C47 x7.x1.x3.CLK x7.x3.B2 0.095485f
C48 x7.x1.x2.Q x7.x3.B2 0.012057f
C49 avss standby_33 1.55838f
C50 x7.x5.TE_B x7.x2.x2.CLK 0.012819f
C51 dvdd ena 0.377442f
C52 inv_in dout_filt 0.016514f
C53 inv_m1 dout_ip 0.086642f
C54 x7.x3.B2 standby_ip 0.121072f
C55 x7.x5.TE_B x7.x3.A2 0.724301f
C56 x7.x1.x3.CLK x7.x1.x2.Q 0.040893f
C57 dvdd dout_filt 1.76157f
C58 ena_ip standby 0.035742f
C59 x7.x2.x4.CLK x7.x2.x3.Q 0.040893f
C60 x7.x1.x4.CLK x7.x2.x4.CLK 0.0262f
C61 x7.x1.x4.CLK x7.x3.B2 0.095442f
C62 dvss_ip x7.x3.A2 1.50207f
C63 x7.x3.B2 dout_ip 0.187422f
C64 x7.x2.x2.CLK x4.in_b 0.073414f
C65 dvdd standby 0.386478f
C66 x7.x2.x2.Q x4.in_b 0.035311f
C67 inv_m2 dout_ip 0.58911f
C68 dvss_ip dout 6.66227f
C69 avdd ena_33 9.25241f
C70 x7.x3.A2 x4.in_b 0.752988f
C71 avdd x4.out_b 7.47211f
C72 xin xout 12.4713f
C73 dvdd x7.x2.x2.CLK 0.367738f
C74 dvdd x7.x2.x2.Q 0.11753f
C75 vg1 vrb 0.41458f
C76 xin vg2 6.28706f
C77 standby_ip dout_ip 0.055907f
C78 dvss_ip xin 1.63134f
C79 ena_ip x7.x1.x3.Q 0.035311f
C80 x7.x2.x3.CLK x4.in_b 0.347492f
C81 vn xin 2.31407f
C82 dvdd x7.x3.A2 5.3536f
C83 ena_33 avss 5.31495f
C84 dvdd x7.x1.x3.Q 0.112744f
C85 dvdd x7.x1.x4.Q 0.117621f
C86 vbp dvss_ip 1.29294f
C87 x4.out_b avss 1.60459f
C88 dvdd dout 0.550876f
C89 xout vg2 0.938912f
C90 dvss_ip xout 14.1458f
C91 avdd_ip xin 6.15688f
C92 dvss_ip vg2 3.94057f
C93 dvdd x7.x2.x3.CLK 1.15446f
C94 avdd_ip ena_b_33 2.29698f
C95 vn xout 0.040555f
C96 standby standby_ip 0.045124f
C97 dout_ip dout_filt 3.64627f
C98 avdd ena_b_33 11.963599f
C99 inv_in xin 0.323721f
C100 dvdd x7.x2.x4.Q 0.117611f
C101 vn dvss_ip 6.67609f
C102 x7.x2.x4.CLK x7.x3.A2 0.099468f
C103 x7.x2.x2.CLK x7.x1.x2.CLK 0.011009f
C104 x7.x5.TE_B x4.in_b 0.01498f
C105 x7.x3.A2 x7.x3.B2 1.61077f
C106 x7.x1.x3.Q x7.x3.B2 0.012117f
C107 ena_ip ena_b_33 0.931668f
C108 x7.x1.x4.Q x7.x3.B2 0.061065f
C109 avdd_ip xout 6.8108f
C110 vg2 icnode 0.421477f
C111 dvss_ip x4.in_b 3.69012f
C112 inv_in vbp 0.307286f
C113 avdd_ip vg2 0.280688f
C114 dvss_ip avdd_ip 20.4556f
C115 standby ena 0.095384f
C116 inv_in xout 1.30855f
C117 dvss_ip ibias 0.014158f
C118 ena_b_33 avss 1.7988f
C119 inv_in vg2 0.137694f
C120 ena_ip dvss_ip 0.012218f
C121 dvdd x7.x5.TE_B 0.382951f
C122 inv_in dvss_ip 15.0668f
C123 x4.out_b standby_ip 0.931668f
C124 inv_in vn 0.109718f
C125 avdd_ip icnode 43.4983f
C126 dvdd dvss_ip 20.229f
C127 x7.x2.x3.CLK x7.x1.x3.CLK 0.0262f
C128 x4.out_b standby_33 0.696369f
C129 avdd x4.in_b 0.805158f
C130 avdd icnode 0.341154f
C131 ibias x4.in_b 0.300759f
C132 avdd avdd_ip 9.31081f
C133 x7.x3.A2 x7.x2.x3.Q 0.012117f
C134 ena_ip x4.in_b 3.80832f
C135 x7.x1.x4.CLK x7.x1.x3.Q 0.040893f
C136 x7.x3.A2 dout_ip 0.251518f
C137 inv_in icnode 0.110238f
C138 inv_in avdd_ip 0.669037f
C139 inv_m1 dvss_ip 3.10116f
C140 ena_ip avdd 0.709432f
C141 avdd inv_in 0.024554f
C142 dvdd x4.in_b 6.03413f
C143 ena_ip ibias 0.172379f
C144 dvdd avdd 0.136618f
C145 dvss_ip x7.x2.x4.CLK 0.073361f
C146 avss x4.in_b 1.88593f
C147 avss icnode 0.021172f
C148 dvss_ip x7.x3.B2 1.48709f
C149 dvdd ibias 0.083154f
C150 tail xin 1.67389f
C151 avdd_ip avss 0.575284f
C152 x7.x3.A2 dout_filt 0.193457f
C153 dvdd ena_ip 7.75581f
C154 dvdd inv_in 0.696511f
C155 avdd avss 0.108894p
C156 inv_m2 dvss_ip 1.69984f
C157 ena_ip avss 1.87875f
C158 dout dout_filt 0.639323f
C159 inv_in avss 0.144174f
C160 tail vbp 9.31212f
C161 x7.x2.x4.CLK x4.in_b 0.347451f
C162 vrb vg2 4.64004f
C163 x4.in_b x7.x3.B2 0.017099f
C164 inv_in inv_m1 0.243271f
C165 dvss_ip vrb 1.19104f
C166 dvdd avss 0.230646f
C167 vg1 xin 0.215332p
C168 tail xout 1.22898f
C169 tail dvss_ip 0.410396f
C170 x7.x5.TE_B dout_ip 0.153671f
C171 ena_ip x7.x3.B2 0.701454f
C172 dvss_ip standby_33 3.43223f
C173 tail vn 0.561519f
C174 x7.x2.x2.CLK x7.x3.A2 0.055466f
C175 x7.x2.x2.Q x7.x3.A2 0.012057f
C176 xout dvss 31.328293f
C177 xin dvss 85.24696f
C178 dout dvss 4.99223f
C179 standby dvss 1.31811f
C180 ena dvss 1.29717f
C181 avss dvss 16.730371f
C182 ibias dvss 5.70727f
C183 dvdd dvss 0.137133p
C184 avdd dvss 96.62521f
C185 vg1 dvss 19.553183f
C186 vrb dvss 7.274848f
C187 icnode dvss 37.841305f
C188 vg2 dvss 0.160023p
C189 tail dvss 0.488561f
C190 inv_m2 dvss 0.561945f
C191 inv_m1 dvss -0.317498f
C192 inv_in dvss 8.245181f
C193 vn dvss 5.99695f
C194 vbp dvss 18.663542f
C195 x4.out_b dvss 1.060882f
C196 ena_b_33 dvss 1.758028f
C197 ena_33 dvss 4.924316f
C198 x7.x2.x4.Q dvss 0.100179f
C199 x7.x2.x3.Q dvss 0.092032f
C200 x7.x2.x4.CLK dvss 0.510343f
C201 x7.x2.x2.Q dvss 0.092454f
C202 dout_filt dvss 13.912813f
C203 x7.x2.x3.CLK dvss 0.539804f
C204 x7.x2.x2.CLK dvss 0.389657f
C205 x7.x5.TE_B dvss 4.59445f
C206 x7.x1.x4.Q dvss 0.100179f
C207 x7.x1.x3.Q dvss 0.092032f
C208 x7.x1.x2.Q dvss 0.092454f
C209 x7.x3.A2 dvss 5.765015f
C210 standby_33 dvss 11.159889f
C211 x4.in_b dvss 30.171328f
C212 x7.x1.x4.CLK dvss 0.511115f
C213 x7.x1.x3.CLK dvss 0.528314f
C214 x7.x1.x2.CLK dvss 0.382316f
C215 x7.x3.B2 dvss 5.822032f
C216 dout_ip dvss 15.022734f
C217 standby_ip dvss 21.272581f
C218 ena_ip dvss 23.378262f
C219 avdd_ip dvss 0.207998p
C220 dvss_ip dvss 60.189896f
C221 a_22601_n15524.t1 dvss 1.45f
C222 a_22601_n15524.t0 dvss 1.45f
C223 dout.t1 dvss 0.040138f
C224 dout.t0 dvss 0.223213f
C225 dout.n0 dvss 3.29562f
C226 x4.out_b.n0 dvss 5.53652f
C227 x4.out_b.t3 dvss 1.30743f
C228 x4.out_b.t1 dvss 0.044437f
C229 x4.out_b.t2 dvss 0.044437f
C230 x4.out_b.n1 dvss 0.140668f
C231 x4.out_b.t0 dvss 0.055178f
C232 dout_filt.n0 dvss 3.37345f
C233 dout_filt.t0 dvss 0.033084f
C234 dout_filt.n1 dvss 0.063466f
C235 dout_filt.t1 dvss 0.020119f
C236 dout_filt.n2 dvss 0.064349f
C237 dout_filt.t2 dvss 0.028544f
C238 dout_filt.t3 dvss 0.296603f
C239 dout_filt.t4 dvss 0.738515f
C240 vn.n1 dvss 1.00977f
C241 vn.n2 dvss 0.659335f
C242 vn.n3 dvss 0.85526f
C243 vn.t3 dvss 1.05137f
C244 vn.t5 dvss 1.15294f
C245 vn.t9 dvss 1.23617f
C246 vn.t8 dvss 1.05137f
C247 vn.n4 dvss 0.38691f
C248 vn.t2 dvss 0.047578f
C249 vn.t0 dvss 0.047578f
C250 vn.n5 dvss 0.099929f
C251 vn.t1 dvss 0.175661f
C252 vn.n6 dvss 0.536235f
C253 vn.t4 dvss 0.047578f
C254 vn.t6 dvss 0.047578f
C255 vn.n7 dvss 0.095156f
C256 vn.t7 dvss 0.166434f
C257 ena_33.n0 dvss 6.315629f
C258 ena_33.n1 dvss 0.292187f
C259 ena_33.n2 dvss 0.292479f
C260 ena_33.t5 dvss 0.411695f
C261 ena_33.t8 dvss 0.391709f
C262 ena_33.n3 dvss 0.294838f
C263 ena_33.t3 dvss 0.411399f
C264 ena_33.t6 dvss 0.391709f
C265 ena_33.n4 dvss 0.292479f
C266 ena_33.n5 dvss 0.557916f
C267 ena_33.t7 dvss 0.391709f
C268 ena_33.n6 dvss 0.126403f
C269 ena_33.n7 dvss 0.352232f
C270 ena_33.n8 dvss 0.884488f
C271 ena_33.t4 dvss 1.50033f
C272 ena_33.t0 dvss 0.050995f
C273 ena_33.t1 dvss 0.050995f
C274 ena_33.n9 dvss 0.161368f
C275 ena_33.t2 dvss 0.06332f
C276 vrb.t2 dvss 0.112245f
C277 vrb.t4 dvss 0.137391f
C278 vrb.n0 dvss 1.23688f
C279 vrb.t3 dvss 0.112257f
C280 vrb.t1 dvss 0.136226f
C281 vrb.n1 dvss 1.23886f
C282 vrb.t0 dvss 0.036259f
C283 vrb.n2 dvss 1.03965f
C284 vrb.n3 dvss 0.533375f
C285 vg2.n0 dvss 0.03576f
C286 vg2.n1 dvss 0.032988f
C287 vg2.t5 dvss 0.080953f
C288 vg2.n2 dvss 0.148193f
C289 vg2.n3 dvss 0.030952f
C290 vg2.n4 dvss 0.065976f
C291 vg2.t7 dvss 0.07945f
C292 vg2.n5 dvss 0.039561f
C293 vg2.n6 dvss 0.020508f
C294 vg2.n7 dvss 0.03576f
C295 vg2.n8 dvss 0.032988f
C296 vg2.t9 dvss 0.080949f
C297 vg2.n9 dvss 0.148053f
C298 vg2.n10 dvss 0.030952f
C299 vg2.n11 dvss 0.065976f
C300 vg2.t6 dvss 0.07945f
C301 vg2.n12 dvss 0.039706f
C302 vg2.n13 dvss 0.020508f
C303 vg2.n14 dvss 0.022657f
C304 vg2.t8 dvss 0.063882f
C305 vg2.t2 dvss 4.94472f
C306 vg2.t1 dvss 4.97221f
C307 vg2.t4 dvss 4.97221f
C308 vg2.t3 dvss 4.94281f
C309 vg2.n15 dvss 1.13816f
C310 vg2.n16 dvss 0.438266f
C311 vg2.n18 dvss 0.028457f
C312 xin.t21 dvss 0.018527f
C313 xin.t8 dvss 0.018041f
C314 xin.n0 dvss 0.133592f
C315 xin.n1 dvss 0.074808f
C316 xin.n2 dvss 0.074808f
C317 xin.n3 dvss 0.074808f
C318 xin.n4 dvss 0.074808f
C319 xin.n5 dvss 0.142348f
C320 xin.t18 dvss 0.148572f
C321 xin.t15 dvss 0.148502f
C322 xin.n6 dvss 0.142348f
C323 xin.n7 dvss 0.074808f
C324 xin.t13 dvss 0.148502f
C325 xin.n8 dvss 0.074808f
C326 xin.t19 dvss 0.148502f
C327 xin.n9 dvss 0.074808f
C328 xin.n10 dvss 0.074808f
C329 xin.t16 dvss 0.148502f
C330 xin.n11 dvss 0.074808f
C331 xin.t11 dvss 0.148502f
C332 xin.n12 dvss 0.074808f
C333 xin.n13 dvss 0.074808f
C334 xin.t10 dvss 0.148502f
C335 xin.n14 dvss 0.074808f
C336 xin.t17 dvss 0.148502f
C337 xin.n15 dvss 0.074808f
C338 xin.n16 dvss 0.074808f
C339 xin.t14 dvss 0.148502f
C340 xin.n17 dvss 0.074808f
C341 xin.t12 dvss 0.148502f
C342 xin.n18 dvss 0.074808f
C343 xin.n19 dvss 0.074808f
C344 xin.t9 dvss 0.148502f
C345 xin.n20 dvss 0.074808f
C346 xin.t6 dvss 0.148502f
C347 xin.n21 dvss 0.135448f
C348 xin.n22 dvss 0.606785f
C349 xin.n23 dvss 0.238527f
C350 xin.n24 dvss 0.241646f
C351 xin.n25 dvss 0.276924f
C352 xin.t20 dvss 0.570521f
C353 xin.n26 dvss 0.244557f
C354 xin.t7 dvss 0.570521f
C355 xin.n27 dvss 0.217057f
C356 xin.n28 dvss 0.161022f
C357 xin.n29 dvss 2.90223f
C358 xin.n30 dvss 3.49329f
C359 xin.n31 dvss 2.79271f
C360 xin.t2 dvss 44.0798f
C361 xin.t4 dvss 34.1562f
C362 xin.t1 dvss 34.0215f
C363 xin.t0 dvss 0.096027f
C364 xin.n32 dvss 3.69079f
C365 xin.n33 dvss 21.082699f
C366 xin.t5 dvss 24.1119f
C367 xin.n34 dvss 21.077301f
C368 xin.t3 dvss 24.088f
C369 xin.n35 dvss 21.08f
C370 xin.n36 dvss 2.91967f
C371 xin.n37 dvss 1.43525f
C372 xin.n38 dvss 0.571166f
C373 vg1.t3 dvss 0.052096f
C374 vg1.n0 dvss 0.412053f
C375 vg1.n1 dvss 0.135013f
C376 vg1.t1 dvss 0.248955f
C377 vg1.t5 dvss 0.32393f
C378 vg1.n2 dvss 0.210078f
C379 vg1.t2 dvss 0.044909f
C380 vg1.n3 dvss 0.263389f
C381 vg1.n4 dvss 0.067733f
C382 vg1.t8 dvss 42.208103f
C383 vg1.t9 dvss 42.9209f
C384 vg1.t4 dvss 21.9912f
C385 vg1.n5 dvss 21.955198f
C386 vg1.t7 dvss 21.9912f
C387 vg1.n6 dvss 21.5232f
C388 vg1.t6 dvss 21.9912f
C389 vg1.n7 dvss 11.900599f
C390 vg1.n8 dvss 13.9559f
C391 vg1.t0 dvss 0.012376f
C392 vg1.n9 dvss 2.83328f
C393 vg1.n10 dvss 1.38457f
C394 vg1.n11 dvss 0.103037f
C395 vg1.n12 dvss 0.393913f
C396 ena_b_33.n0 dvss 0.984134f
C397 ena_b_33.n1 dvss 6.57801f
C398 ena_b_33.n2 dvss 0.299431f
C399 ena_b_33.t6 dvss 0.400911f
C400 ena_b_33.t8 dvss 0.421207f
C401 ena_b_33.t4 dvss 0.420861f
C402 ena_b_33.t7 dvss 0.400911f
C403 ena_b_33.n3 dvss 0.299431f
C404 ena_b_33.n4 dvss 0.565594f
C405 ena_b_33.n5 dvss 0.30181f
C406 ena_b_33.t3 dvss 0.400911f
C407 ena_b_33.n6 dvss 0.30181f
C408 ena_b_33.n7 dvss 0.482654f
C409 ena_b_33.t5 dvss 1.5126f
C410 ena_b_33.t0 dvss 0.05141f
C411 ena_b_33.t1 dvss 0.05141f
C412 ena_b_33.n8 dvss 0.162741f
C413 ena_b_33.t2 dvss 0.063836f
C414 avdd.n0 dvss 0.482001f
C415 avdd.t5 dvss 0.033339f
C416 avdd.n1 dvss 1.66082f
C417 avdd.n2 dvss 0.05952f
C418 avdd.n3 dvss 0.055259f
C419 avdd.n4 dvss 0.08282f
C420 avdd.n5 dvss 0.57254f
C421 avdd.n6 dvss 1.01205f
C422 avdd.n7 dvss 1.01205f
C423 avdd.t2 dvss 0.875283f
C424 avdd.t17 dvss 0.687077f
C425 avdd.t6 dvss 0.875283f
C426 avdd.t13 dvss 0.687077f
C427 avdd.n8 dvss 0.452172f
C428 avdd.t9 dvss 7.37116f
C429 avdd.n9 dvss 7.35034f
C430 avdd.t8 dvss 8.92008f
C431 avdd.t11 dvss 7.09459f
C432 avdd.n10 dvss 7.54853f
C433 avdd.t10 dvss 8.96278f
C434 avdd.n11 dvss 3.6056f
C435 avdd.n12 dvss 0.751718f
C436 avdd.n13 dvss 0.567021f
C437 avdd.n14 dvss 0.547944f
C438 avdd.n15 dvss 0.345317f
C439 avdd.n16 dvss 0.477166f
C440 avdd.n17 dvss 3.66554f
C441 avdd.n18 dvss 0.715165f
C442 avdd.t14 dvss 0.036186f
C443 avdd.t7 dvss 0.036186f
C444 avdd.n19 dvss 0.088691f
C445 avdd.t18 dvss 0.036186f
C446 avdd.t16 dvss 0.036186f
C447 avdd.n20 dvss 0.088691f
C448 avdd.n21 dvss 1.89167f
C449 avdd.n22 dvss 0.946075f
C450 avdd.t3 dvss 0.13224f
C451 avdd.n23 dvss 0.335803f
C452 avdd.n24 dvss 5.54098f
C453 avdd.n25 dvss 0.872611f
C454 avdd.n26 dvss 1.16121f
C455 avdd.n27 dvss 1.16121f
C456 avdd.n28 dvss 4.35756f
C457 avdd.n29 dvss 1.29639f
C458 avdd.n30 dvss 0.088681f
C459 avdd.n31 dvss 0.070403f
C460 avdd.n32 dvss 0.532281f
C461 avdd.n33 dvss 1.52809f
C462 avdd.t1 dvss 0.033339f
C463 avdd.n34 dvss 1.43378f
C464 avdd.n35 dvss 0.105027f
C465 avdd.n36 dvss 0.105573f
C466 avdd.n37 dvss 0.154685f
C467 avdd.t0 dvss 2.45528f
C468 avdd.n38 dvss 0.070403f
C469 avdd.n39 dvss 0.101864f
C470 avdd.n40 dvss 0.105573f
C471 avdd.n41 dvss 0.54455f
C472 avdd.t12 dvss 0.033339f
C473 avdd.n42 dvss 0.022804f
C474 avdd.n43 dvss 0.672007f
C475 avdd.n44 dvss 1.4511f
C476 avdd.n45 dvss 1.11231f
C477 avdd.n46 dvss 0.724468f
C478 avdd.n47 dvss 2.40543f
C479 avdd.n48 dvss 3.34797f
C480 avdd.n49 dvss 1.13035f
C481 avdd.n50 dvss 0.352457f
C482 avdd.n51 dvss 0.307059f
C483 avdd.n52 dvss 0.10386f
C484 avdd.n53 dvss 1.64194f
C485 avdd.n54 dvss 0.10386f
C486 avdd.n55 dvss 0.154685f
C487 avdd.n56 dvss 0.088681f
C488 avdd.n57 dvss 0.061522f
C489 avdd.n58 dvss 0.10386f
C490 avdd.n59 dvss 1.64194f
C491 avdd.n60 dvss 0.10386f
C492 avdd.n61 dvss 0.05952f
C493 avdd.n62 dvss 0.114361f
C494 avdd.n63 dvss 0.703461f
C495 avdd.n64 dvss 1.34899f
C496 avdd.n65 dvss 1.44f
C497 avdd.t19 dvss 0.033339f
C498 avdd.n66 dvss 1.40397f
C499 avdd.n67 dvss 0.355639f
C500 avdd.n68 dvss 0.105573f
C501 avdd.n69 dvss 0.154685f
C502 avdd.t4 dvss 2.45528f
C503 avdd.n70 dvss 0.101864f
C504 avdd.n71 dvss 0.105573f
C505 avdd.n72 dvss 0.105027f
C506 avdd.n73 dvss 0.061522f
C507 avdd.n74 dvss 0.10386f
C508 avdd.n75 dvss 1.64194f
C509 avdd.n76 dvss 0.10386f
C510 avdd.n77 dvss 0.154685f
C511 avdd.n78 dvss 0.10386f
C512 avdd.n79 dvss 1.64194f
C513 avdd.n80 dvss 0.10386f
C514 avdd.n81 dvss 0.303824f
C515 avdd.n82 dvss 0.711278f
C516 avdd.n83 dvss 1.90791f
C517 avdd.n84 dvss 4.04344f
C518 avdd.n85 dvss 0.691895f
C519 avdd.n86 dvss 0.469079f
C520 avdd.n87 dvss 1.29149f
C521 avdd.n88 dvss 1.28783f
C522 avdd.n89 dvss 0.441283f
C523 avdd.n90 dvss 1.16292f
C524 avdd.n91 dvss 4.37865f
C525 avdd.n92 dvss 4.35756f
C526 avdd.n93 dvss 4.37865f
C527 avdd.n94 dvss 1.16292f
C528 avdd.n95 dvss 0.641325f
C529 avdd.n96 dvss 3.16932f
C530 avdd.n97 dvss 0.204843f
C531 avdd.t15 dvss 0.687077f
C532 avdd.n98 dvss 0.204843f
C533 avdd.n99 dvss 0.715578f
C534 avdd.n100 dvss 0.611329f
C535 avdd.n101 dvss 0.143723f
C536 avdd.n102 dvss 0.056349f
C537 avdd.n103 dvss 0.296365f
C538 avss.n0 dvss 0.259025f
C539 avss.n1 dvss 0.275848f
C540 avss.t25 dvss 0.059315f
C541 avss.n2 dvss 0.188304f
C542 avss.n3 dvss 0.025591f
C543 avss.n4 dvss 0.097042f
C544 avss.n5 dvss 0.087001f
C545 avss.n6 dvss 0.087001f
C546 avss.t24 dvss 0.417521f
C547 avss.t22 dvss 0.417521f
C548 avss.n7 dvss 0.041818f
C549 avss.n8 dvss 0.074102f
C550 avss.t23 dvss 0.059553f
C551 avss.t11 dvss 0.059553f
C552 avss.n9 dvss 0.784978f
C553 avss.n10 dvss 0.110883f
C554 avss.t17 dvss 0.059315f
C555 avss.t13 dvss 0.059315f
C556 avss.n11 dvss 0.472749f
C557 avss.n12 dvss 0.04178f
C558 avss.n13 dvss 0.088476f
C559 avss.n14 dvss 0.088476f
C560 avss.n15 dvss 0.479005f
C561 avss.n16 dvss 0.087001f
C562 avss.n17 dvss 0.479005f
C563 avss.t10 dvss 0.417521f
C564 avss.n18 dvss 0.225919f
C565 avss.t12 dvss 0.417521f
C566 avss.n19 dvss 3.07761f
C567 avss.n20 dvss 6.9069f
C568 avss.t16 dvss 0.417521f
C569 avss.n21 dvss 0.088476f
C570 avss.n22 dvss 0.088476f
C571 avss.n23 dvss 0.074102f
C572 avss.n24 dvss 0.14364f
C573 avss.n25 dvss 0.087001f
C574 avss.n26 dvss 0.087001f
C575 avss.n27 dvss 0.225919f
C576 avss.t18 dvss 0.417521f
C577 avss.n28 dvss 0.087001f
C578 avss.n29 dvss 0.479005f
C579 avss.n30 dvss 0.479005f
C580 avss.t0 dvss 0.417521f
C581 avss.t2 dvss 0.417521f
C582 avss.n31 dvss 0.041818f
C583 avss.t19 dvss 0.059553f
C584 avss.t1 dvss 0.059553f
C585 avss.t3 dvss 0.059315f
C586 avss.n32 dvss 0.075425f
C587 avss.n33 dvss 0.453458f
C588 avss.n34 dvss 0.073465f
C589 avss.n35 dvss 0.1253f
C590 avss.n36 dvss 2.78849f
C591 avss.t20 dvss 0.809304f
C592 avss.t14 dvss 0.689326f
C593 avss.n37 dvss 2.02175f
C594 avss.n38 dvss 1.63265f
C595 avss.t6 dvss 0.783127f
C596 avss.t4 dvss 0.689326f
C597 avss.n39 dvss 0.125508f
C598 avss.t8 dvss 0.689326f
C599 avss.n40 dvss 0.125508f
C600 avss.n41 dvss 0.075425f
C601 avss.t7 dvss 0.076187f
C602 avss.n42 dvss 0.481111f
C603 avss.t9 dvss 0.022354f
C604 avss.t5 dvss 0.022354f
C605 avss.n43 dvss 0.07455f
C606 avss.t21 dvss 0.022354f
C607 avss.t15 dvss 0.022354f
C608 avss.n44 dvss 0.081002f
C609 avss.n45 dvss 1.28451f
C610 avss.n46 dvss 0.976711f
C611 avss.t26 dvss 7.70817f
C612 avss.n47 dvss 7.26208f
C613 avss.t29 dvss 7.70817f
C614 avss.n48 dvss 7.55356f
C615 avss.t28 dvss 7.70817f
C616 avss.n49 dvss 7.45534f
C617 avss.n50 dvss 3.788f
C618 avss.t27 dvss 7.70817f
C619 avss.n51 dvss 2.0569f
C620 avss.n52 dvss 4.69347f
C621 avss.n53 dvss 1.74716f
C622 avss.n54 dvss 1.83304f
C623 avss.n55 dvss 1.74559f
C624 avss.n56 dvss 0.089885f
C625 avss.n57 dvss 0.214326f
C626 avss.n58 dvss 0.250065f
C627 avss.n59 dvss 0.607011f
C628 avss.n60 dvss 0.259025f
C629 avss.n61 dvss 0.33435f
C630 avss.n62 dvss 0.074102f
C631 avss.n63 dvss 0.09708f
C632 avss.n64 dvss 0.025591f
C633 avss.n65 dvss 0.034883f
C634 avss.n66 dvss 0.088476f
C635 avss.n67 dvss 0.225919f
C636 avss.n68 dvss 0.088476f
C637 avss.n69 dvss 0.03485f
C638 avss.n70 dvss 0.097042f
C639 avss.n71 dvss 0.04178f
C640 avss.n72 dvss 0.110805f
C641 avss.n73 dvss 0.087001f
C642 avss.n74 dvss 0.752109f
C643 avss.n75 dvss 1.87691f
C644 avss.n76 dvss 0.752109f
C645 avss.n77 dvss 0.087001f
C646 avss.n78 dvss 0.110805f
C647 avss.n79 dvss 0.110883f
C648 avss.n80 dvss 0.429808f
C649 avss.n81 dvss 1.13806f
C650 avss.n82 dvss 0.538123f
C651 avss.n83 dvss 0.33435f
C652 avss.n84 dvss 0.074102f
C653 avss.n85 dvss 0.09708f
C654 avss.n86 dvss 0.034883f
C655 avss.n87 dvss 0.088476f
C656 avss.n88 dvss 0.225919f
C657 avss.n89 dvss 0.088476f
C658 avss.n90 dvss 0.03485f
C659 avss.n91 dvss 0.14364f
C660 avss.n92 dvss 0.083634f
C661 avss.n93 dvss 0.15294f
C662 avss.n94 dvss 0.227923f
C663 standby_ip.n0 dvss 3.29304f
C664 standby_ip.n1 dvss 0.852877f
C665 standby_ip.n2 dvss 0.630392f
C666 standby_ip.n3 dvss 0.097579f
C667 standby_ip.n7 dvss 0.113896f
C668 standby_ip.n9 dvss 0.109598f
C669 standby_ip.n11 dvss 0.113896f
C670 standby_ip.n14 dvss 0.108447f
C671 standby_ip.t0 dvss 0.020746f
C672 standby_ip.t1 dvss 0.029835f
C673 standby_ip.t3 dvss 0.019244f
C674 standby_ip.t14 dvss 0.012026f
C675 standby_ip.n15 dvss 0.034453f
C676 standby_ip.n16 dvss 0.061012f
C677 standby_ip.t10 dvss 0.94678f
C678 standby_ip.n17 dvss 0.113896f
C679 standby_ip.t6 dvss 0.291364f
C680 standby_ip.n18 dvss 0.113896f
C681 standby_ip.t5 dvss 0.291364f
C682 standby_ip.t17 dvss 0.291364f
C683 standby_ip.n19 dvss 0.113896f
C684 standby_ip.n20 dvss 0.113896f
C685 standby_ip.t12 dvss 0.291364f
C686 standby_ip.n21 dvss 0.113896f
C687 standby_ip.n22 dvss 0.116158f
C688 standby_ip.n23 dvss 0.113896f
C689 standby_ip.t9 dvss 0.291364f
C690 standby_ip.n24 dvss 0.113896f
C691 standby_ip.t15 dvss 0.294612f
C692 standby_ip.n25 dvss 0.116227f
C693 standby_ip.n26 dvss 0.113896f
C694 standby_ip.t8 dvss 0.291364f
C695 standby_ip.n27 dvss 0.113896f
C696 standby_ip.n28 dvss 0.113896f
C697 standby_ip.t11 dvss 0.291364f
C698 standby_ip.n29 dvss 0.113896f
C699 standby_ip.n30 dvss 0.113896f
C700 standby_ip.t18 dvss 0.291364f
C701 standby_ip.n31 dvss 0.113896f
C702 standby_ip.n32 dvss 0.113896f
C703 standby_ip.t4 dvss 0.294685f
C704 standby_ip.t2 dvss 0.26673f
C705 standby_ip.n33 dvss 0.230886f
C706 standby_ip.t13 dvss 0.241192f
C707 standby_ip.t7 dvss 0.241004f
C708 standby_ip.n34 dvss 0.202569f
C709 standby_ip.n35 dvss 0.931655f
C710 standby_ip.t16 dvss 0.275696f
C711 standby_ip.n36 dvss 0.125129f
C712 a_17576_n6897.t0 dvss 0.195122p
C713 a_17576_n6897.n0 dvss 0.083483f
C714 a_17576_n6897.t1 dvss 0.184195f
C715 a_17576_n6897.t2 dvss 0.067412f
C716 a_17576_n6897.n1 dvss 0.085831f
C717 a_17576_n6897.t3 dvss 0.190371f
C718 a_17576_n6897.t4 dvss 0.066238f
C719 dout_ip.t0 dvss 0.022607f
C720 dout_ip.t3 dvss 0.021864f
C721 dout_ip.t2 dvss 0.021852f
C722 dout_ip.t4 dvss 0.023836f
C723 dout_ip.t10 dvss 0.01616f
C724 dout_ip.n0 dvss 0.038785f
C725 dout_ip.t7 dvss 0.012534f
C726 dout_ip.n1 dvss 0.033243f
C727 dout_ip.n2 dvss 0.027616f
C728 dout_ip.n3 dvss 0.027616f
C729 dout_ip.t6 dvss 0.012534f
C730 dout_ip.n4 dvss 0.033243f
C731 dout_ip.n5 dvss 0.35872f
C732 dout_ip.n6 dvss 0.352547f
C733 dout_ip.t1 dvss 0.022607f
C734 inv_m1.t0 dvss 0.046283f
C735 inv_m1.n0 dvss 0.469196f
C736 inv_m1.n1 dvss 0.129403f
C737 inv_m1.t5 dvss 0.362679f
C738 inv_m1.t2 dvss 0.36268f
C739 inv_m1.n2 dvss 0.117551f
C740 inv_m1.t4 dvss 0.340571f
C741 inv_m1.t3 dvss 0.340573f
C742 inv_m1.n3 dvss 3.00164f
C743 inv_m1.t1 dvss 0.044738f
C744 inv_m1.n4 dvss 0.57064f
C745 inv_m1.n5 dvss 0.723313f
C746 inv_m1.n6 dvss 0.280865f
C747 inv_m1.n7 dvss 0.038196f
C748 inv_m1.n8 dvss 0.093067f
C749 inv_in.t3 dvss 0.656506f
C750 inv_in.t11 dvss 5.66972f
C751 inv_in.n0 dvss 5.16758f
C752 inv_in.t5 dvss 5.51881f
C753 inv_in.n1 dvss 2.61945f
C754 inv_in.t6 dvss 5.51881f
C755 inv_in.n2 dvss 2.65659f
C756 inv_in.n3 dvss 2.79157f
C757 inv_in.t14 dvss 5.51881f
C758 inv_in.n4 dvss 5.28337f
C759 inv_in.t12 dvss 5.54244f
C760 inv_in.n5 dvss 5.27646f
C761 inv_in.t13 dvss 5.51881f
C762 inv_in.n6 dvss 2.65659f
C763 inv_in.t9 dvss 5.57337f
C764 inv_in.n7 dvss 5.38886f
C765 inv_in.t10 dvss 5.57337f
C766 inv_in.t2 dvss 5.57337f
C767 inv_in.n8 dvss 5.25688f
C768 inv_in.n9 dvss 5.39873f
C769 inv_in.t4 dvss 5.51881f
C770 inv_in.n10 dvss 2.65659f
C771 inv_in.n11 dvss 2.89677f
C772 inv_in.n12 dvss 2.75493f
C773 inv_in.t8 dvss 5.51881f
C774 inv_in.n13 dvss 2.61945f
C775 inv_in.n14 dvss 2.75985f
C776 inv_in.n15 dvss 2.75985f
C777 inv_in.n16 dvss 2.75695f
C778 inv_in.t7 dvss 5.51881f
C779 inv_in.n17 dvss 5.4492f
C780 inv_in.n18 dvss 0.821552f
C781 inv_in.t0 dvss 0.112287f
C782 inv_in.t1 dvss 0.646679f
C783 inv_in.n19 dvss 2.21037f
C784 xout.t26 dvss 0.031623f
C785 xout.t24 dvss 0.032499f
C786 xout.t18 dvss 0.162965f
C787 xout.t20 dvss 0.162965f
C788 xout.n0 dvss 1.30069f
C789 xout.t17 dvss 0.162965f
C790 xout.t19 dvss 0.162965f
C791 xout.n1 dvss 0.919705f
C792 xout.n2 dvss 3.69834f
C793 xout.t16 dvss 0.164923f
C794 xout.n3 dvss 0.36174f
C795 xout.t14 dvss 0.164923f
C796 xout.n4 dvss 0.36234f
C797 xout.t21 dvss 0.162965f
C798 xout.n5 dvss 0.557313f
C799 xout.t22 dvss 0.162965f
C800 xout.n6 dvss 0.557313f
C801 xout.n7 dvss 0.711321f
C802 xout.n8 dvss 0.782198f
C803 xout.n9 dvss 0.780269f
C804 xout.n10 dvss 4.25798f
C805 xout.n11 dvss 2.51745f
C806 xout.t12 dvss 0.162965f
C807 xout.t11 dvss 0.162965f
C808 xout.n12 dvss 0.776049f
C809 xout.n13 dvss 0.782941f
C810 xout.t15 dvss 0.162965f
C811 xout.t13 dvss 0.162965f
C812 xout.n14 dvss 0.776049f
C813 xout.n15 dvss 0.781535f
C814 xout.n16 dvss 0.833328f
C815 xout.t6 dvss 0.044594f
C816 xout.t7 dvss 0.044594f
C817 xout.n17 dvss 0.151768f
C818 xout.t9 dvss 0.044594f
C819 xout.t4 dvss 0.044594f
C820 xout.n18 dvss 0.145391f
C821 xout.t8 dvss 0.044594f
C822 xout.t0 dvss 0.044594f
C823 xout.n19 dvss 0.153068f
C824 xout.n20 dvss 2.99948f
C825 xout.t10 dvss 0.044594f
C826 xout.t2 dvss 0.044594f
C827 xout.n21 dvss 0.145391f
C828 xout.t5 dvss 0.044594f
C829 xout.t3 dvss 0.044594f
C830 xout.n22 dvss 0.099654f
C831 xout.n23 dvss 1.98386f
C832 xout.n24 dvss 2.32242f
C833 xout.n25 dvss 2.77708f
C834 xout.t1 dvss 0.060812f
C835 xout.n26 dvss 2.6875f
C836 xout.n27 dvss 0.418318f
C837 xout.n28 dvss 0.423788f
C838 xout.n29 dvss 0.485658f
C839 xout.t23 dvss 1.00055f
C840 xout.n30 dvss 0.428893f
C841 xout.t25 dvss 1.00055f
C842 xout.n31 dvss 0.380665f
C843 xout.n32 dvss 0.282855f
C844 xout.n33 dvss 5.34696f
C845 xout.n34 dvss 6.45162f
C846 xout.n35 dvss 1.6717f
C847 avdd_ip.n0 dvss 0.60907f
C848 avdd_ip.n1 dvss 0.975189f
C849 avdd_ip.n2 dvss 0.568516f
C850 avdd_ip.n3 dvss 1.23782f
C851 avdd_ip.n4 dvss 1.23782f
C852 avdd_ip.n5 dvss 4.75695f
C853 avdd_ip.n6 dvss 0.785548f
C854 avdd_ip.t20 dvss 0.039571f
C855 avdd_ip.n7 dvss 0.146289f
C856 avdd_ip.n8 dvss 0.169741f
C857 avdd_ip.n9 dvss 2.27671f
C858 avdd_ip.t28 dvss 0.039571f
C859 avdd_ip.t22 dvss 0.039571f
C860 avdd_ip.n10 dvss 0.311255f
C861 avdd_ip.t27 dvss 0.039571f
C862 avdd_ip.t19 dvss 0.039571f
C863 avdd_ip.n11 dvss 0.188441f
C864 avdd_ip.n12 dvss 0.239694f
C865 avdd_ip.t5 dvss 0.010828f
C866 avdd_ip.t3 dvss 0.010828f
C867 avdd_ip.n13 dvss 0.02654f
C868 avdd_ip.t0 dvss 0.010828f
C869 avdd_ip.t6 dvss 0.010828f
C870 avdd_ip.n14 dvss 0.028004f
C871 avdd_ip.t1 dvss 0.044012f
C872 avdd_ip.n15 dvss 0.302781f
C873 avdd_ip.n16 dvss 0.649109f
C874 avdd_ip.t33 dvss 29.2301f
C875 avdd_ip.n17 dvss 6.11247f
C876 avdd_ip.n18 dvss 4.52625f
C877 avdd_ip.t30 dvss 1.82962f
C878 avdd_ip.n19 dvss 1.16812f
C879 avdd_ip.t31 dvss 1.82962f
C880 avdd_ip.n20 dvss 1.12616f
C881 avdd_ip.n21 dvss 1.48398f
C882 avdd_ip.t29 dvss 1.82962f
C883 avdd_ip.n22 dvss 1.64206f
C884 avdd_ip.t32 dvss 1.82962f
C885 avdd_ip.n23 dvss 1.63866f
C886 avdd_ip.n24 dvss 1.60189f
C887 avdd_ip.n25 dvss 4.18817f
C888 avdd_ip.n26 dvss 6.1263f
C889 avdd_ip.n27 dvss 0.072597f
C890 avdd_ip.n28 dvss 1.02884f
C891 avdd_ip.t21 dvss 0.039571f
C892 avdd_ip.n29 dvss 0.1983f
C893 avdd_ip.t23 dvss 0.040722f
C894 avdd_ip.n30 dvss 0.238511f
C895 avdd_ip.t25 dvss 0.039571f
C896 avdd_ip.n31 dvss 0.146289f
C897 avdd_ip.t26 dvss 0.039571f
C898 avdd_ip.n32 dvss 0.197546f
C899 avdd_ip.t24 dvss 0.040771f
C900 avdd_ip.n33 dvss 0.116402f
C901 avdd_ip.n34 dvss 0.239694f
C902 avdd_ip.n35 dvss 1.71745f
C903 avdd_ip.n36 dvss 0.946073f
C904 avdd_ip.t18 dvss 0.039571f
C905 avdd_ip.t17 dvss 0.039571f
C906 avdd_ip.n37 dvss 0.311247f
C907 avdd_ip.t16 dvss 0.039571f
C908 avdd_ip.t14 dvss 0.039571f
C909 avdd_ip.n38 dvss 0.188729f
C910 avdd_ip.n39 dvss 0.239802f
C911 avdd_ip.n40 dvss 0.977469f
C912 avdd_ip.n41 dvss 0.780191f
C913 avdd_ip.n42 dvss 1.81869f
C914 avdd_ip.n43 dvss 1.22909f
C915 avdd_ip.n44 dvss 1.11439f
C916 avdd_ip.n45 dvss 2.2026f
C917 avdd_ip.n46 dvss 2.2026f
C918 avdd_ip.t7 dvss 2.80357f
C919 avdd_ip.t8 dvss 0.039571f
C920 avdd_ip.t9 dvss 0.039571f
C921 avdd_ip.t10 dvss 0.039571f
C922 avdd_ip.n47 dvss 0.499823f
C923 avdd_ip.t12 dvss 0.039571f
C924 avdd_ip.t13 dvss 0.039571f
C925 avdd_ip.t15 dvss 0.039571f
C926 avdd_ip.n48 dvss 0.239694f
C927 avdd_ip.n49 dvss 1.0546f
C928 avdd_ip.n50 dvss 0.110378f
C929 avdd_ip.n51 dvss 0.203213f
C930 avdd_ip.t11 dvss 2.80357f
C931 avdd_ip.n52 dvss 2.39957f
C932 avdd_ip.n53 dvss 0.203213f
C933 avdd_ip.n54 dvss 0.41208f
C934 avdd_ip.n55 dvss 0.629324f
C935 avdd_ip.n56 dvss 1.0246f
C936 avdd_ip.n57 dvss 0.419429f
C937 avdd_ip.n58 dvss 1.23612f
C938 avdd_ip.n59 dvss 4.73082f
C939 avdd_ip.n60 dvss 4.75695f
C940 avdd_ip.n61 dvss 4.73082f
C941 avdd_ip.n62 dvss 1.23612f
C942 avdd_ip.n63 dvss 0.40817f
C943 avdd_ip.n64 dvss 0.011754f
C944 avdd_ip.n70 dvss 0.039931f
C945 avdd_ip.t4 dvss 0.061763f
C946 avdd_ip.n73 dvss 0.039931f
C947 avdd_ip.n76 dvss 0.381639f
C948 avdd_ip.n77 dvss 0.011227f
C949 avdd_ip.t2 dvss 0.053089f
C950 avdd_ip.n82 dvss -3.33095f
C951 avdd_ip.n83 dvss 3.37127f
C952 avdd_ip.n87 dvss 0.039931f
C953 avdd_ip.n90 dvss 0.339621f
C954 avdd_ip.n91 dvss 0.447224f
C955 avdd_ip.n92 dvss 0.881006f
C956 avdd_ip.n93 dvss 3.97624f
C957 a_10658_n5446.n0 dvss 12.804701f
C958 a_10658_n5446.t13 dvss 0.728619f
C959 a_10658_n5446.t2 dvss 0.719247f
C960 a_10658_n5446.t3 dvss 0.086698f
C961 a_10658_n5446.t7 dvss 0.086698f
C962 a_10658_n5446.t1 dvss 0.086698f
C963 a_10658_n5446.t0 dvss 0.719247f
C964 a_10658_n5446.t11 dvss 0.728627f
C965 a_10658_n5446.t4 dvss 0.71925f
C966 a_10658_n5446.t5 dvss 0.086698f
C967 a_10658_n5446.t9 dvss 0.086698f
C968 a_10658_n5446.t8 dvss 0.71925f
C969 a_10658_n5446.t12 dvss 0.72111f
C970 a_10658_n5446.t6 dvss 0.719247f
C971 a_10658_n5446.t10 dvss 0.287197f
C972 standby_33.n0 dvss 7.35104f
C973 standby_33.t3 dvss 0.807828f
C974 standby_33.t4 dvss 1.63225f
C975 standby_33.t2 dvss 0.055479f
C976 standby_33.t1 dvss 0.055479f
C977 standby_33.n1 dvss 0.175556f
C978 standby_33.t0 dvss 0.068888f
C979 x7.x3.B2.t1 dvss 0.052533f
C980 x7.x3.B2.t0 dvss 0.066515f
C981 x7.x3.B2.t3 dvss 0.032856f
C982 x7.x3.B2.t2 dvss 0.020632f
C983 x7.x3.B2.n0 dvss 0.044446f
C984 x7.x3.B2.n1 dvss 0.160205f
C985 x7.x3.B2.t4 dvss 0.017992f
C986 x7.x3.B2.n2 dvss 0.051591f
C987 x7.x3.B2.t7 dvss 0.018195f
C988 x7.x3.B2.n3 dvss 0.056022f
C989 x7.x3.B2.n4 dvss 0.0112f
C990 x7.x3.B2.n5 dvss 0.058083f
C991 x7.x3.B2.t6 dvss 0.024488f
C992 x7.x3.B2.t5 dvss 0.026956f
C993 x7.x3.B2.n6 dvss 0.077088f
C994 x7.x3.B2.n7 dvss 1.89977f
C995 x7.x3.B2.n8 dvss 0.075188f
C996 a_9120_n9346.t3 dvss 0.027446f
C997 a_9120_n9346.t2 dvss 1.80482f
C998 a_9120_n9346.n0 dvss 2.79699f
C999 a_9120_n9346.t0 dvss 2.03504f
C1000 a_9120_n9346.t1 dvss 0.02735f
C1001 a_9120_n9346.n1 dvss 4.42071f
C1002 a_9120_n9346.t4 dvss 0.087656f
C1003 x4.in_b.n0 dvss 4.20129f
C1004 x4.in_b.n1 dvss 0.195939f
C1005 x4.in_b.n2 dvss 0.166239f
C1006 x4.in_b.n3 dvss 0.166517f
C1007 x4.in_b.n4 dvss 0.155263f
C1008 x4.in_b.t12 dvss 0.184865f
C1009 x4.in_b.t4 dvss 0.184721f
C1010 x4.in_b.t16 dvss 0.222927f
C1011 x4.in_b.t3 dvss 0.223807f
C1012 x4.in_b.t18 dvss 0.222094f
C1013 x4.in_b.t23 dvss 0.223668f
C1014 x4.in_b.t17 dvss 0.222037f
C1015 x4.in_b.t19 dvss 0.222448f
C1016 x4.in_b.t7 dvss 0.222043f
C1017 x4.in_b.t21 dvss 0.223667f
C1018 x4.in_b.t0 dvss 0.223807f
C1019 x4.in_b.t6 dvss 0.222526f
C1020 x4.in_b.t14 dvss 0.014284f
C1021 x4.in_b.n5 dvss 0.025334f
C1022 x4.in_b.t25 dvss 0.014284f
C1023 x4.in_b.n7 dvss 0.025334f
C1024 x4.in_b.t11 dvss 0.014284f
C1025 x4.in_b.n9 dvss 0.025334f
C1026 x4.in_b.t2 dvss 0.012433f
C1027 x4.in_b.n11 dvss 0.024252f
C1028 x4.in_b.t15 dvss 0.012433f
C1029 x4.in_b.n12 dvss 0.024252f
C1030 x4.in_b.t13 dvss 0.012433f
C1031 x4.in_b.n13 dvss 0.024252f
C1032 x4.in_b.t24 dvss 0.014864f
C1033 x4.in_b.n14 dvss 0.022789f
C1034 tail.n0 dvss 1.91477f
C1035 tail.t0 dvss 0.059783f
C1036 tail.t1 dvss 0.059783f
C1037 tail.n1 dvss 0.130872f
C1038 tail.n2 dvss 10.8565f
C1039 tail.t2 dvss 0.109992f
C1040 tail.t7 dvss 0.109992f
C1041 tail.n3 dvss 0.398074f
C1042 tail.t9 dvss 0.109992f
C1043 tail.t4 dvss 0.109992f
C1044 tail.n4 dvss 0.440953f
C1045 tail.t6 dvss 0.109992f
C1046 tail.t11 dvss 0.109992f
C1047 tail.n5 dvss 0.454375f
C1048 tail.t5 dvss 0.109992f
C1049 tail.t10 dvss 0.109992f
C1050 tail.n6 dvss 0.434225f
C1051 tail.t8 dvss 0.109992f
C1052 tail.t3 dvss 0.109992f
C1053 tail.n7 dvss 0.399316f
C1054 dvdd_ip.n0 dvss 0.105612f
C1055 dvdd_ip.n1 dvss 0.107411f
C1056 dvdd_ip.n2 dvss 0.170539f
C1057 dvdd_ip.n3 dvss 27.5155f
C1058 dvdd_ip.n4 dvss 8.99732f
C1059 dvdd_ip.n5 dvss 13.391299f
C1060 dvdd_ip.n6 dvss 9.85327f
C1061 dvdd_ip.n7 dvss 9.74982f
C1062 dvdd_ip.n8 dvss 9.74982f
C1063 dvdd_ip.n9 dvss 0.971823f
C1064 dvdd_ip.n10 dvss 9.85327f
C1065 dvdd_ip.n11 dvss 0.748792f
C1066 dvdd_ip.t56 dvss 0.423533p
C1067 dvdd_ip.n12 dvss 0.295713f
C1068 dvdd_ip.n13 dvss 0.708023f
C1069 dvdd_ip.t46 dvss 0.160415f
C1070 dvdd_ip.n14 dvss 12.7264f
C1071 dvdd_ip.n15 dvss 0.17054f
C1072 dvdd_ip.n16 dvss 0.112539f
C1073 dvdd_ip.n17 dvss 0.852304f
C1074 dvdd_ip.n18 dvss 0.528217f
C1075 dvdd_ip.n19 dvss 0.713054f
C1076 dvdd_ip.n20 dvss 6.80705f
C1077 dvdd_ip.n21 dvss 0.853678f
C1078 dvdd_ip.n22 dvss 0.45297f
C1079 dvdd_ip.n23 dvss 1.39412f
C1080 dvdd_ip.n24 dvss 0.538522f
C1081 dvdd_ip.n25 dvss 0.62375f
C1082 dvdd_ip.n26 dvss 0.013162f
C1083 dvdd_ip.n27 dvss 0.62919f
C1084 dvdd_ip.n29 dvss 3.02381f
C1085 dvdd_ip.n30 dvss 1.62374f
C1086 dvdd_ip.t31 dvss 0.05161f
C1087 dvdd_ip.n31 dvss 0.277899f
C1088 dvdd_ip.n32 dvss 1.12529f
C1089 dvdd_ip.t30 dvss 0.310004f
C1090 dvdd_ip.t39 dvss 0.160415f
C1091 dvdd_ip.t49 dvss 0.310004f
C1092 dvdd_ip.t50 dvss 0.32951f
C1093 dvdd_ip.n33 dvss 0.883458f
C1094 dvdd_ip.n34 dvss 0.248032f
C1095 dvdd_ip.t25 dvss 0.05161f
C1096 dvdd_ip.n35 dvss 0.524291f
C1097 dvdd_ip.t26 dvss 0.05161f
C1098 dvdd_ip.n36 dvss 0.258886f
C1099 dvdd_ip.t41 dvss 0.052512f
C1100 dvdd_ip.t32 dvss 0.05161f
C1101 dvdd_ip.n37 dvss 0.277899f
C1102 dvdd_ip.t33 dvss 0.05161f
C1103 dvdd_ip.n38 dvss 0.258748f
C1104 dvdd_ip.t47 dvss 0.05248f
C1105 dvdd_ip.t51 dvss 0.05251f
C1106 dvdd_ip.t37 dvss 0.05251f
C1107 dvdd_ip.n39 dvss 0.227267f
C1108 dvdd_ip.t35 dvss 0.05251f
C1109 dvdd_ip.t45 dvss 0.05251f
C1110 dvdd_ip.t43 dvss 0.05161f
C1111 dvdd_ip.n40 dvss 0.281525f
C1112 dvdd_ip.t44 dvss 0.05161f
C1113 dvdd_ip.n41 dvss 0.264717f
C1114 dvdd_ip.t48 dvss 0.052501f
C1115 dvdd_ip.t52 dvss 0.052518f
C1116 dvdd_ip.t28 dvss 0.052501f
C1117 dvdd_ip.n42 dvss 0.331183f
C1118 dvdd_ip.n43 dvss 0.234525f
C1119 dvdd_ip.n44 dvss 0.234525f
C1120 dvdd_ip.n45 dvss 0.7519f
C1121 dvdd_ip.t7 dvss 0.013318f
C1122 dvdd_ip.n47 dvss 0.773381f
C1123 dvdd_ip.n48 dvss 0.773381f
C1124 dvdd_ip.t13 dvss 0.013318f
C1125 dvdd_ip.n49 dvss 0.076958f
C1126 dvdd_ip.n50 dvss 0.058601f
C1127 dvdd_ip.n51 dvss 0.058601f
C1128 dvdd_ip.n52 dvss 0.538522f
C1129 dvdd_ip.n53 dvss 0.818296f
C1130 dvdd_ip.t21 dvss 0.013323f
C1131 dvdd_ip.n54 dvss 0.162119f
C1132 dvdd_ip.n55 dvss 0.097837f
C1133 dvdd_ip.n57 dvss 0.097837f
C1134 dvdd_ip.n58 dvss 0.088173f
C1135 dvdd_ip.n59 dvss 0.832248f
C1136 dvdd_ip.t20 dvss 1.16439f
C1137 dvdd_ip.n61 dvss 0.097837f
C1138 dvdd_ip.n62 dvss 0.832248f
C1139 dvdd_ip.n63 dvss 0.105489f
C1140 dvdd_ip.n64 dvss 0.635974f
C1141 dvdd_ip.t11 dvss 0.02854f
C1142 dvdd_ip.t16 dvss 0.02854f
C1143 dvdd_ip.n65 dvss 0.068444f
C1144 dvdd_ip.t53 dvss 0.02854f
C1145 dvdd_ip.t55 dvss 0.02854f
C1146 dvdd_ip.n66 dvss 0.068465f
C1147 dvdd_ip.t8 dvss 0.02854f
C1148 dvdd_ip.t54 dvss 0.02854f
C1149 dvdd_ip.n67 dvss 0.068444f
C1150 dvdd_ip.t14 dvss 0.02854f
C1151 dvdd_ip.t19 dvss 0.02854f
C1152 dvdd_ip.n68 dvss 0.068444f
C1153 dvdd_ip.t15 dvss 0.02854f
C1154 dvdd_ip.t18 dvss 0.02854f
C1155 dvdd_ip.n69 dvss 0.068465f
C1156 dvdd_ip.n70 dvss 2.09697f
C1157 dvdd_ip.n71 dvss 1.7395f
C1158 dvdd_ip.t1 dvss 0.104024f
C1159 dvdd_ip.n72 dvss 0.688131f
C1160 dvdd_ip.n73 dvss 0.067064f
C1161 dvdd_ip.t0 dvss 0.862706f
C1162 dvdd_ip.n76 dvss 0.067064f
C1163 dvdd_ip.n77 dvss 0.553603f
C1164 dvdd_ip.n80 dvss 0.503725f
C1165 dvdd_ip.n81 dvss 0.299443f
C1166 dvdd_ip.n82 dvss 0.361199f
C1167 dvdd_ip.t2 dvss 0.377055f
C1168 dvdd_ip.n83 dvss 0.243117f
C1169 dvdd_ip.t4 dvss 0.377055f
C1170 dvdd_ip.n84 dvss 0.361199f
C1171 dvdd_ip.n85 dvss 0.033188f
C1172 dvdd_ip.n86 dvss 0.3512f
C1173 dvdd_ip.n87 dvss 0.241382f
C1174 dvdd_ip.n88 dvss 0.105556f
C1175 dvdd_ip.n89 dvss 0.671287f
C1176 dvdd_ip.n90 dvss 0.509632f
C1177 dvdd_ip.n91 dvss 0.096026f
C1178 dvdd_ip.t6 dvss 1.28574f
C1179 dvdd_ip.n94 dvss 0.499573f
C1180 dvdd_ip.n95 dvss 0.307876f
C1181 dvdd_ip.n96 dvss 1.14024f
C1182 dvdd_ip.t22 dvss 1.45294f
C1183 dvdd_ip.t9 dvss 1.17811f
C1184 dvdd_ip.n97 dvss 0.785408f
C1185 dvdd_ip.t23 dvss 1.17811f
C1186 dvdd_ip.t10 dvss 1.45294f
C1187 dvdd_ip.n98 dvss 1.14024f
C1188 dvdd_ip.n99 dvss 0.044176f
C1189 dvdd_ip.n100 dvss 0.584225f
C1190 dvdd_ip.n101 dvss 0.833014f
C1191 dvdd_ip.n102 dvss 0.275953f
C1192 dvdd_ip.n103 dvss 0.969324f
C1193 dvdd_ip.t24 dvss 1.57246f
C1194 dvdd_ip.t40 dvss 1.9224f
C1195 dvdd_ip.t34 dvss 1.9224f
C1196 dvdd_ip.t36 dvss 1.4418f
C1197 dvdd_ip.n104 dvss 0.9612f
C1198 dvdd_ip.t42 dvss 1.4418f
C1199 dvdd_ip.t27 dvss 1.9224f
C1200 dvdd_ip.t38 dvss 1.9224f
C1201 dvdd_ip.t29 dvss 1.57246f
C1202 dvdd_ip.n105 dvss 0.969324f
C1203 vbp.n0 dvss 8.12052f
C1204 vbp.n1 dvss 0.149433f
C1205 vbp.n2 dvss 0.278043f
C1206 vbp.n3 dvss 0.309746f
C1207 vbp.t13 dvss 0.703868f
C1208 vbp.t12 dvss 0.614226f
C1209 vbp.n5 dvss 0.650619f
C1210 vbp.t5 dvss 0.752574f
C1211 vbp.n6 dvss 0.61948f
C1212 vbp.t2 dvss 0.090599f
C1213 vbp.t4 dvss 0.595378f
C1214 vbp.t7 dvss 0.595378f
C1215 vbp.n7 dvss 0.456086f
C1216 vbp.t17 dvss 0.608214f
C1217 vbp.n8 dvss 0.470076f
C1218 vbp.t11 dvss 0.705712f
C1219 vbp.n9 dvss 0.456086f
C1220 vbp.t14 dvss 0.595378f
C1221 vbp.t15 dvss 0.881413f
C1222 vbp.t8 dvss 0.683861f
C1223 vbp.t16 dvss 0.70411f
C1224 vbp.t6 dvss 0.724452f
C1225 vbp.t10 dvss 0.595378f
C1226 vbp.n10 dvss 0.456086f
C1227 vbp.t3 dvss 0.595378f
C1228 vbp.t1 dvss 0.64127f
C1229 vbp.t9 dvss 0.595378f
C1230 vbp.n11 dvss 0.456086f
C1231 vbp.t0 dvss 0.098789f
C1232 vbreg.n0 dvss 1.81217f
C1233 vbreg.n1 dvss 0.851099f
C1234 vbreg.n2 dvss 0.467546f
C1235 vbreg.n3 dvss 1.15478f
C1236 vbreg.n4 dvss 4.16667f
C1237 vbreg.n5 dvss 0.97222f
C1238 vbreg.n6 dvss 0.496926f
C1239 vbreg.n7 dvss 8.82024f
C1240 vbreg.n8 dvss 1.1584f
C1241 vbreg.n9 dvss 0.155057f
C1242 vbreg.n11 dvss 1.01043f
C1243 vbreg.n12 dvss 1.04968f
C1244 vbreg.n13 dvss 0.794925f
C1245 vbreg.n15 dvss 0.514068f
C1246 vbreg.n16 dvss 0.746492f
C1247 vbreg.n17 dvss 0.747813f
C1248 vbreg.n18 dvss 0.323996f
C1249 vbreg.n19 dvss 0.747813f
C1250 vbreg.t11 dvss 0.962705f
C1251 vbreg.n20 dvss 0.746492f
C1252 vbreg.n21 dvss 0.643449f
C1253 vbreg.n22 dvss 0.643449f
C1254 vbreg.n23 dvss 2.31728f
C1255 vbreg.n24 dvss 0.57718f
C1256 vbreg.n25 dvss 2.33154f
C1257 vbreg.n26 dvss 0.980351f
C1258 vbreg.t6 dvss 0.962705f
C1259 vbreg.n27 dvss 0.463288f
C1260 vbreg.t19 dvss 0.962705f
C1261 vbreg.n28 dvss 0.323996f
C1262 vbreg.n29 dvss 0.321619f
C1263 vbreg.t20 dvss 0.962705f
C1264 vbreg.t18 dvss 0.962705f
C1265 vbreg.t15 dvss 0.962705f
C1266 vbreg.n30 dvss 0.801483f
C1267 vbreg.t16 dvss 0.962705f
C1268 vbreg.n31 dvss 0.549792f
C1269 vbreg.n32 dvss 0.533473f
C1270 vbreg.n33 dvss 0.425139f
C1271 vbreg.n34 dvss 0.323996f
C1272 vbreg.t10 dvss 0.962705f
C1273 vbreg.t13 dvss 0.962705f
C1274 vbreg.n35 dvss 0.801483f
C1275 vbreg.n36 dvss 0.06842f
C1276 vbreg.n37 dvss 0.48842f
C1277 vbreg.t12 dvss 0.962705f
C1278 vbreg.n38 dvss 0.801483f
C1279 vbreg.t14 dvss 0.962705f
C1280 vbreg.n39 dvss 0.462848f
C1281 vbreg.n40 dvss 0.801483f
C1282 vbreg.t9 dvss 0.962705f
C1283 vbreg.n41 dvss 0.425139f
C1284 vbreg.n42 dvss 0.57343f
C1285 vbreg.t17 dvss 0.962705f
C1286 vbreg.n43 dvss 0.801483f
C1287 vbreg.n44 dvss 0.137064f
C1288 vbreg.n45 dvss 0.801483f
C1289 vbreg.t7 dvss 0.18306f
C1290 vbreg.n46 dvss 0.57105f
C1291 vbreg.n47 dvss 0.423817f
C1292 vbreg.n48 dvss 0.323996f
C1293 vbreg.n49 dvss 0.801483f
C1294 vbreg.t22 dvss 0.962705f
C1295 vbreg.n50 dvss 0.467693f
C1296 vbreg.t24 dvss 0.962705f
C1297 vbreg.t25 dvss 0.962705f
C1298 vbreg.n51 dvss 0.801483f
C1299 vbreg.t21 dvss 0.962705f
C1300 vbreg.n52 dvss 0.42602f
C1301 vbreg.n53 dvss 0.487245f
C1302 vbreg.t23 dvss 0.962705f
C1303 vbreg.n54 dvss 0.801483f
C1304 vbreg.n55 dvss 0.06886f
C1305 vbreg.n56 dvss 0.57483f
C1306 vbreg.n57 dvss 0.42602f
C1307 vbreg.n58 dvss 0.323996f
C1308 vbreg.n59 dvss 0.422936f
C1309 vbreg.n60 dvss 0.422936f
C1310 vbreg.n61 dvss 0.323996f
C1311 vbreg.n62 dvss 0.660032f
C1312 vbreg.t8 dvss 0.170945f
C1313 vbreg.t5 dvss 0.175683f
C1314 vbreg.t1 dvss 0.180252f
C1315 vbreg.t3 dvss 0.217084f
C1316 vbreg.t4 dvss 0.175417f
C1317 vbreg.t0 dvss 0.113684f
C1318 vbreg.t2 dvss 0.191737f
C1319 icnode.t1 dvss 0.024737f
C1320 icnode.t3 dvss 0.809758f
C1321 icnode.n0 dvss 3.30319f
C1322 icnode.t2 dvss 1.1318f
C1323 icnode.n1 dvss 1.04269f
C1324 icnode.n2 dvss 1.26325f
C1325 icnode.t0 dvss 39.8957f
C1326 icnode.n3 dvss 0.021984f
C1327 ena_ip.n0 dvss 0.816565f
C1328 ena_ip.n1 dvss 0.052729f
C1329 ena_ip.t1 dvss 0.038646f
C1330 ena_ip.n2 dvss 0.299073f
C1331 ena_ip.t14 dvss 0.312422f
C1332 ena_ip.t17 dvss 0.312179f
C1333 ena_ip.n3 dvss 0.262394f
C1334 ena_ip.n4 dvss 1.2068f
C1335 ena_ip.t2 dvss 0.357117f
C1336 ena_ip.t12 dvss 0.343909f
C1337 ena_ip.t18 dvss 0.013233f
C1338 ena_ip.t16 dvss 0.021012f
C1339 ena_ip.n5 dvss 0.040986f
C1340 ena_ip.t15 dvss 0.010303f
C1341 ena_ip.t4 dvss 0.024139f
C1342 ena_ip.n8 dvss 0.042815f
C1343 ena_ip.t10 dvss 0.013233f
C1344 ena_ip.t8 dvss 0.021012f
C1345 ena_ip.n9 dvss 0.040986f
C1346 ena_ip.t5 dvss 0.010303f
C1347 ena_ip.t13 dvss 0.024139f
C1348 ena_ip.n12 dvss 0.042815f
C1349 ena_ip.t9 dvss 0.013233f
C1350 ena_ip.t6 dvss 0.021012f
C1351 ena_ip.n13 dvss 0.040986f
C1352 ena_ip.t3 dvss 0.010303f
C1353 ena_ip.t7 dvss 0.024139f
C1354 ena_ip.n16 dvss 0.042815f
C1355 ena_ip.t19 dvss 0.025235f
C1356 ena_ip.t11 dvss 0.015832f
C1357 ena_ip.n17 dvss 0.036079f
C1358 ena_ip.n18 dvss 0.024525f
C1359 ena_ip.n19 dvss 0.153572f
C1360 ena_ip.t0 dvss 0.026873f
C1361 dvdd.t126 dvss 0.010255f
C1362 dvdd.t114 dvss 0.010255f
C1363 dvdd.n0 dvss 0.232741f
C1364 dvdd.n1 dvss 0.072395f
C1365 dvdd.n3 dvss 0.016649f
C1366 dvdd.n4 dvss 0.115384f
C1367 dvdd.n5 dvss 0.115384f
C1368 dvdd.t41 dvss 0.054374f
C1369 dvdd.t147 dvss 0.018382f
C1370 dvdd.n9 dvss 0.013708f
C1371 dvdd.n11 dvss 0.045003f
C1372 dvdd.n14 dvss 0.023574f
C1373 dvdd.n15 dvss 0.028089f
C1374 dvdd.n16 dvss 0.018614f
C1375 dvdd.t137 dvss 0.054374f
C1376 dvdd.t32 dvss 0.018382f
C1377 dvdd.n18 dvss 0.045003f
C1378 dvdd.n23 dvss 0.013708f
C1379 dvdd.n25 dvss 0.028989f
C1380 dvdd.n26 dvss 0.0118f
C1381 dvdd.n27 dvss 0.115384f
C1382 dvdd.n28 dvss 0.016649f
C1383 dvdd.n29 dvss 0.115384f
C1384 dvdd.n30 dvss 0.016663f
C1385 dvdd.t113 dvss 0.166037f
C1386 dvdd.n33 dvss 0.016663f
C1387 dvdd.n34 dvss 0.0118f
C1388 dvdd.n38 dvss 0.47509f
C1389 dvdd.n39 dvss 0.250837f
C1390 dvdd.n41 dvss 0.0118f
C1391 dvdd.n42 dvss 0.016663f
C1392 dvdd.t125 dvss 0.166037f
C1393 dvdd.n45 dvss 0.016663f
C1394 dvdd.n46 dvss 0.0118f
C1395 dvdd.n48 dvss 0.098284f
C1396 dvdd.n49 dvss 1.85368f
C1397 dvdd.t175 dvss 3.84974f
C1398 dvdd.n50 dvss 3.24063f
C1399 dvdd.n51 dvss 1.77951f
C1400 dvdd.n53 dvss 0.032035f
C1401 dvdd.n54 dvss 0.032035f
C1402 dvdd.n55 dvss 0.032035f
C1403 dvdd.n56 dvss 0.013403f
C1404 dvdd.n57 dvss 0.011326f
C1405 dvdd.n67 dvss 0.018622f
C1406 dvdd.n71 dvss 0.012463f
C1407 dvdd.n88 dvss 0.018622f
C1408 dvdd.n92 dvss 0.012463f
C1409 dvdd.n109 dvss 0.018622f
C1410 dvdd.n113 dvss 0.012463f
C1411 dvdd.n123 dvss 0.015374f
C1412 dvdd.n129 dvss 0.026036f
C1413 dvdd.n142 dvss 0.013299f
C1414 dvdd.n149 dvss 0.013074f
C1415 dvdd.n154 dvss 0.016521f
C1416 dvdd.n161 dvss 0.015374f
C1417 dvdd.n167 dvss 0.026036f
C1418 dvdd.n180 dvss 0.013299f
C1419 dvdd.n187 dvss 0.013074f
C1420 dvdd.n192 dvss 0.016521f
C1421 dvdd.n199 dvss 0.015374f
C1422 dvdd.n205 dvss 0.026036f
C1423 dvdd.n218 dvss 0.013299f
C1424 dvdd.n225 dvss 0.013074f
C1425 dvdd.n230 dvss 0.016521f
C1426 dvdd.n238 dvss 0.037612f
C1427 dvdd.n240 dvss 0.011337f
C1428 dvdd.t62 dvss 0.05252f
C1429 dvdd.t37 dvss 0.027032f
C1430 dvdd.t39 dvss 0.021162f
C1431 dvdd.t130 dvss 0.039081f
C1432 dvdd.t10 dvss 0.029194f
C1433 dvdd.t141 dvss 0.04387f
C1434 dvdd.t158 dvss 0.042016f
C1435 dvdd.t98 dvss 0.025951f
C1436 dvdd.t19 dvss 0.01761f
C1437 dvdd.n245 dvss 0.045201f
C1438 dvdd.n246 dvss 0.046181f
C1439 dvdd.n254 dvss 0.010815f
C1440 dvdd.n257 dvss 0.013065f
C1441 dvdd.n265 dvss 0.013257f
C1442 dvdd.n267 dvss 0.032892f
C1443 dvdd.n269 dvss 0.071148f
C1444 dvdd.t52 dvss 0.045486f
C1445 dvdd.t12 dvss 0.065913f
C1446 dvdd.t82 dvss 0.084434f
C1447 dvdd.n270 dvss 0.072307f
C1448 dvdd.t28 dvss 0.040583f
C1449 dvdd.t24 dvss 0.095601f
C1450 dvdd.t123 dvss 0.09778f
C1451 dvdd.t136 dvss 0.052023f
C1452 dvdd.t89 dvss 0.065096f
C1453 dvdd.t43 dvss 0.064551f
C1454 dvdd.t91 dvss 0.080077f
C1455 dvdd.t121 dvss 0.080621f
C1456 dvdd.t104 dvss 0.050388f
C1457 dvdd.t26 dvss 0.046303f
C1458 dvdd.t58 dvss 0.052295f
C1459 dvdd.t65 dvss 0.052295f
C1460 dvdd.t8 dvss 0.067548f
C1461 dvdd.t101 dvss 0.104317f
C1462 dvdd.t2 dvss 0.086069f
C1463 dvdd.t4 dvss 0.067548f
C1464 dvdd.n271 dvss 0.070945f
C1465 dvdd.t46 dvss 0.040583f
C1466 dvdd.t20 dvss 0.095601f
C1467 dvdd.t68 dvss 0.09778f
C1468 dvdd.t18 dvss 0.052023f
C1469 dvdd.t36 dvss 0.065096f
C1470 dvdd.t60 dvss 0.064551f
C1471 dvdd.t111 dvss 0.080077f
C1472 dvdd.t79 dvss 0.080621f
C1473 dvdd.t34 dvss 0.050388f
C1474 dvdd.t45 dvss 0.046303f
C1475 dvdd.t86 dvss 0.052295f
C1476 dvdd.t94 dvss 0.052295f
C1477 dvdd.t63 dvss 0.067548f
C1478 dvdd.t84 dvss 0.104317f
C1479 dvdd.t48 dvss 0.086069f
C1480 dvdd.t108 dvss 0.067548f
C1481 dvdd.n272 dvss 0.070945f
C1482 dvdd.t119 dvss 0.040583f
C1483 dvdd.t145 dvss 0.095601f
C1484 dvdd.t14 dvss 0.09778f
C1485 dvdd.t105 dvss 0.052023f
C1486 dvdd.t103 dvss 0.065096f
C1487 dvdd.t0 dvss 0.064551f
C1488 dvdd.t134 dvss 0.080077f
C1489 dvdd.t6 dvss 0.080621f
C1490 dvdd.t144 dvss 0.050388f
C1491 dvdd.t106 dvss 0.046303f
C1492 dvdd.t54 dvss 0.052295f
C1493 dvdd.t30 dvss 0.052295f
C1494 dvdd.t50 dvss 0.067548f
C1495 dvdd.t56 dvss 0.104317f
C1496 dvdd.t132 dvss 0.086069f
C1497 dvdd.t16 dvss 0.096045f
C1498 dvdd.n273 dvss 0.098227f
C1499 dvdd.n274 dvss 2.52168f
C1500 dvdd.n275 dvss 12.367001f
C1501 dvdd.t178 dvss 3.84974f
C1502 dvdd.n276 dvss 6.82163f
C1503 dvdd.t177 dvss 3.84974f
C1504 dvdd.n277 dvss 3.74301f
C1505 dvdd.t176 dvss 3.84974f
C1506 dvdd.n278 dvss 3.62059f
C1507 dvdd.n279 dvss 2.58506f
C1508 dvdd.n280 dvss 0.391933f
C1509 dvdd.t167 dvss 0.011164f
C1510 dvdd.t74 dvss 0.011164f
C1511 dvdd.n281 dvss 0.026774f
C1512 dvdd.t116 dvss 0.011164f
C1513 dvdd.t23 dvss 0.011164f
C1514 dvdd.n282 dvss 0.026774f
C1515 dvdd.n283 dvss 0.052444f
C1516 dvdd.t165 dvss 0.040692f
C1517 dvdd.n284 dvss 0.048107f
C1518 dvdd.n285 dvss 0.047967f
C1519 dvdd.n286 dvss 0.047967f
C1520 dvdd.t71 dvss 0.040692f
C1521 dvdd.t78 dvss 0.011164f
C1522 dvdd.t76 dvss 0.011164f
C1523 dvdd.n287 dvss 0.026774f
C1524 dvdd.t97 dvss 0.011164f
C1525 dvdd.t162 dvss 0.011164f
C1526 dvdd.n288 dvss 0.026774f
C1527 dvdd.n289 dvss 0.467698f
C1528 dvdd.n290 dvss 0.872117f
C1529 dvdd.n291 dvss 0.243934f
C1530 dvdd.n292 dvss 0.211775f
C1531 dvdd.t70 dvss 0.223699f
C1532 dvdd.t77 dvss 0.188256f
C1533 dvdd.t75 dvss 0.188256f
C1534 dvdd.t96 dvss 0.188256f
C1535 dvdd.t161 dvss 0.141192f
C1536 dvdd.n293 dvss 0.094128f
C1537 dvdd.t166 dvss 0.141192f
C1538 dvdd.t73 dvss 0.188256f
C1539 dvdd.t115 dvss 0.188256f
C1540 dvdd.t22 dvss 0.188256f
C1541 dvdd.t164 dvss 0.223699f
C1542 dvdd.n294 dvss 0.211775f
C1543 dvdd.n295 dvss 0.256858f
C1544 dvdd.n296 dvss 0.776554f
C1545 dvdd.n297 dvss 0.376011f
C1546 dvdd.n298 dvss 0.088779f
C1547 x7.x3.A2.t1 dvss 0.057884f
C1548 x7.x3.A2.t5 dvss 0.028593f
C1549 x7.x3.A2.t7 dvss 0.017955f
C1550 x7.x3.A2.n0 dvss 0.038437f
C1551 x7.x3.A2.n1 dvss 0.153155f
C1552 x7.x3.A2.t4 dvss 0.015834f
C1553 x7.x3.A2.n2 dvss 0.048959f
C1554 x7.x3.A2.t3 dvss 0.015657f
C1555 x7.x3.A2.n3 dvss 0.044896f
C1556 x7.x3.A2.n4 dvss 0.047435f
C1557 x7.x3.A2.t2 dvss 0.02131f
C1558 x7.x3.A2.t6 dvss 0.023458f
C1559 x7.x3.A2.n5 dvss 0.067085f
C1560 x7.x3.A2.n6 dvss 1.6639f
C1561 x7.x3.A2.n7 dvss 0.069954f
C1562 x7.x3.A2.t0 dvss 0.043534f
.ends

