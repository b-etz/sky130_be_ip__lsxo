magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< metal4 >>
rect -7545 7039 -4847 7080
rect -7545 4961 -5103 7039
rect -4867 4961 -4847 7039
rect -7545 4920 -4847 4961
rect -4447 7039 -1749 7080
rect -4447 4961 -2005 7039
rect -1769 4961 -1749 7039
rect -4447 4920 -1749 4961
rect -1349 7039 1349 7080
rect -1349 4961 1093 7039
rect 1329 4961 1349 7039
rect -1349 4920 1349 4961
rect 1749 7039 4447 7080
rect 1749 4961 4191 7039
rect 4427 4961 4447 7039
rect 1749 4920 4447 4961
rect 4847 7039 7545 7080
rect 4847 4961 7289 7039
rect 7525 4961 7545 7039
rect 4847 4920 7545 4961
rect -7545 4639 -4847 4680
rect -7545 2561 -5103 4639
rect -4867 2561 -4847 4639
rect -7545 2520 -4847 2561
rect -4447 4639 -1749 4680
rect -4447 2561 -2005 4639
rect -1769 2561 -1749 4639
rect -4447 2520 -1749 2561
rect -1349 4639 1349 4680
rect -1349 2561 1093 4639
rect 1329 2561 1349 4639
rect -1349 2520 1349 2561
rect 1749 4639 4447 4680
rect 1749 2561 4191 4639
rect 4427 2561 4447 4639
rect 1749 2520 4447 2561
rect 4847 4639 7545 4680
rect 4847 2561 7289 4639
rect 7525 2561 7545 4639
rect 4847 2520 7545 2561
rect -7545 2239 -4847 2280
rect -7545 161 -5103 2239
rect -4867 161 -4847 2239
rect -7545 120 -4847 161
rect -4447 2239 -1749 2280
rect -4447 161 -2005 2239
rect -1769 161 -1749 2239
rect -4447 120 -1749 161
rect -1349 2239 1349 2280
rect -1349 161 1093 2239
rect 1329 161 1349 2239
rect -1349 120 1349 161
rect 1749 2239 4447 2280
rect 1749 161 4191 2239
rect 4427 161 4447 2239
rect 1749 120 4447 161
rect 4847 2239 7545 2280
rect 4847 161 7289 2239
rect 7525 161 7545 2239
rect 4847 120 7545 161
rect -7545 -161 -4847 -120
rect -7545 -2239 -5103 -161
rect -4867 -2239 -4847 -161
rect -7545 -2280 -4847 -2239
rect -4447 -161 -1749 -120
rect -4447 -2239 -2005 -161
rect -1769 -2239 -1749 -161
rect -4447 -2280 -1749 -2239
rect -1349 -161 1349 -120
rect -1349 -2239 1093 -161
rect 1329 -2239 1349 -161
rect -1349 -2280 1349 -2239
rect 1749 -161 4447 -120
rect 1749 -2239 4191 -161
rect 4427 -2239 4447 -161
rect 1749 -2280 4447 -2239
rect 4847 -161 7545 -120
rect 4847 -2239 7289 -161
rect 7525 -2239 7545 -161
rect 4847 -2280 7545 -2239
rect -7545 -2561 -4847 -2520
rect -7545 -4639 -5103 -2561
rect -4867 -4639 -4847 -2561
rect -7545 -4680 -4847 -4639
rect -4447 -2561 -1749 -2520
rect -4447 -4639 -2005 -2561
rect -1769 -4639 -1749 -2561
rect -4447 -4680 -1749 -4639
rect -1349 -2561 1349 -2520
rect -1349 -4639 1093 -2561
rect 1329 -4639 1349 -2561
rect -1349 -4680 1349 -4639
rect 1749 -2561 4447 -2520
rect 1749 -4639 4191 -2561
rect 4427 -4639 4447 -2561
rect 1749 -4680 4447 -4639
rect 4847 -2561 7545 -2520
rect 4847 -4639 7289 -2561
rect 7525 -4639 7545 -2561
rect 4847 -4680 7545 -4639
rect -7545 -4961 -4847 -4920
rect -7545 -7039 -5103 -4961
rect -4867 -7039 -4847 -4961
rect -7545 -7080 -4847 -7039
rect -4447 -4961 -1749 -4920
rect -4447 -7039 -2005 -4961
rect -1769 -7039 -1749 -4961
rect -4447 -7080 -1749 -7039
rect -1349 -4961 1349 -4920
rect -1349 -7039 1093 -4961
rect 1329 -7039 1349 -4961
rect -1349 -7080 1349 -7039
rect 1749 -4961 4447 -4920
rect 1749 -7039 4191 -4961
rect 4427 -7039 4447 -4961
rect 1749 -7080 4447 -7039
rect 4847 -4961 7545 -4920
rect 4847 -7039 7289 -4961
rect 7525 -7039 7545 -4961
rect 4847 -7080 7545 -7039
<< via4 >>
rect -5103 4961 -4867 7039
rect -2005 4961 -1769 7039
rect 1093 4961 1329 7039
rect 4191 4961 4427 7039
rect 7289 4961 7525 7039
rect -5103 2561 -4867 4639
rect -2005 2561 -1769 4639
rect 1093 2561 1329 4639
rect 4191 2561 4427 4639
rect 7289 2561 7525 4639
rect -5103 161 -4867 2239
rect -2005 161 -1769 2239
rect 1093 161 1329 2239
rect 4191 161 4427 2239
rect 7289 161 7525 2239
rect -5103 -2239 -4867 -161
rect -2005 -2239 -1769 -161
rect 1093 -2239 1329 -161
rect 4191 -2239 4427 -161
rect 7289 -2239 7525 -161
rect -5103 -4639 -4867 -2561
rect -2005 -4639 -1769 -2561
rect 1093 -4639 1329 -2561
rect 4191 -4639 4427 -2561
rect 7289 -4639 7525 -2561
rect -5103 -7039 -4867 -4961
rect -2005 -7039 -1769 -4961
rect 1093 -7039 1329 -4961
rect 4191 -7039 4427 -4961
rect 7289 -7039 7525 -4961
<< mimcap2 >>
rect -7465 6960 -5465 7000
rect -7465 5040 -7425 6960
rect -5505 5040 -5465 6960
rect -7465 5000 -5465 5040
rect -4367 6960 -2367 7000
rect -4367 5040 -4327 6960
rect -2407 5040 -2367 6960
rect -4367 5000 -2367 5040
rect -1269 6960 731 7000
rect -1269 5040 -1229 6960
rect 691 5040 731 6960
rect -1269 5000 731 5040
rect 1829 6960 3829 7000
rect 1829 5040 1869 6960
rect 3789 5040 3829 6960
rect 1829 5000 3829 5040
rect 4927 6960 6927 7000
rect 4927 5040 4967 6960
rect 6887 5040 6927 6960
rect 4927 5000 6927 5040
rect -7465 4560 -5465 4600
rect -7465 2640 -7425 4560
rect -5505 2640 -5465 4560
rect -7465 2600 -5465 2640
rect -4367 4560 -2367 4600
rect -4367 2640 -4327 4560
rect -2407 2640 -2367 4560
rect -4367 2600 -2367 2640
rect -1269 4560 731 4600
rect -1269 2640 -1229 4560
rect 691 2640 731 4560
rect -1269 2600 731 2640
rect 1829 4560 3829 4600
rect 1829 2640 1869 4560
rect 3789 2640 3829 4560
rect 1829 2600 3829 2640
rect 4927 4560 6927 4600
rect 4927 2640 4967 4560
rect 6887 2640 6927 4560
rect 4927 2600 6927 2640
rect -7465 2160 -5465 2200
rect -7465 240 -7425 2160
rect -5505 240 -5465 2160
rect -7465 200 -5465 240
rect -4367 2160 -2367 2200
rect -4367 240 -4327 2160
rect -2407 240 -2367 2160
rect -4367 200 -2367 240
rect -1269 2160 731 2200
rect -1269 240 -1229 2160
rect 691 240 731 2160
rect -1269 200 731 240
rect 1829 2160 3829 2200
rect 1829 240 1869 2160
rect 3789 240 3829 2160
rect 1829 200 3829 240
rect 4927 2160 6927 2200
rect 4927 240 4967 2160
rect 6887 240 6927 2160
rect 4927 200 6927 240
rect -7465 -240 -5465 -200
rect -7465 -2160 -7425 -240
rect -5505 -2160 -5465 -240
rect -7465 -2200 -5465 -2160
rect -4367 -240 -2367 -200
rect -4367 -2160 -4327 -240
rect -2407 -2160 -2367 -240
rect -4367 -2200 -2367 -2160
rect -1269 -240 731 -200
rect -1269 -2160 -1229 -240
rect 691 -2160 731 -240
rect -1269 -2200 731 -2160
rect 1829 -240 3829 -200
rect 1829 -2160 1869 -240
rect 3789 -2160 3829 -240
rect 1829 -2200 3829 -2160
rect 4927 -240 6927 -200
rect 4927 -2160 4967 -240
rect 6887 -2160 6927 -240
rect 4927 -2200 6927 -2160
rect -7465 -2640 -5465 -2600
rect -7465 -4560 -7425 -2640
rect -5505 -4560 -5465 -2640
rect -7465 -4600 -5465 -4560
rect -4367 -2640 -2367 -2600
rect -4367 -4560 -4327 -2640
rect -2407 -4560 -2367 -2640
rect -4367 -4600 -2367 -4560
rect -1269 -2640 731 -2600
rect -1269 -4560 -1229 -2640
rect 691 -4560 731 -2640
rect -1269 -4600 731 -4560
rect 1829 -2640 3829 -2600
rect 1829 -4560 1869 -2640
rect 3789 -4560 3829 -2640
rect 1829 -4600 3829 -4560
rect 4927 -2640 6927 -2600
rect 4927 -4560 4967 -2640
rect 6887 -4560 6927 -2640
rect 4927 -4600 6927 -4560
rect -7465 -5040 -5465 -5000
rect -7465 -6960 -7425 -5040
rect -5505 -6960 -5465 -5040
rect -7465 -7000 -5465 -6960
rect -4367 -5040 -2367 -5000
rect -4367 -6960 -4327 -5040
rect -2407 -6960 -2367 -5040
rect -4367 -7000 -2367 -6960
rect -1269 -5040 731 -5000
rect -1269 -6960 -1229 -5040
rect 691 -6960 731 -5040
rect -1269 -7000 731 -6960
rect 1829 -5040 3829 -5000
rect 1829 -6960 1869 -5040
rect 3789 -6960 3829 -5040
rect 1829 -7000 3829 -6960
rect 4927 -5040 6927 -5000
rect 4927 -6960 4967 -5040
rect 6887 -6960 6927 -5040
rect 4927 -7000 6927 -6960
<< mimcap2contact >>
rect -7425 5040 -5505 6960
rect -4327 5040 -2407 6960
rect -1229 5040 691 6960
rect 1869 5040 3789 6960
rect 4967 5040 6887 6960
rect -7425 2640 -5505 4560
rect -4327 2640 -2407 4560
rect -1229 2640 691 4560
rect 1869 2640 3789 4560
rect 4967 2640 6887 4560
rect -7425 240 -5505 2160
rect -4327 240 -2407 2160
rect -1229 240 691 2160
rect 1869 240 3789 2160
rect 4967 240 6887 2160
rect -7425 -2160 -5505 -240
rect -4327 -2160 -2407 -240
rect -1229 -2160 691 -240
rect 1869 -2160 3789 -240
rect 4967 -2160 6887 -240
rect -7425 -4560 -5505 -2640
rect -4327 -4560 -2407 -2640
rect -1229 -4560 691 -2640
rect 1869 -4560 3789 -2640
rect 4967 -4560 6887 -2640
rect -7425 -6960 -5505 -5040
rect -4327 -6960 -2407 -5040
rect -1229 -6960 691 -5040
rect 1869 -6960 3789 -5040
rect 4967 -6960 6887 -5040
<< metal5 >>
rect -6625 6984 -6305 7200
rect -5145 7039 -4825 7200
rect -7449 6960 -5481 6984
rect -7449 5040 -7425 6960
rect -5505 5040 -5481 6960
rect -7449 5016 -5481 5040
rect -6625 4584 -6305 5016
rect -5145 4961 -5103 7039
rect -4867 4961 -4825 7039
rect -3527 6984 -3207 7200
rect -2047 7039 -1727 7200
rect -4351 6960 -2383 6984
rect -4351 5040 -4327 6960
rect -2407 5040 -2383 6960
rect -4351 5016 -2383 5040
rect -5145 4639 -4825 4961
rect -7449 4560 -5481 4584
rect -7449 2640 -7425 4560
rect -5505 2640 -5481 4560
rect -7449 2616 -5481 2640
rect -6625 2184 -6305 2616
rect -5145 2561 -5103 4639
rect -4867 2561 -4825 4639
rect -3527 4584 -3207 5016
rect -2047 4961 -2005 7039
rect -1769 4961 -1727 7039
rect -429 6984 -109 7200
rect 1051 7039 1371 7200
rect -1253 6960 715 6984
rect -1253 5040 -1229 6960
rect 691 5040 715 6960
rect -1253 5016 715 5040
rect -2047 4639 -1727 4961
rect -4351 4560 -2383 4584
rect -4351 2640 -4327 4560
rect -2407 2640 -2383 4560
rect -4351 2616 -2383 2640
rect -5145 2239 -4825 2561
rect -7449 2160 -5481 2184
rect -7449 240 -7425 2160
rect -5505 240 -5481 2160
rect -7449 216 -5481 240
rect -6625 -216 -6305 216
rect -5145 161 -5103 2239
rect -4867 161 -4825 2239
rect -3527 2184 -3207 2616
rect -2047 2561 -2005 4639
rect -1769 2561 -1727 4639
rect -429 4584 -109 5016
rect 1051 4961 1093 7039
rect 1329 4961 1371 7039
rect 2669 6984 2989 7200
rect 4149 7039 4469 7200
rect 1845 6960 3813 6984
rect 1845 5040 1869 6960
rect 3789 5040 3813 6960
rect 1845 5016 3813 5040
rect 1051 4639 1371 4961
rect -1253 4560 715 4584
rect -1253 2640 -1229 4560
rect 691 2640 715 4560
rect -1253 2616 715 2640
rect -2047 2239 -1727 2561
rect -4351 2160 -2383 2184
rect -4351 240 -4327 2160
rect -2407 240 -2383 2160
rect -4351 216 -2383 240
rect -5145 -161 -4825 161
rect -7449 -240 -5481 -216
rect -7449 -2160 -7425 -240
rect -5505 -2160 -5481 -240
rect -7449 -2184 -5481 -2160
rect -6625 -2616 -6305 -2184
rect -5145 -2239 -5103 -161
rect -4867 -2239 -4825 -161
rect -3527 -216 -3207 216
rect -2047 161 -2005 2239
rect -1769 161 -1727 2239
rect -429 2184 -109 2616
rect 1051 2561 1093 4639
rect 1329 2561 1371 4639
rect 2669 4584 2989 5016
rect 4149 4961 4191 7039
rect 4427 4961 4469 7039
rect 5767 6984 6087 7200
rect 7247 7039 7567 7200
rect 4943 6960 6911 6984
rect 4943 5040 4967 6960
rect 6887 5040 6911 6960
rect 4943 5016 6911 5040
rect 4149 4639 4469 4961
rect 1845 4560 3813 4584
rect 1845 2640 1869 4560
rect 3789 2640 3813 4560
rect 1845 2616 3813 2640
rect 1051 2239 1371 2561
rect -1253 2160 715 2184
rect -1253 240 -1229 2160
rect 691 240 715 2160
rect -1253 216 715 240
rect -2047 -161 -1727 161
rect -4351 -240 -2383 -216
rect -4351 -2160 -4327 -240
rect -2407 -2160 -2383 -240
rect -4351 -2184 -2383 -2160
rect -5145 -2561 -4825 -2239
rect -7449 -2640 -5481 -2616
rect -7449 -4560 -7425 -2640
rect -5505 -4560 -5481 -2640
rect -7449 -4584 -5481 -4560
rect -6625 -5016 -6305 -4584
rect -5145 -4639 -5103 -2561
rect -4867 -4639 -4825 -2561
rect -3527 -2616 -3207 -2184
rect -2047 -2239 -2005 -161
rect -1769 -2239 -1727 -161
rect -429 -216 -109 216
rect 1051 161 1093 2239
rect 1329 161 1371 2239
rect 2669 2184 2989 2616
rect 4149 2561 4191 4639
rect 4427 2561 4469 4639
rect 5767 4584 6087 5016
rect 7247 4961 7289 7039
rect 7525 4961 7567 7039
rect 7247 4639 7567 4961
rect 4943 4560 6911 4584
rect 4943 2640 4967 4560
rect 6887 2640 6911 4560
rect 4943 2616 6911 2640
rect 4149 2239 4469 2561
rect 1845 2160 3813 2184
rect 1845 240 1869 2160
rect 3789 240 3813 2160
rect 1845 216 3813 240
rect 1051 -161 1371 161
rect -1253 -240 715 -216
rect -1253 -2160 -1229 -240
rect 691 -2160 715 -240
rect -1253 -2184 715 -2160
rect -2047 -2561 -1727 -2239
rect -4351 -2640 -2383 -2616
rect -4351 -4560 -4327 -2640
rect -2407 -4560 -2383 -2640
rect -4351 -4584 -2383 -4560
rect -5145 -4961 -4825 -4639
rect -7449 -5040 -5481 -5016
rect -7449 -6960 -7425 -5040
rect -5505 -6960 -5481 -5040
rect -7449 -6984 -5481 -6960
rect -6625 -7200 -6305 -6984
rect -5145 -7039 -5103 -4961
rect -4867 -7039 -4825 -4961
rect -3527 -5016 -3207 -4584
rect -2047 -4639 -2005 -2561
rect -1769 -4639 -1727 -2561
rect -429 -2616 -109 -2184
rect 1051 -2239 1093 -161
rect 1329 -2239 1371 -161
rect 2669 -216 2989 216
rect 4149 161 4191 2239
rect 4427 161 4469 2239
rect 5767 2184 6087 2616
rect 7247 2561 7289 4639
rect 7525 2561 7567 4639
rect 7247 2239 7567 2561
rect 4943 2160 6911 2184
rect 4943 240 4967 2160
rect 6887 240 6911 2160
rect 4943 216 6911 240
rect 4149 -161 4469 161
rect 1845 -240 3813 -216
rect 1845 -2160 1869 -240
rect 3789 -2160 3813 -240
rect 1845 -2184 3813 -2160
rect 1051 -2561 1371 -2239
rect -1253 -2640 715 -2616
rect -1253 -4560 -1229 -2640
rect 691 -4560 715 -2640
rect -1253 -4584 715 -4560
rect -2047 -4961 -1727 -4639
rect -4351 -5040 -2383 -5016
rect -4351 -6960 -4327 -5040
rect -2407 -6960 -2383 -5040
rect -4351 -6984 -2383 -6960
rect -5145 -7200 -4825 -7039
rect -3527 -7200 -3207 -6984
rect -2047 -7039 -2005 -4961
rect -1769 -7039 -1727 -4961
rect -429 -5016 -109 -4584
rect 1051 -4639 1093 -2561
rect 1329 -4639 1371 -2561
rect 2669 -2616 2989 -2184
rect 4149 -2239 4191 -161
rect 4427 -2239 4469 -161
rect 5767 -216 6087 216
rect 7247 161 7289 2239
rect 7525 161 7567 2239
rect 7247 -161 7567 161
rect 4943 -240 6911 -216
rect 4943 -2160 4967 -240
rect 6887 -2160 6911 -240
rect 4943 -2184 6911 -2160
rect 4149 -2561 4469 -2239
rect 1845 -2640 3813 -2616
rect 1845 -4560 1869 -2640
rect 3789 -4560 3813 -2640
rect 1845 -4584 3813 -4560
rect 1051 -4961 1371 -4639
rect -1253 -5040 715 -5016
rect -1253 -6960 -1229 -5040
rect 691 -6960 715 -5040
rect -1253 -6984 715 -6960
rect -2047 -7200 -1727 -7039
rect -429 -7200 -109 -6984
rect 1051 -7039 1093 -4961
rect 1329 -7039 1371 -4961
rect 2669 -5016 2989 -4584
rect 4149 -4639 4191 -2561
rect 4427 -4639 4469 -2561
rect 5767 -2616 6087 -2184
rect 7247 -2239 7289 -161
rect 7525 -2239 7567 -161
rect 7247 -2561 7567 -2239
rect 4943 -2640 6911 -2616
rect 4943 -4560 4967 -2640
rect 6887 -4560 6911 -2640
rect 4943 -4584 6911 -4560
rect 4149 -4961 4469 -4639
rect 1845 -5040 3813 -5016
rect 1845 -6960 1869 -5040
rect 3789 -6960 3813 -5040
rect 1845 -6984 3813 -6960
rect 1051 -7200 1371 -7039
rect 2669 -7200 2989 -6984
rect 4149 -7039 4191 -4961
rect 4427 -7039 4469 -4961
rect 5767 -5016 6087 -4584
rect 7247 -4639 7289 -2561
rect 7525 -4639 7567 -2561
rect 7247 -4961 7567 -4639
rect 4943 -5040 6911 -5016
rect 4943 -6960 4967 -5040
rect 6887 -6960 6911 -5040
rect 4943 -6984 6911 -6960
rect 4149 -7200 4469 -7039
rect 5767 -7200 6087 -6984
rect 7247 -7039 7289 -4961
rect 7525 -7039 7567 -4961
rect 7247 -7200 7567 -7039
<< properties >>
string FIXED_BBOX 4847 4920 7007 7080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 5 ny 6 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
