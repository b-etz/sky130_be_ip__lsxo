magic
tech sky130A
magscale 1 2
timestamp 1712888116
<< pwell >>
rect -2193 -11782 2193 11782
<< psubdiff >>
rect -2157 11712 -2061 11746
rect 2061 11712 2157 11746
rect -2157 11650 -2123 11712
rect 2123 11650 2157 11712
rect -2157 -11712 -2123 -11650
rect 2123 -11712 2157 -11650
rect -2157 -11746 -2061 -11712
rect 2061 -11746 2157 -11712
<< psubdiffcont >>
rect -2061 11712 2061 11746
rect -2157 -11650 -2123 11650
rect 2123 -11650 2157 11650
rect -2061 -11746 2061 -11712
<< xpolycontact >>
rect -2027 11184 -1957 11616
rect -2027 -11616 -1957 -11184
rect -1861 11184 -1791 11616
rect -1861 -11616 -1791 -11184
rect -1695 11184 -1625 11616
rect -1695 -11616 -1625 -11184
rect -1529 11184 -1459 11616
rect -1529 -11616 -1459 -11184
rect -1363 11184 -1293 11616
rect -1363 -11616 -1293 -11184
rect -1197 11184 -1127 11616
rect -1197 -11616 -1127 -11184
rect -1031 11184 -961 11616
rect -1031 -11616 -961 -11184
rect -865 11184 -795 11616
rect -865 -11616 -795 -11184
rect -699 11184 -629 11616
rect -699 -11616 -629 -11184
rect -533 11184 -463 11616
rect -533 -11616 -463 -11184
rect -367 11184 -297 11616
rect -367 -11616 -297 -11184
rect -201 11184 -131 11616
rect -201 -11616 -131 -11184
rect -35 11184 35 11616
rect -35 -11616 35 -11184
rect 131 11184 201 11616
rect 131 -11616 201 -11184
rect 297 11184 367 11616
rect 297 -11616 367 -11184
rect 463 11184 533 11616
rect 463 -11616 533 -11184
rect 629 11184 699 11616
rect 629 -11616 699 -11184
rect 795 11184 865 11616
rect 795 -11616 865 -11184
rect 961 11184 1031 11616
rect 961 -11616 1031 -11184
rect 1127 11184 1197 11616
rect 1127 -11616 1197 -11184
rect 1293 11184 1363 11616
rect 1293 -11616 1363 -11184
rect 1459 11184 1529 11616
rect 1459 -11616 1529 -11184
rect 1625 11184 1695 11616
rect 1625 -11616 1695 -11184
rect 1791 11184 1861 11616
rect 1791 -11616 1861 -11184
rect 1957 11184 2027 11616
rect 1957 -11616 2027 -11184
<< xpolyres >>
rect -2027 -11184 -1957 11184
rect -1861 -11184 -1791 11184
rect -1695 -11184 -1625 11184
rect -1529 -11184 -1459 11184
rect -1363 -11184 -1293 11184
rect -1197 -11184 -1127 11184
rect -1031 -11184 -961 11184
rect -865 -11184 -795 11184
rect -699 -11184 -629 11184
rect -533 -11184 -463 11184
rect -367 -11184 -297 11184
rect -201 -11184 -131 11184
rect -35 -11184 35 11184
rect 131 -11184 201 11184
rect 297 -11184 367 11184
rect 463 -11184 533 11184
rect 629 -11184 699 11184
rect 795 -11184 865 11184
rect 961 -11184 1031 11184
rect 1127 -11184 1197 11184
rect 1293 -11184 1363 11184
rect 1459 -11184 1529 11184
rect 1625 -11184 1695 11184
rect 1791 -11184 1861 11184
rect 1957 -11184 2027 11184
<< locali >>
rect -2157 11712 -2061 11746
rect 2061 11712 2157 11746
rect -2157 11650 -2123 11712
rect 2123 11650 2157 11712
rect -2157 -11712 -2123 -11650
rect 2123 -11712 2157 -11650
rect -2157 -11746 -2061 -11712
rect 2061 -11746 2157 -11712
<< viali >>
rect -2011 11201 -1973 11598
rect -1845 11201 -1807 11598
rect -1679 11201 -1641 11598
rect -1513 11201 -1475 11598
rect -1347 11201 -1309 11598
rect -1181 11201 -1143 11598
rect -1015 11201 -977 11598
rect -849 11201 -811 11598
rect -683 11201 -645 11598
rect -517 11201 -479 11598
rect -351 11201 -313 11598
rect -185 11201 -147 11598
rect -19 11201 19 11598
rect 147 11201 185 11598
rect 313 11201 351 11598
rect 479 11201 517 11598
rect 645 11201 683 11598
rect 811 11201 849 11598
rect 977 11201 1015 11598
rect 1143 11201 1181 11598
rect 1309 11201 1347 11598
rect 1475 11201 1513 11598
rect 1641 11201 1679 11598
rect 1807 11201 1845 11598
rect 1973 11201 2011 11598
rect -2011 -11598 -1973 -11201
rect -1845 -11598 -1807 -11201
rect -1679 -11598 -1641 -11201
rect -1513 -11598 -1475 -11201
rect -1347 -11598 -1309 -11201
rect -1181 -11598 -1143 -11201
rect -1015 -11598 -977 -11201
rect -849 -11598 -811 -11201
rect -683 -11598 -645 -11201
rect -517 -11598 -479 -11201
rect -351 -11598 -313 -11201
rect -185 -11598 -147 -11201
rect -19 -11598 19 -11201
rect 147 -11598 185 -11201
rect 313 -11598 351 -11201
rect 479 -11598 517 -11201
rect 645 -11598 683 -11201
rect 811 -11598 849 -11201
rect 977 -11598 1015 -11201
rect 1143 -11598 1181 -11201
rect 1309 -11598 1347 -11201
rect 1475 -11598 1513 -11201
rect 1641 -11598 1679 -11201
rect 1807 -11598 1845 -11201
rect 1973 -11598 2011 -11201
<< metal1 >>
rect -2017 11598 -1967 11610
rect -2017 11201 -2011 11598
rect -1973 11201 -1967 11598
rect -2017 11189 -1967 11201
rect -1851 11598 -1801 11610
rect -1851 11201 -1845 11598
rect -1807 11201 -1801 11598
rect -1851 11189 -1801 11201
rect -1685 11598 -1635 11610
rect -1685 11201 -1679 11598
rect -1641 11201 -1635 11598
rect -1685 11189 -1635 11201
rect -1519 11598 -1469 11610
rect -1519 11201 -1513 11598
rect -1475 11201 -1469 11598
rect -1519 11189 -1469 11201
rect -1353 11598 -1303 11610
rect -1353 11201 -1347 11598
rect -1309 11201 -1303 11598
rect -1353 11189 -1303 11201
rect -1187 11598 -1137 11610
rect -1187 11201 -1181 11598
rect -1143 11201 -1137 11598
rect -1187 11189 -1137 11201
rect -1021 11598 -971 11610
rect -1021 11201 -1015 11598
rect -977 11201 -971 11598
rect -1021 11189 -971 11201
rect -855 11598 -805 11610
rect -855 11201 -849 11598
rect -811 11201 -805 11598
rect -855 11189 -805 11201
rect -689 11598 -639 11610
rect -689 11201 -683 11598
rect -645 11201 -639 11598
rect -689 11189 -639 11201
rect -523 11598 -473 11610
rect -523 11201 -517 11598
rect -479 11201 -473 11598
rect -523 11189 -473 11201
rect -357 11598 -307 11610
rect -357 11201 -351 11598
rect -313 11201 -307 11598
rect -357 11189 -307 11201
rect -191 11598 -141 11610
rect -191 11201 -185 11598
rect -147 11201 -141 11598
rect -191 11189 -141 11201
rect -25 11598 25 11610
rect -25 11201 -19 11598
rect 19 11201 25 11598
rect -25 11189 25 11201
rect 141 11598 191 11610
rect 141 11201 147 11598
rect 185 11201 191 11598
rect 141 11189 191 11201
rect 307 11598 357 11610
rect 307 11201 313 11598
rect 351 11201 357 11598
rect 307 11189 357 11201
rect 473 11598 523 11610
rect 473 11201 479 11598
rect 517 11201 523 11598
rect 473 11189 523 11201
rect 639 11598 689 11610
rect 639 11201 645 11598
rect 683 11201 689 11598
rect 639 11189 689 11201
rect 805 11598 855 11610
rect 805 11201 811 11598
rect 849 11201 855 11598
rect 805 11189 855 11201
rect 971 11598 1021 11610
rect 971 11201 977 11598
rect 1015 11201 1021 11598
rect 971 11189 1021 11201
rect 1137 11598 1187 11610
rect 1137 11201 1143 11598
rect 1181 11201 1187 11598
rect 1137 11189 1187 11201
rect 1303 11598 1353 11610
rect 1303 11201 1309 11598
rect 1347 11201 1353 11598
rect 1303 11189 1353 11201
rect 1469 11598 1519 11610
rect 1469 11201 1475 11598
rect 1513 11201 1519 11598
rect 1469 11189 1519 11201
rect 1635 11598 1685 11610
rect 1635 11201 1641 11598
rect 1679 11201 1685 11598
rect 1635 11189 1685 11201
rect 1801 11598 1851 11610
rect 1801 11201 1807 11598
rect 1845 11201 1851 11598
rect 1801 11189 1851 11201
rect 1967 11598 2017 11610
rect 1967 11201 1973 11598
rect 2011 11201 2017 11598
rect 1967 11189 2017 11201
rect -2017 -11201 -1967 -11189
rect -2017 -11598 -2011 -11201
rect -1973 -11598 -1967 -11201
rect -2017 -11610 -1967 -11598
rect -1851 -11201 -1801 -11189
rect -1851 -11598 -1845 -11201
rect -1807 -11598 -1801 -11201
rect -1851 -11610 -1801 -11598
rect -1685 -11201 -1635 -11189
rect -1685 -11598 -1679 -11201
rect -1641 -11598 -1635 -11201
rect -1685 -11610 -1635 -11598
rect -1519 -11201 -1469 -11189
rect -1519 -11598 -1513 -11201
rect -1475 -11598 -1469 -11201
rect -1519 -11610 -1469 -11598
rect -1353 -11201 -1303 -11189
rect -1353 -11598 -1347 -11201
rect -1309 -11598 -1303 -11201
rect -1353 -11610 -1303 -11598
rect -1187 -11201 -1137 -11189
rect -1187 -11598 -1181 -11201
rect -1143 -11598 -1137 -11201
rect -1187 -11610 -1137 -11598
rect -1021 -11201 -971 -11189
rect -1021 -11598 -1015 -11201
rect -977 -11598 -971 -11201
rect -1021 -11610 -971 -11598
rect -855 -11201 -805 -11189
rect -855 -11598 -849 -11201
rect -811 -11598 -805 -11201
rect -855 -11610 -805 -11598
rect -689 -11201 -639 -11189
rect -689 -11598 -683 -11201
rect -645 -11598 -639 -11201
rect -689 -11610 -639 -11598
rect -523 -11201 -473 -11189
rect -523 -11598 -517 -11201
rect -479 -11598 -473 -11201
rect -523 -11610 -473 -11598
rect -357 -11201 -307 -11189
rect -357 -11598 -351 -11201
rect -313 -11598 -307 -11201
rect -357 -11610 -307 -11598
rect -191 -11201 -141 -11189
rect -191 -11598 -185 -11201
rect -147 -11598 -141 -11201
rect -191 -11610 -141 -11598
rect -25 -11201 25 -11189
rect -25 -11598 -19 -11201
rect 19 -11598 25 -11201
rect -25 -11610 25 -11598
rect 141 -11201 191 -11189
rect 141 -11598 147 -11201
rect 185 -11598 191 -11201
rect 141 -11610 191 -11598
rect 307 -11201 357 -11189
rect 307 -11598 313 -11201
rect 351 -11598 357 -11201
rect 307 -11610 357 -11598
rect 473 -11201 523 -11189
rect 473 -11598 479 -11201
rect 517 -11598 523 -11201
rect 473 -11610 523 -11598
rect 639 -11201 689 -11189
rect 639 -11598 645 -11201
rect 683 -11598 689 -11201
rect 639 -11610 689 -11598
rect 805 -11201 855 -11189
rect 805 -11598 811 -11201
rect 849 -11598 855 -11201
rect 805 -11610 855 -11598
rect 971 -11201 1021 -11189
rect 971 -11598 977 -11201
rect 1015 -11598 1021 -11201
rect 971 -11610 1021 -11598
rect 1137 -11201 1187 -11189
rect 1137 -11598 1143 -11201
rect 1181 -11598 1187 -11201
rect 1137 -11610 1187 -11598
rect 1303 -11201 1353 -11189
rect 1303 -11598 1309 -11201
rect 1347 -11598 1353 -11201
rect 1303 -11610 1353 -11598
rect 1469 -11201 1519 -11189
rect 1469 -11598 1475 -11201
rect 1513 -11598 1519 -11201
rect 1469 -11610 1519 -11598
rect 1635 -11201 1685 -11189
rect 1635 -11598 1641 -11201
rect 1679 -11598 1685 -11201
rect 1635 -11610 1685 -11598
rect 1801 -11201 1851 -11189
rect 1801 -11598 1807 -11201
rect 1845 -11598 1851 -11201
rect 1801 -11610 1851 -11598
rect 1967 -11201 2017 -11189
rect 1967 -11598 1973 -11201
rect 2011 -11598 2017 -11201
rect 1967 -11610 2017 -11598
<< properties >>
string FIXED_BBOX -2140 -11729 2140 11729
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 112 m 1 nx 25 wmin 0.350 lmin 0.50 rho 2000 val 641.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
