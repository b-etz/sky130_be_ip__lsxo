magic
tech sky130A
magscale 1 2
timestamp 1712782684
<< nwell >>
rect -458 -5359 458 5359
<< mvpmos >>
rect -200 4262 200 5062
rect -200 3226 200 4026
rect -200 2190 200 2990
rect -200 1154 200 1954
rect -200 118 200 918
rect -200 -918 200 -118
rect -200 -1954 200 -1154
rect -200 -2990 200 -2190
rect -200 -4026 200 -3226
rect -200 -5062 200 -4262
<< mvpdiff >>
rect -258 5050 -200 5062
rect -258 4274 -246 5050
rect -212 4274 -200 5050
rect -258 4262 -200 4274
rect 200 5050 258 5062
rect 200 4274 212 5050
rect 246 4274 258 5050
rect 200 4262 258 4274
rect -258 4014 -200 4026
rect -258 3238 -246 4014
rect -212 3238 -200 4014
rect -258 3226 -200 3238
rect 200 4014 258 4026
rect 200 3238 212 4014
rect 246 3238 258 4014
rect 200 3226 258 3238
rect -258 2978 -200 2990
rect -258 2202 -246 2978
rect -212 2202 -200 2978
rect -258 2190 -200 2202
rect 200 2978 258 2990
rect 200 2202 212 2978
rect 246 2202 258 2978
rect 200 2190 258 2202
rect -258 1942 -200 1954
rect -258 1166 -246 1942
rect -212 1166 -200 1942
rect -258 1154 -200 1166
rect 200 1942 258 1954
rect 200 1166 212 1942
rect 246 1166 258 1942
rect 200 1154 258 1166
rect -258 906 -200 918
rect -258 130 -246 906
rect -212 130 -200 906
rect -258 118 -200 130
rect 200 906 258 918
rect 200 130 212 906
rect 246 130 258 906
rect 200 118 258 130
rect -258 -130 -200 -118
rect -258 -906 -246 -130
rect -212 -906 -200 -130
rect -258 -918 -200 -906
rect 200 -130 258 -118
rect 200 -906 212 -130
rect 246 -906 258 -130
rect 200 -918 258 -906
rect -258 -1166 -200 -1154
rect -258 -1942 -246 -1166
rect -212 -1942 -200 -1166
rect -258 -1954 -200 -1942
rect 200 -1166 258 -1154
rect 200 -1942 212 -1166
rect 246 -1942 258 -1166
rect 200 -1954 258 -1942
rect -258 -2202 -200 -2190
rect -258 -2978 -246 -2202
rect -212 -2978 -200 -2202
rect -258 -2990 -200 -2978
rect 200 -2202 258 -2190
rect 200 -2978 212 -2202
rect 246 -2978 258 -2202
rect 200 -2990 258 -2978
rect -258 -3238 -200 -3226
rect -258 -4014 -246 -3238
rect -212 -4014 -200 -3238
rect -258 -4026 -200 -4014
rect 200 -3238 258 -3226
rect 200 -4014 212 -3238
rect 246 -4014 258 -3238
rect 200 -4026 258 -4014
rect -258 -4274 -200 -4262
rect -258 -5050 -246 -4274
rect -212 -5050 -200 -4274
rect -258 -5062 -200 -5050
rect 200 -4274 258 -4262
rect 200 -5050 212 -4274
rect 246 -5050 258 -4274
rect 200 -5062 258 -5050
<< mvpdiffc >>
rect -246 4274 -212 5050
rect 212 4274 246 5050
rect -246 3238 -212 4014
rect 212 3238 246 4014
rect -246 2202 -212 2978
rect 212 2202 246 2978
rect -246 1166 -212 1942
rect 212 1166 246 1942
rect -246 130 -212 906
rect 212 130 246 906
rect -246 -906 -212 -130
rect 212 -906 246 -130
rect -246 -1942 -212 -1166
rect 212 -1942 246 -1166
rect -246 -2978 -212 -2202
rect 212 -2978 246 -2202
rect -246 -4014 -212 -3238
rect 212 -4014 246 -3238
rect -246 -5050 -212 -4274
rect 212 -5050 246 -4274
<< mvnsubdiff >>
rect -392 5281 392 5293
rect -392 5247 -284 5281
rect 284 5247 392 5281
rect -392 5235 392 5247
rect -392 5185 -334 5235
rect -392 -5185 -380 5185
rect -346 -5185 -334 5185
rect 334 5185 392 5235
rect -392 -5235 -334 -5185
rect 334 -5185 346 5185
rect 380 -5185 392 5185
rect 334 -5235 392 -5185
rect -392 -5247 392 -5235
rect -392 -5281 -284 -5247
rect 284 -5281 392 -5247
rect -392 -5293 392 -5281
<< mvnsubdiffcont >>
rect -284 5247 284 5281
rect -380 -5185 -346 5185
rect 346 -5185 380 5185
rect -284 -5281 284 -5247
<< poly >>
rect -200 5143 200 5159
rect -200 5109 -184 5143
rect 184 5109 200 5143
rect -200 5062 200 5109
rect -200 4215 200 4262
rect -200 4181 -184 4215
rect 184 4181 200 4215
rect -200 4165 200 4181
rect -200 4107 200 4123
rect -200 4073 -184 4107
rect 184 4073 200 4107
rect -200 4026 200 4073
rect -200 3179 200 3226
rect -200 3145 -184 3179
rect 184 3145 200 3179
rect -200 3129 200 3145
rect -200 3071 200 3087
rect -200 3037 -184 3071
rect 184 3037 200 3071
rect -200 2990 200 3037
rect -200 2143 200 2190
rect -200 2109 -184 2143
rect 184 2109 200 2143
rect -200 2093 200 2109
rect -200 2035 200 2051
rect -200 2001 -184 2035
rect 184 2001 200 2035
rect -200 1954 200 2001
rect -200 1107 200 1154
rect -200 1073 -184 1107
rect 184 1073 200 1107
rect -200 1057 200 1073
rect -200 999 200 1015
rect -200 965 -184 999
rect 184 965 200 999
rect -200 918 200 965
rect -200 71 200 118
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -118 200 -71
rect -200 -965 200 -918
rect -200 -999 -184 -965
rect 184 -999 200 -965
rect -200 -1015 200 -999
rect -200 -1073 200 -1057
rect -200 -1107 -184 -1073
rect 184 -1107 200 -1073
rect -200 -1154 200 -1107
rect -200 -2001 200 -1954
rect -200 -2035 -184 -2001
rect 184 -2035 200 -2001
rect -200 -2051 200 -2035
rect -200 -2109 200 -2093
rect -200 -2143 -184 -2109
rect 184 -2143 200 -2109
rect -200 -2190 200 -2143
rect -200 -3037 200 -2990
rect -200 -3071 -184 -3037
rect 184 -3071 200 -3037
rect -200 -3087 200 -3071
rect -200 -3145 200 -3129
rect -200 -3179 -184 -3145
rect 184 -3179 200 -3145
rect -200 -3226 200 -3179
rect -200 -4073 200 -4026
rect -200 -4107 -184 -4073
rect 184 -4107 200 -4073
rect -200 -4123 200 -4107
rect -200 -4181 200 -4165
rect -200 -4215 -184 -4181
rect 184 -4215 200 -4181
rect -200 -4262 200 -4215
rect -200 -5109 200 -5062
rect -200 -5143 -184 -5109
rect 184 -5143 200 -5109
rect -200 -5159 200 -5143
<< polycont >>
rect -184 5109 184 5143
rect -184 4181 184 4215
rect -184 4073 184 4107
rect -184 3145 184 3179
rect -184 3037 184 3071
rect -184 2109 184 2143
rect -184 2001 184 2035
rect -184 1073 184 1107
rect -184 965 184 999
rect -184 37 184 71
rect -184 -71 184 -37
rect -184 -999 184 -965
rect -184 -1107 184 -1073
rect -184 -2035 184 -2001
rect -184 -2143 184 -2109
rect -184 -3071 184 -3037
rect -184 -3179 184 -3145
rect -184 -4107 184 -4073
rect -184 -4215 184 -4181
rect -184 -5143 184 -5109
<< locali >>
rect -380 5247 -284 5281
rect 284 5247 380 5281
rect -380 5185 -346 5247
rect 346 5185 380 5247
rect -200 5109 -184 5143
rect 184 5109 200 5143
rect -246 5050 -212 5066
rect -246 4258 -212 4274
rect 212 5050 246 5066
rect 212 4258 246 4274
rect -200 4181 -184 4215
rect 184 4181 200 4215
rect -200 4073 -184 4107
rect 184 4073 200 4107
rect -246 4014 -212 4030
rect -246 3222 -212 3238
rect 212 4014 246 4030
rect 212 3222 246 3238
rect -200 3145 -184 3179
rect 184 3145 200 3179
rect -200 3037 -184 3071
rect 184 3037 200 3071
rect -246 2978 -212 2994
rect -246 2186 -212 2202
rect 212 2978 246 2994
rect 212 2186 246 2202
rect -200 2109 -184 2143
rect 184 2109 200 2143
rect -200 2001 -184 2035
rect 184 2001 200 2035
rect -246 1942 -212 1958
rect -246 1150 -212 1166
rect 212 1942 246 1958
rect 212 1150 246 1166
rect -200 1073 -184 1107
rect 184 1073 200 1107
rect -200 965 -184 999
rect 184 965 200 999
rect -246 906 -212 922
rect -246 114 -212 130
rect 212 906 246 922
rect 212 114 246 130
rect -200 37 -184 71
rect 184 37 200 71
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -246 -130 -212 -114
rect -246 -922 -212 -906
rect 212 -130 246 -114
rect 212 -922 246 -906
rect -200 -999 -184 -965
rect 184 -999 200 -965
rect -200 -1107 -184 -1073
rect 184 -1107 200 -1073
rect -246 -1166 -212 -1150
rect -246 -1958 -212 -1942
rect 212 -1166 246 -1150
rect 212 -1958 246 -1942
rect -200 -2035 -184 -2001
rect 184 -2035 200 -2001
rect -200 -2143 -184 -2109
rect 184 -2143 200 -2109
rect -246 -2202 -212 -2186
rect -246 -2994 -212 -2978
rect 212 -2202 246 -2186
rect 212 -2994 246 -2978
rect -200 -3071 -184 -3037
rect 184 -3071 200 -3037
rect -200 -3179 -184 -3145
rect 184 -3179 200 -3145
rect -246 -3238 -212 -3222
rect -246 -4030 -212 -4014
rect 212 -3238 246 -3222
rect 212 -4030 246 -4014
rect -200 -4107 -184 -4073
rect 184 -4107 200 -4073
rect -200 -4215 -184 -4181
rect 184 -4215 200 -4181
rect -246 -4274 -212 -4258
rect -246 -5066 -212 -5050
rect 212 -4274 246 -4258
rect 212 -5066 246 -5050
rect -200 -5143 -184 -5109
rect 184 -5143 200 -5109
rect -380 -5247 -346 -5185
rect 346 -5247 380 -5185
rect -380 -5281 -284 -5247
rect 284 -5281 380 -5247
<< viali >>
rect -184 5109 184 5143
rect -246 4274 -212 5050
rect 212 4274 246 5050
rect -184 4181 184 4215
rect -184 4073 184 4107
rect -246 3238 -212 4014
rect 212 3238 246 4014
rect -184 3145 184 3179
rect -184 3037 184 3071
rect -246 2202 -212 2978
rect 212 2202 246 2978
rect -184 2109 184 2143
rect -184 2001 184 2035
rect -246 1166 -212 1942
rect 212 1166 246 1942
rect -184 1073 184 1107
rect -184 965 184 999
rect -246 130 -212 906
rect 212 130 246 906
rect -184 37 184 71
rect -184 -71 184 -37
rect -246 -906 -212 -130
rect 212 -906 246 -130
rect -184 -999 184 -965
rect -184 -1107 184 -1073
rect -246 -1942 -212 -1166
rect 212 -1942 246 -1166
rect -184 -2035 184 -2001
rect -184 -2143 184 -2109
rect -246 -2978 -212 -2202
rect 212 -2978 246 -2202
rect -184 -3071 184 -3037
rect -184 -3179 184 -3145
rect -246 -4014 -212 -3238
rect 212 -4014 246 -3238
rect -184 -4107 184 -4073
rect -184 -4215 184 -4181
rect -246 -5050 -212 -4274
rect 212 -5050 246 -4274
rect -184 -5143 184 -5109
<< metal1 >>
rect -196 5143 196 5149
rect -196 5109 -184 5143
rect 184 5109 196 5143
rect -196 5103 196 5109
rect -252 5050 -206 5062
rect -252 4274 -246 5050
rect -212 4274 -206 5050
rect -252 4262 -206 4274
rect 206 5050 252 5062
rect 206 4274 212 5050
rect 246 4274 252 5050
rect 206 4262 252 4274
rect -196 4215 196 4221
rect -196 4181 -184 4215
rect 184 4181 196 4215
rect -196 4175 196 4181
rect -196 4107 196 4113
rect -196 4073 -184 4107
rect 184 4073 196 4107
rect -196 4067 196 4073
rect -252 4014 -206 4026
rect -252 3238 -246 4014
rect -212 3238 -206 4014
rect -252 3226 -206 3238
rect 206 4014 252 4026
rect 206 3238 212 4014
rect 246 3238 252 4014
rect 206 3226 252 3238
rect -196 3179 196 3185
rect -196 3145 -184 3179
rect 184 3145 196 3179
rect -196 3139 196 3145
rect -196 3071 196 3077
rect -196 3037 -184 3071
rect 184 3037 196 3071
rect -196 3031 196 3037
rect -252 2978 -206 2990
rect -252 2202 -246 2978
rect -212 2202 -206 2978
rect -252 2190 -206 2202
rect 206 2978 252 2990
rect 206 2202 212 2978
rect 246 2202 252 2978
rect 206 2190 252 2202
rect -196 2143 196 2149
rect -196 2109 -184 2143
rect 184 2109 196 2143
rect -196 2103 196 2109
rect -196 2035 196 2041
rect -196 2001 -184 2035
rect 184 2001 196 2035
rect -196 1995 196 2001
rect -252 1942 -206 1954
rect -252 1166 -246 1942
rect -212 1166 -206 1942
rect -252 1154 -206 1166
rect 206 1942 252 1954
rect 206 1166 212 1942
rect 246 1166 252 1942
rect 206 1154 252 1166
rect -196 1107 196 1113
rect -196 1073 -184 1107
rect 184 1073 196 1107
rect -196 1067 196 1073
rect -196 999 196 1005
rect -196 965 -184 999
rect 184 965 196 999
rect -196 959 196 965
rect -252 906 -206 918
rect -252 130 -246 906
rect -212 130 -206 906
rect -252 118 -206 130
rect 206 906 252 918
rect 206 130 212 906
rect 246 130 252 906
rect 206 118 252 130
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect -252 -130 -206 -118
rect -252 -906 -246 -130
rect -212 -906 -206 -130
rect -252 -918 -206 -906
rect 206 -130 252 -118
rect 206 -906 212 -130
rect 246 -906 252 -130
rect 206 -918 252 -906
rect -196 -965 196 -959
rect -196 -999 -184 -965
rect 184 -999 196 -965
rect -196 -1005 196 -999
rect -196 -1073 196 -1067
rect -196 -1107 -184 -1073
rect 184 -1107 196 -1073
rect -196 -1113 196 -1107
rect -252 -1166 -206 -1154
rect -252 -1942 -246 -1166
rect -212 -1942 -206 -1166
rect -252 -1954 -206 -1942
rect 206 -1166 252 -1154
rect 206 -1942 212 -1166
rect 246 -1942 252 -1166
rect 206 -1954 252 -1942
rect -196 -2001 196 -1995
rect -196 -2035 -184 -2001
rect 184 -2035 196 -2001
rect -196 -2041 196 -2035
rect -196 -2109 196 -2103
rect -196 -2143 -184 -2109
rect 184 -2143 196 -2109
rect -196 -2149 196 -2143
rect -252 -2202 -206 -2190
rect -252 -2978 -246 -2202
rect -212 -2978 -206 -2202
rect -252 -2990 -206 -2978
rect 206 -2202 252 -2190
rect 206 -2978 212 -2202
rect 246 -2978 252 -2202
rect 206 -2990 252 -2978
rect -196 -3037 196 -3031
rect -196 -3071 -184 -3037
rect 184 -3071 196 -3037
rect -196 -3077 196 -3071
rect -196 -3145 196 -3139
rect -196 -3179 -184 -3145
rect 184 -3179 196 -3145
rect -196 -3185 196 -3179
rect -252 -3238 -206 -3226
rect -252 -4014 -246 -3238
rect -212 -4014 -206 -3238
rect -252 -4026 -206 -4014
rect 206 -3238 252 -3226
rect 206 -4014 212 -3238
rect 246 -4014 252 -3238
rect 206 -4026 252 -4014
rect -196 -4073 196 -4067
rect -196 -4107 -184 -4073
rect 184 -4107 196 -4073
rect -196 -4113 196 -4107
rect -196 -4181 196 -4175
rect -196 -4215 -184 -4181
rect 184 -4215 196 -4181
rect -196 -4221 196 -4215
rect -252 -4274 -206 -4262
rect -252 -5050 -246 -4274
rect -212 -5050 -206 -4274
rect -252 -5062 -206 -5050
rect 206 -4274 252 -4262
rect 206 -5050 212 -4274
rect 246 -5050 252 -4274
rect 206 -5062 252 -5050
rect -196 -5109 196 -5103
rect -196 -5143 -184 -5109
rect 184 -5143 196 -5109
rect -196 -5149 196 -5143
<< properties >>
string FIXED_BBOX -363 -5264 363 5264
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 2.0 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
