magic
tech sky130A
magscale 1 2
timestamp 1712849042
<< pwell >>
rect -201 -17922 201 17922
<< psubdiff >>
rect -165 17852 -69 17886
rect 69 17852 165 17886
rect -165 17790 -131 17852
rect 131 17790 165 17852
rect -165 -17852 -131 -17790
rect 131 -17852 165 -17790
rect -165 -17886 -69 -17852
rect 69 -17886 165 -17852
<< psubdiffcont >>
rect -69 17852 69 17886
rect -165 -17790 -131 17790
rect 131 -17790 165 17790
rect -69 -17886 69 -17852
<< xpolycontact >>
rect -35 17324 35 17756
rect -35 11924 35 12356
rect -35 11388 35 11820
rect -35 5988 35 6420
rect -35 5452 35 5884
rect -35 52 35 484
rect -35 -484 35 -52
rect -35 -5884 35 -5452
rect -35 -6420 35 -5988
rect -35 -11820 35 -11388
rect -35 -12356 35 -11924
rect -35 -17756 35 -17324
<< xpolyres >>
rect -35 12356 35 17324
rect -35 6420 35 11388
rect -35 484 35 5452
rect -35 -5452 35 -484
rect -35 -11388 35 -6420
rect -35 -17324 35 -12356
<< locali >>
rect -165 17852 -69 17886
rect 69 17852 165 17886
rect -165 17790 -131 17852
rect 131 17790 165 17852
rect -165 -17852 -131 -17790
rect 131 -17852 165 -17790
rect -165 -17886 -69 -17852
rect 69 -17886 165 -17852
<< viali >>
rect -19 17341 19 17738
rect -19 11942 19 12339
rect -19 11405 19 11802
rect -19 6006 19 6403
rect -19 5469 19 5866
rect -19 70 19 467
rect -19 -467 19 -70
rect -19 -5866 19 -5469
rect -19 -6403 19 -6006
rect -19 -11802 19 -11405
rect -19 -12339 19 -11942
rect -19 -17738 19 -17341
<< metal1 >>
rect -25 17738 25 17750
rect -25 17341 -19 17738
rect 19 17341 25 17738
rect -25 17329 25 17341
rect -25 12339 25 12351
rect -25 11942 -19 12339
rect 19 11942 25 12339
rect -25 11930 25 11942
rect -25 11802 25 11814
rect -25 11405 -19 11802
rect 19 11405 25 11802
rect -25 11393 25 11405
rect -25 6403 25 6415
rect -25 6006 -19 6403
rect 19 6006 25 6403
rect -25 5994 25 6006
rect -25 5866 25 5878
rect -25 5469 -19 5866
rect 19 5469 25 5866
rect -25 5457 25 5469
rect -25 467 25 479
rect -25 70 -19 467
rect 19 70 25 467
rect -25 58 25 70
rect -25 -70 25 -58
rect -25 -467 -19 -70
rect 19 -467 25 -70
rect -25 -479 25 -467
rect -25 -5469 25 -5457
rect -25 -5866 -19 -5469
rect 19 -5866 25 -5469
rect -25 -5878 25 -5866
rect -25 -6006 25 -5994
rect -25 -6403 -19 -6006
rect 19 -6403 25 -6006
rect -25 -6415 25 -6403
rect -25 -11405 25 -11393
rect -25 -11802 -19 -11405
rect 19 -11802 25 -11405
rect -25 -11814 25 -11802
rect -25 -11942 25 -11930
rect -25 -12339 -19 -11942
rect 19 -12339 25 -11942
rect -25 -12351 25 -12339
rect -25 -17341 25 -17329
rect -25 -17738 -19 -17341
rect 19 -17738 25 -17341
rect -25 -17750 25 -17738
<< properties >>
string FIXED_BBOX -148 -17869 148 17869
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 25 m 6 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 143.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
