magic
tech sky130A
magscale 1 2
timestamp 1712946411
<< pwell >>
rect -1825 -260 1825 260
<< nmos >>
rect -1629 -50 -29 50
rect 29 -50 1629 50
<< ndiff >>
rect -1687 38 -1629 50
rect -1687 -38 -1675 38
rect -1641 -38 -1629 38
rect -1687 -50 -1629 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 1629 38 1687 50
rect 1629 -38 1641 38
rect 1675 -38 1687 38
rect 1629 -50 1687 -38
<< ndiffc >>
rect -1675 -38 -1641 38
rect -17 -38 17 38
rect 1641 -38 1675 38
<< psubdiff >>
rect -1789 190 -1693 224
rect 1693 190 1789 224
rect -1789 128 -1755 190
rect 1755 128 1789 190
rect -1789 -190 -1755 -128
rect 1755 -190 1789 -128
rect -1789 -224 -1693 -190
rect 1693 -224 1789 -190
<< psubdiffcont >>
rect -1693 190 1693 224
rect -1789 -128 -1755 128
rect 1755 -128 1789 128
rect -1693 -224 1693 -190
<< poly >>
rect -1629 122 -29 138
rect -1629 88 -1613 122
rect -45 88 -29 122
rect -1629 50 -29 88
rect 29 122 1629 138
rect 29 88 45 122
rect 1613 88 1629 122
rect 29 50 1629 88
rect -1629 -88 -29 -50
rect -1629 -122 -1613 -88
rect -45 -122 -29 -88
rect -1629 -138 -29 -122
rect 29 -88 1629 -50
rect 29 -122 45 -88
rect 1613 -122 1629 -88
rect 29 -138 1629 -122
<< polycont >>
rect -1613 88 -45 122
rect 45 88 1613 122
rect -1613 -122 -45 -88
rect 45 -122 1613 -88
<< locali >>
rect -1789 190 -1693 224
rect 1693 190 1789 224
rect -1789 128 -1755 190
rect 1755 128 1789 190
rect -1629 88 -1613 122
rect -45 88 -29 122
rect 29 88 45 122
rect 1613 88 1629 122
rect -1675 38 -1641 54
rect -1675 -54 -1641 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 1641 38 1675 54
rect 1641 -54 1675 -38
rect -1629 -122 -1613 -88
rect -45 -122 -29 -88
rect 29 -122 45 -88
rect 1613 -122 1629 -88
rect -1789 -190 -1755 -128
rect 1755 -190 1789 -128
rect -1789 -224 -1693 -190
rect 1693 -224 1789 -190
<< viali >>
rect -1613 88 -45 122
rect 45 88 1613 122
rect -1675 -38 -1641 38
rect -17 -38 17 38
rect 1641 -38 1675 38
rect -1613 -122 -45 -88
rect 45 -122 1613 -88
<< metal1 >>
rect -1625 122 -33 128
rect -1625 88 -1613 122
rect -45 88 -33 122
rect -1625 82 -33 88
rect 33 122 1625 128
rect 33 88 45 122
rect 1613 88 1625 122
rect 33 82 1625 88
rect -1681 38 -1635 50
rect -1681 -38 -1675 38
rect -1641 -38 -1635 38
rect -1681 -50 -1635 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 1635 38 1681 50
rect 1635 -38 1641 38
rect 1675 -38 1681 38
rect 1635 -50 1681 -38
rect -1625 -88 -33 -82
rect -1625 -122 -1613 -88
rect -45 -122 -33 -88
rect -1625 -128 -33 -122
rect 33 -88 1625 -82
rect 33 -122 45 -88
rect 1613 -122 1625 -88
rect 33 -128 1625 -122
<< properties >>
string FIXED_BBOX -1772 -207 1772 207
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 8 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
