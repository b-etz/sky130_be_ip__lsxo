magic
tech sky130A
magscale 1 2
timestamp 1713210209
<< pwell >>
rect -296 -285 296 285
<< nmos >>
rect -100 -75 100 75
<< ndiff >>
rect -158 63 -100 75
rect -158 -63 -146 63
rect -112 -63 -100 63
rect -158 -75 -100 -63
rect 100 63 158 75
rect 100 -63 112 63
rect 146 -63 158 63
rect 100 -75 158 -63
<< ndiffc >>
rect -146 -63 -112 63
rect 112 -63 146 63
<< psubdiff >>
rect -260 215 -164 249
rect 164 215 260 249
rect -260 153 -226 215
rect 226 153 260 215
rect -260 -215 -226 -153
rect 226 -215 260 -153
rect -260 -249 -164 -215
rect 164 -249 260 -215
<< psubdiffcont >>
rect -164 215 164 249
rect -260 -153 -226 153
rect 226 -153 260 153
rect -164 -249 164 -215
<< poly >>
rect -100 147 100 163
rect -100 113 -84 147
rect 84 113 100 147
rect -100 75 100 113
rect -100 -113 100 -75
rect -100 -147 -84 -113
rect 84 -147 100 -113
rect -100 -163 100 -147
<< polycont >>
rect -84 113 84 147
rect -84 -147 84 -113
<< locali >>
rect -260 215 -164 249
rect 164 215 260 249
rect -260 153 -226 215
rect 226 153 260 215
rect -100 113 -84 147
rect 84 113 100 147
rect -146 63 -112 79
rect -146 -79 -112 -63
rect 112 63 146 79
rect 112 -79 146 -63
rect -100 -147 -84 -113
rect 84 -147 100 -113
rect -260 -215 -226 -153
rect 226 -215 260 -153
rect -260 -249 -164 -215
rect 164 -249 260 -215
<< viali >>
rect -84 113 84 147
rect -146 -63 -112 63
rect 112 -63 146 63
rect -84 -147 84 -113
<< metal1 >>
rect -96 147 96 153
rect -96 113 -84 147
rect 84 113 96 147
rect -96 107 96 113
rect -152 63 -106 75
rect -152 -63 -146 63
rect -112 -63 -106 63
rect -152 -75 -106 -63
rect 106 63 152 75
rect 106 -63 112 63
rect 146 -63 152 63
rect 106 -75 152 -63
rect -96 -113 96 -107
rect -96 -147 -84 -113
rect 84 -147 96 -113
rect -96 -153 96 -147
<< properties >>
string FIXED_BBOX -243 -232 243 232
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.75 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
