magic
tech sky130A
timestamp 1713210209
<< pwell >>
rect -297 -329 297 329
<< mvnmos >>
rect -183 -200 -133 200
rect -104 -200 -54 200
rect -25 -200 25 200
rect 54 -200 104 200
rect 133 -200 183 200
<< mvndiff >>
rect -212 194 -183 200
rect -212 -194 -206 194
rect -189 -194 -183 194
rect -212 -200 -183 -194
rect -133 194 -104 200
rect -133 -194 -127 194
rect -110 -194 -104 194
rect -133 -200 -104 -194
rect -54 194 -25 200
rect -54 -194 -48 194
rect -31 -194 -25 194
rect -54 -200 -25 -194
rect 25 194 54 200
rect 25 -194 31 194
rect 48 -194 54 194
rect 25 -200 54 -194
rect 104 194 133 200
rect 104 -194 110 194
rect 127 -194 133 194
rect 104 -200 133 -194
rect 183 194 212 200
rect 183 -194 189 194
rect 206 -194 212 194
rect 183 -200 212 -194
<< mvndiffc >>
rect -206 -194 -189 194
rect -127 -194 -110 194
rect -48 -194 -31 194
rect 31 -194 48 194
rect 110 -194 127 194
rect 189 -194 206 194
<< mvpsubdiff >>
rect -279 305 279 311
rect -279 288 -225 305
rect 225 288 279 305
rect -279 282 279 288
rect -279 257 -250 282
rect -279 -257 -273 257
rect -256 -257 -250 257
rect 250 257 279 282
rect -279 -282 -250 -257
rect 250 -257 256 257
rect 273 -257 279 257
rect 250 -282 279 -257
rect -279 -288 279 -282
rect -279 -305 -225 -288
rect 225 -305 279 -288
rect -279 -311 279 -305
<< mvpsubdiffcont >>
rect -225 288 225 305
rect -273 -257 -256 257
rect 256 -257 273 257
rect -225 -305 225 -288
<< poly >>
rect -183 236 -133 244
rect -183 219 -175 236
rect -141 219 -133 236
rect -183 200 -133 219
rect -104 236 -54 244
rect -104 219 -96 236
rect -62 219 -54 236
rect -104 200 -54 219
rect -25 236 25 244
rect -25 219 -17 236
rect 17 219 25 236
rect -25 200 25 219
rect 54 236 104 244
rect 54 219 62 236
rect 96 219 104 236
rect 54 200 104 219
rect 133 236 183 244
rect 133 219 141 236
rect 175 219 183 236
rect 133 200 183 219
rect -183 -219 -133 -200
rect -183 -236 -175 -219
rect -141 -236 -133 -219
rect -183 -244 -133 -236
rect -104 -219 -54 -200
rect -104 -236 -96 -219
rect -62 -236 -54 -219
rect -104 -244 -54 -236
rect -25 -219 25 -200
rect -25 -236 -17 -219
rect 17 -236 25 -219
rect -25 -244 25 -236
rect 54 -219 104 -200
rect 54 -236 62 -219
rect 96 -236 104 -219
rect 54 -244 104 -236
rect 133 -219 183 -200
rect 133 -236 141 -219
rect 175 -236 183 -219
rect 133 -244 183 -236
<< polycont >>
rect -175 219 -141 236
rect -96 219 -62 236
rect -17 219 17 236
rect 62 219 96 236
rect 141 219 175 236
rect -175 -236 -141 -219
rect -96 -236 -62 -219
rect -17 -236 17 -219
rect 62 -236 96 -219
rect 141 -236 175 -219
<< locali >>
rect -273 288 -225 305
rect 225 288 273 305
rect -273 257 -256 288
rect 256 257 273 288
rect -183 219 -175 236
rect -141 219 -133 236
rect -104 219 -96 236
rect -62 219 -54 236
rect -25 219 -17 236
rect 17 219 25 236
rect 54 219 62 236
rect 96 219 104 236
rect 133 219 141 236
rect 175 219 183 236
rect -206 194 -189 202
rect -206 -202 -189 -194
rect -127 194 -110 202
rect -127 -202 -110 -194
rect -48 194 -31 202
rect -48 -202 -31 -194
rect 31 194 48 202
rect 31 -202 48 -194
rect 110 194 127 202
rect 110 -202 127 -194
rect 189 194 206 202
rect 189 -202 206 -194
rect -183 -236 -175 -219
rect -141 -236 -133 -219
rect -104 -236 -96 -219
rect -62 -236 -54 -219
rect -25 -236 -17 -219
rect 17 -236 25 -219
rect 54 -236 62 -219
rect 96 -236 104 -219
rect 133 -236 141 -219
rect 175 -236 183 -219
rect -273 -288 -256 -257
rect 256 -288 273 -257
rect -273 -305 -225 -288
rect 225 -305 273 -288
<< properties >>
string FIXED_BBOX -264 -296 264 296
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 0.5 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
