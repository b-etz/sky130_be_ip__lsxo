magic
tech sky130A
magscale 1 2
timestamp 1713104671
<< metal3 >>
rect -2186 -2040 1882 2040
<< mimcap >>
rect -2146 1960 1854 2000
rect -2146 -1960 -2106 1960
rect 1814 -1960 1854 1960
rect -2146 -2000 1854 -1960
<< mimcapcontact >>
rect -2106 -1960 1814 1960
<< metal4 >>
rect -2107 1960 1815 1961
rect -2107 -1960 -2106 1960
rect 1814 -1960 1815 1960
rect -2107 -1961 1815 -1960
<< properties >>
string FIXED_BBOX -2186 -2040 1894 2040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 20 l 20 val 815.2 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
