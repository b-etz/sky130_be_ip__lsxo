* NGSPICE file created from sky130_be_ip__lsxo_rcx.ext - technology: sky130A

.subckt sky130_be_ip__lsxo_rcx ibias dout xout xin ena avss avdd standby dvss dvdd
X0 a_16620_n1869# a_15705_n2241# a_16273_n2273# dvss.t4 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1 a_20376_n2791# x7.stby_done_b dvdd.t109 dvdd.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_21036_n1869# a_19955_n2241# a_20689_n2273# dvdd.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3 a_10620_n8338# a_24220_n8172# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X4 a_16795_n2817# a_16620_n2791# a_16974_n2791# dvss.t146 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5 dvdd.t74 ena_ip x3.in_b dvdd.t73 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X6 dvdd.t164 a_21036_n1869# a_21211_n1943# dvdd.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_18828_n2791# a_17913_n2791# a_18481_n2549# dvss.t159 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X8 a_2130_n19848# a_24530_n20014# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X9 vbreg icnode a_11526_n12394# avss_ip.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X10 x7.x2.x2.CLK a_15000_n2791# dvss.t24 dvss.t23 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X11 a_18168_n1881# x7.x1.Qb2 dvss.t81 dvss.t80 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X12 tail vbp dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X13 a_16317_n2791# a_16273_n2549# a_16151_n2791# dvss.t147 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X14 dvss.t74 standby_b dvss_ip dvss.t73 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X15 a_9120_n9346.t0 a_24220_n9832# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X16 a_16795_n1943# a_16620_n1869# a_16974_n1881# dvss.t179 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X17 x7.ena_done_b a_21775_n2247# dvdd.t133 dvdd.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X18 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X19 a_20121_n2241# a_19955_n2241# dvdd.t85 dvdd.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_2130_n21176# a_24530_n21342# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X21 ibias_ip standby_33 ibias.t1 ibias.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X22 xout.t19 vbreg avdd_ip.t26 avdd_ip.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X23 inv_m1 inv_in.t1 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X24 a_2132_n15590# a_18932_n15756# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X25 dout_ip inv_m2 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X26 a_20733_n2791# a_20689_n2549# a_20567_n2791# dvss.t2 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X27 inv_in.t2 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X28 x7.x1.x2.CLK a_15000_n1881# dvss.t1 dvss.t0 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X29 avdd_ip.t29 avss_ip.t52 sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X30 a_16317_n1881# a_16273_n2273# a_16151_n1869# dvss.t101 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X31 x7.stby_done_b a_21775_n2791# dvss.t26 dvss.t25 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X32 a_14009_n2701# x7.clk_disable dvss.t208 dvss.t82 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.07665 ps=0.785 w=0.42 l=0.15
X33 dvss.t196 standby_ip standby_b dvss.t195 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X34 dvss.t205 a_2971_n1521# ena_ip dvss.t204 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X35 dvss.t72 standby_b a_16317_n2791# dvss.t71 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X36 avdd_ip.t30 avss_ip.t33 sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X37 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X38 dvss.t22 x7.ena_done_b a_14035_n1997# dvss.t21 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X39 x7.stby_done_b a_21775_n2791# dvdd.t24 dvdd.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X40 a_2132_n17582# a_18932_n17416# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X41 inv_m1 inv_in.t3 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X42 avss.t26 avdd.t19 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X43 a_10620_n9666# a_24220_n9832# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X44 a_20733_n1881# a_20689_n2273# a_20567_n1869# dvss.t153 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X45 dvdd.t9 x7.x2.x2.CLK a_15539_n2791# dvdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X46 a_16782_n2425# a_15705_n2791# a_16620_n2791# dvdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X47 dvdd_ip inv_m1 inv_m2 dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X48 a_4857_n1521# standby.t0 dvdd.t132 dvdd.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X49 avdd_ip.t2 x3.out_b.t3 avdd.t9 avdd.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X50 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X51 a_20121_n2791# a_19955_n2791# dvss.t169 dvss.t168 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X52 dvss.t98 ena_ip a_16317_n1881# dvss.t97 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X53 x7.x1.Qb2 a_19567_n2247# dvss.t76 dvss.t75 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X54 dvss.t185 ena.t0 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X55 dvdd.t80 a_19003_n2817# a_19567_n2791# dvdd.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X56 avss_ip.t57 vg1.t2 vg1.t3 avss_ip.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X57 a_21145_n1869# a_19955_n2241# a_21036_n1869# dvss.t113 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X58 avdd_ip.t25 vbreg avdd_ip.t24 avdd_ip.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X59 a_21211_n2817# standby_b dvdd.t55 dvdd.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X60 avss_ip.t30 xin.t6 avss_ip.t29 avss_ip.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0 ps=0 w=4 l=0.5
X61 a_19003_n2817# a_18828_n2791# a_19182_n2791# dvss.t180 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X62 a_15000_n1881# dout_ip dvdd.t65 dvdd.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
X63 a_2132_n17250# a_18932_n17416# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X64 a_20121_n2241# a_19955_n2241# dvss.t112 dvss.t111 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X65 dvss_ip ibias_ip dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=5.8 ps=45.8 w=2 l=2
X66 a_10620_n9666# a_24220_n9500# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X67 a_18359_n1869# a_17913_n2241# a_18263_n1869# dvss.t152 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X68 xout.t18 vbreg avdd_ip.t23 avdd_ip.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X69 avss_ip.t11 avss_ip.t12 avss_ip.t0 sky130_fd_pr__res_xhigh_po_0p35 l=75
X70 vbreg vg2.t5 vrb.t4 avss_ip.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X71 a_18525_n2791# a_18481_n2549# a_18359_n2791# dvss.t186 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X72 a_2130_n20844# a_24530_n21010# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X73 a_15083_n2791# dout_ip a_15000_n2791# dvss.t84 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X74 a_21036_n1869# a_20121_n2241# a_20689_n2273# dvss.t182 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X75 dvss_ip standby_b dvss.t70 dvss.t69 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X76 a_2132_n15590# a_18932_n15424# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X77 a_14285_n2079# x7.ena_done_b a_14285_n2281# dvdd.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X78 a_19003_n1943# a_18828_n1869# a_19182_n1881# dvss.t150 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X79 vn xin.t7 vn dvdd_ip sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=2.32 ps=17.16 w=4 l=2
X80 avss.t7 standby_b standby_33 avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X81 a_10620_n7674# a_24220_n7840# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X82 ibias_ip ibias_ip dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X83 avdd.t14 x3.out_b.t4 avdd_ip.t27 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X84 a_15960_n2791# x7.x2.Qb1 dvdd.t98 dvdd.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X85 a_2130_n19516# a_24530_n19682# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X86 xin.t8 avdd_ip.t28 sky130_fd_pr__diode_pd2nw_05v5 perim=1.8e+06 area=2.025e+11
X87 a_20579_n2247# ena_ip dvdd.t72 dvdd.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X88 dvdd.t167 a_2971_n1521# ena_ip dvdd.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X89 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X90 a_15083_n1881# dout_ip a_15000_n1881# dvss.t83 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X91 a_18525_n1881# a_18481_n2273# a_18359_n1869# dvss.t33 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X92 a_18168_n2791# x7.x2.Qb2 dvdd.t102 dvdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X93 dvss.t68 standby_b a_18525_n2791# dvss.t67 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X94 xin_buf xout.t23 tail dvdd_ip sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X95 a_16273_n2549# a_16055_n2791# dvdd.t82 dvdd.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X96 dvss.t145 x7.stby_done_b a_15083_n2791# dvss.t144 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X97 xout.t22 xin.t9 avss_ip.t62 avss_ip.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X98 x7.x1.x4.Q a_21211_n1943# dvss.t165 dvss.t164 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X99 dvdd.t108 x7.stby_done_b a_15000_n2791# dvdd.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X100 a_14009_n2404# standby_ip a_14285_n2079# dvdd.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X101 dvss_ip standby_b dvss.t66 dvss.t65 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X102 avdd_ip.t19 vbreg xout.t17 avdd_ip.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X103 tail vbp dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X104 a_2130_n20844# a_24530_n20678# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X105 a_16729_n1869# a_15539_n2241# a_16620_n1869# dvss.t42 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X106 avss_ip.t63 vg2.t4 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X107 dvdd_ip vbp dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=19.865 ps=155.56 w=2 l=2
X108 a_16273_n2273# a_16055_n1869# dvdd.t105 dvdd.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X109 a_2132_n15258# a_18932_n15424# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X110 a_18990_n2425# a_17913_n2791# a_18828_n2791# dvdd.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X111 a_14285_n2281# x7.stby_done_b dvdd.t107 dvdd.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X112 avdd_ip.t22 vbreg avdd_ip.t21 avdd_ip.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X113 dvss.t96 ena_ip a_18525_n1881# dvss.t95 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X114 dvdd.t125 a_21211_n1943# a_21775_n2247# dvdd.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X115 dvss.t20 x7.ena_done_b a_15083_n1881# dvss.t19 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X116 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X117 a_16795_n1943# ena_ip dvdd.t71 dvdd.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X118 dvss.t154 standby.t1 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X119 dvss.t64 standby_b dvss_ip dvss.t63 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X120 a_2130_n19516# a_24530_n19350# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X121 dvdd.t38 a_14009_n2404# x7.clk_disable dvdd.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X122 avss_ip.t9 avss_ip.t10 avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X123 dvdd_ip standby_ip dvdd.t162 dvdd.t161 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X124 a_16163_n2247# ena_ip dvdd.t70 dvdd.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X125 a_2132_n16918# a_18932_n17084# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X126 dvdd.t101 x7.x2.Qb2 a_19955_n2791# dvdd.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X127 a_19003_n1943# ena_ip dvdd.t69 dvdd.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X128 inv_in.t4 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X129 a_10620_n9334# a_24220_n9500# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X130 dvss.t126 a_21211_n2817# a_21775_n2791# dvss.t125 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X131 a_3134_n13324# vrb.t0 avss_ip.t0 sky130_fd_pr__res_xhigh_po_0p35 l=75
X132 dvdd_ip standby_ip dvdd.t160 dvdd.t159 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X133 a_16974_n2791# standby_b dvss.t62 dvss.t61 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X134 x7.x1.x2.Q a_16795_n1943# dvss.t14 dvss.t13 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X135 a_2132_n17582# a_18932_n17748# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X136 dvdd.t16 x7.x1.x2.CLK a_15539_n2241# dvdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X137 dvdd_ip vbp tail dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X138 a_19182_n2791# standby_b dvss.t60 dvss.t59 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X139 dvss.t107 a_19003_n2817# a_18937_n2791# dvss.t106 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X140 avss_ip.t51 avss_ip.t49 avss_ip.t50 avss_ip.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X141 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X142 dout_ip inv_m2 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X143 a_15705_n2791# a_15539_n2791# dvdd.t36 dvdd.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X144 avdd.t15 x3.out_b.t5 x3.out.t2 avdd.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X145 dvdd.t174 a_16795_n2817# a_16782_n2425# dvdd.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X146 dvss.t163 a_21211_n1943# a_21775_n2247# dvss.t162 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X147 xout.t3 xin.t10 avss_ip.t20 avss_ip.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X148 avss_ip.t48 avss_ip.t46 avss_ip.t47 avss_ip.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X149 a_16974_n1881# ena_ip dvss.t94 dvss.t93 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X150 dvdd.t15 a_16795_n1943# a_17359_n2247# dvdd.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X151 xin.t0 a_24530_n22338# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X152 avss_ip.t14 x3.out.t3 avss.t15 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X153 dvss.t207 x7.clk_disable dout_filt dvss.t206 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X154 a_16055_n2791# a_15539_n2791# a_15960_n2791# dvss.t37 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X155 dvdd.t158 standby_ip dvdd_ip dvdd.t157 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X156 standby_33 x4.out_b.t3 avdd.t10 avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X157 a_16055_n1869# a_15705_n2241# a_15960_n1881# dvdd.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X158 dvdd_ip vbp tail dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X159 a_20471_n2791# a_20121_n2791# a_20376_n2791# dvdd.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X160 avss_ip.t25 xout.t24 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
**devattr s=257843176,88584 d=257843176,88584
X161 tail vbp dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X162 dvdd.t79 a_19003_n2817# a_18990_n2425# dvdd.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X163 a_10620_n9334# a_24220_n9168# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X164 a_19182_n1881# ena_ip dvss.t92 dvss.t91 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X165 avdd_ip.t20 vbreg xout.t16 avdd_ip.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X166 avss_ip.t21 xin.t11 xout.t4 avss_ip.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X167 xin_buf xout.t25 xin_buf dvdd_ip sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=2.32 ps=17.16 w=4 l=2
X168 a_3134_n13324# avss_ip.t1 avss_ip.t0 sky130_fd_pr__res_xhigh_po_0p35 l=75
X169 a_21036_n2791# a_19955_n2791# a_20689_n2549# dvdd.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X170 dvss.t32 a_19003_n1943# a_18937_n1869# dvss.t31 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X171 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X172 a_18937_n2791# a_17747_n2791# a_18828_n2791# dvss.t191 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X173 dvss.t214 a_16795_n2817# a_17359_n2791# dvss.t213 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X174 a_16273_n2273# a_16055_n1869# dvss.t140 dvss.t139 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X175 dvdd.t135 a_16620_n1869# a_16795_n1943# dvdd.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X176 x7.x1.x2.Q a_16795_n1943# dvdd.t13 dvdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X177 a_2130_n20512# a_24530_n20678# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X178 avss_ip.t5 xin.t12 xout.t0 avss_ip.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X179 dvdd.t122 a_21036_n2791# a_21211_n2817# dvdd.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X180 x4.out_b.t2 standby_ip avss.t25 avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X181 a_18481_n2549# a_18263_n2791# dvdd.t165 dvdd.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X182 dvss_ip inv_m1 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=7.9025 ps=61.46 w=0.5 l=1
X183 ibias_ip ibias_ip dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X184 dvss.t8 x7.x2.x2.CLK a_15539_n2791# dvss.t7 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X185 xout.t1 xin.t13 avss_ip.t6 avss_ip.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X186 a_2132_n14926# a_18932_n15092# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X187 dvdd.t171 x7.clk_disable a_14357_n2743# dvdd.t170 sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.005 as=0.0672 ps=0.85 w=0.64 l=0.15
X188 vn vn vn dvss_ip sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=2.32 ps=17.16 w=4 l=2
X189 a_20567_n2791# a_20121_n2791# a_20471_n2791# dvss.t184 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X190 dvdd.t156 standby_ip dvdd_ip dvdd.t155 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X191 dvss_ip dout_filt dout.t1 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=1
X192 a_20471_n1869# a_19955_n2241# a_20376_n1881# dvss.t110 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X193 a_18481_n2273# a_18263_n1869# dvdd.t100 dvdd.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X194 avss.t13 x3.out.t4 avss_ip.t13 avss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X195 dvss.t12 a_16795_n1943# a_17359_n2247# dvss.t11 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X196 x7.x1.Qb1 a_17359_n2247# dvdd.t104 dvdd.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X197 dvdd_ip vbp tail dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X198 avss.t27 avdd.t18 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X199 x7.x2.x2.Q a_16795_n2817# dvdd.t173 dvdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X200 a_14035_n2743# dout_ip dout_filt dvss.t82 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X201 dvss.t16 x7.x1.x2.CLK a_15539_n2241# dvss.t15 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X202 dout_ip inv_m2 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X203 xin_buf vn dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X204 avdd_ip.t18 vbreg vg1.t1 avdd_ip.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X205 a_2130_n19848# a_24530_n19682# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X206 vrb.t3 vg2.t6 vbreg avss_ip.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X207 a_18828_n1869# a_17913_n2241# a_18481_n2273# dvss.t151 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X208 x7.x2.Qb1 a_17359_n2791# dvss.t178 dvss.t177 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X209 a_2130_n20512# a_24530_n20346# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X210 dvdd.t118 a_20689_n2273# a_20579_n2247# dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X211 x7.x1.x2.CLK a_15000_n1881# dvdd.t1 dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X212 dvdd_ip standby_ip dvdd.t154 dvdd.t153 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X213 a_2132_n14926# a_18932_n14760# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X214 x7.x2.Qb1 a_17359_n2791# dvdd.t134 dvdd.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X215 x7.x1.x3.Q a_19003_n1943# dvss.t30 dvss.t29 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X216 xout.t8 xin.t14 avss_ip.t38 avss_ip.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X217 avdd.t1 x3.out_b.t6 avdd_ip.t0 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X218 a_16273_n2549# a_16055_n2791# dvss.t109 dvss.t108 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X219 a_16151_n2791# a_15705_n2791# a_16055_n2791# dvss.t203 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X220 vg1.t4 xin.t5 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X221 avss_ip.t39 xin.t15 xout.t9 avss_ip.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X222 dvss_ip inv_m1 inv_m2 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X223 a_2130_n19184# a_24530_n19018# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X224 dvdd_ip vbp dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X225 inv_in.t5 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X226 dvdd.t120 a_4857_n1521# standby_ip dvdd.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X227 a_14035_n1997# ena_ip a_14009_n2404# dvss.t21 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X228 a_17913_n2791# a_17747_n2791# dvdd.t140 dvdd.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X229 a_4857_n1521# standby.t2 dvss.t170 dvss.t155 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X230 a_10620_n9002# a_24220_n9168# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X231 a_18263_n2791# a_17747_n2791# a_18168_n2791# dvss.t190 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X232 a_14009_n2404# standby_b a_14035_n2281# dvss.t21 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X233 a_16620_n1869# a_15539_n2241# a_16273_n2273# dvdd.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X234 a_18263_n1869# a_17913_n2241# a_18168_n1881# dvdd.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X235 a_10620_n9002# a_24220_n8836# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X236 dvdd.t61 x7.x1.Qb2 a_19955_n2241# dvdd.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X237 a_2130_n20180# a_24530_n20346# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X238 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X239 x3.out_b.t2 x3.out.t5 avdd.t7 avdd.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X240 xout.t6 xin.t16 avss_ip.t36 avss_ip.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X241 avdd.t5 standby_33 x4.out_b.t0 avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X242 a_20579_n2247# a_19955_n2241# a_20471_n1869# dvdd.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X243 dvdd.t77 a_16273_n2273# a_16163_n2247# dvdd.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X244 a_15000_n2791# dout_ip dvdd.t64 dvdd.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
X245 dvdd.t115 a_18828_n1869# a_19003_n1943# dvdd.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X246 a_2130_n22172# a_24530_n22006# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X247 avss_ip.t37 xin.t17 xout.t7 avss_ip.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X248 avdd_ip.t31 avss_ip.t34 sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X249 a_15705_n2241# a_15539_n2241# dvdd.t41 dvdd.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X250 a_2130_n21840# a_24530_n22006# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X251 avdd_ip.t17 vbreg xout.t15 avdd_ip.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X252 dvdd.t97 x7.x2.Qb1 a_17747_n2791# dvdd.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X253 a_2132_n16586# a_18932_n16420# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X254 avss_ip.t27 xin.t18 avss_ip.t26 avss_ip.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X255 a_10620_n8670# a_24220_n8836# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X256 xin_buf vn xin_buf dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=2.32 ps=17.16 w=4 l=2
X257 x7.x1.Qb2 a_19567_n2247# dvdd.t57 dvdd.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X258 a_2132_n17250# a_18932_n17084# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X259 a_14009_n2701# x7.clk_disable dvdd.t169 dvdd.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.10855 ps=1.005 w=0.42 l=0.15
X260 dvss.t136 x7.x2.Qb2 a_19955_n2791# dvss.t135 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X261 dvss.t194 standby_ip dout_ip dvss.t193 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X262 dvss_ip ibias_ip vbp dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X263 inv_in.t6 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X264 a_22601_n15524# vbreg a_22601_n15524# avdd_ip.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=2.32 ps=17.16 w=4 l=2
X265 a_20579_n2425# standby_b dvdd.t53 dvdd.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X266 a_16163_n2247# a_15539_n2241# a_16055_n1869# dvdd.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X267 avss_ip.t28 xin.t19 xout.t5 avss_ip.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X268 x7.x2.Qb2 a_19567_n2791# dvss.t149 dvss.t148 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X269 vbreg vg1.t5 vbreg avss_ip.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=7.0818 ps=52.9 w=4 l=2
X270 vg1.t6 xin.t4 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X271 avss_ip.t31 x3.out.t6 avss.t19 avss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X272 x3.in_b ena_ip dvss.t90 dvss.t89 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X273 x7.x2.Qb2 a_19567_n2791# dvdd.t113 dvdd.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X274 dvss.t79 x7.x1.Qb2 a_19955_n2241# dvss.t78 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X275 a_15705_n2791# a_15539_n2791# dvss.t36 dvss.t35 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X276 standby_33 standby_b avss.t5 avss.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X277 vbreg vg2.t7 vrb.t2 avss_ip.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X278 tail xin.t20 vn dvdd_ip sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X279 dout_ip inv_m2 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X280 dvdd.t175 dvss.t77 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X281 dvdd.t124 a_21211_n1943# a_21198_n2247# dvdd.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X282 a_2130_n20180# a_24530_n20014# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X283 dvdd_ip vbp dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X284 a_20376_n2791# x7.stby_done_b dvss.t143 dvss.t142 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X285 a_18828_n1869# a_17747_n2241# a_18481_n2273# dvdd.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X286 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X287 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X288 a_16795_n2817# standby_b dvdd.t51 dvdd.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X289 a_2132_n14594# a_18932_n14428# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X290 a_15705_n2241# a_15539_n2241# dvss.t41 dvss.t40 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X291 x3.out.t1 x3.in_b avss.t3 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X292 a_16163_n2425# standby_b dvdd.t49 dvdd.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X293 inv_in.t7 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X294 a_2132_n15258# a_18932_n15092# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X295 a_19003_n2817# standby_b dvdd.t47 dvdd.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X296 dvdd.t32 a_18481_n2273# a_18371_n2247# dvdd.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X297 avss_ip.t60 avss_ip.t61 avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X298 a_20376_n1881# x7.ena_done_b dvss.t18 dvss.t17 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X299 dvdd_ip inv_m1 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=1
X300 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X301 dvss.t58 standby_b dvss_ip dvss.t57 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X302 vg1.t7 xin.t3 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X303 a_2130_n19184# a_24530_n19350# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X304 a_10620_n8670# a_24220_n8504# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X305 a_17913_n2241# a_17747_n2241# dvdd.t129 dvdd.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X306 x7.x2.x4.Q a_21211_n2817# dvss.t124 dvss.t123 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X307 dvss_ip ibias_ip ibias_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X308 a_21198_n2247# a_20121_n2241# a_21036_n1869# dvdd.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X309 a_20689_n2273# a_20471_n1869# dvss.t6 dvss.t5 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X310 x7.x1.x4.Q a_21211_n1943# dvdd.t123 dvdd.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X311 xout.t21 vbreg xout.t20 avdd_ip.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X312 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X313 a_2132_n16918# a_18932_n16752# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X314 avss_ip.t64 vg2.t3 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X315 a_16055_n2791# a_15705_n2791# a_15960_n2791# dvdd.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X316 avss_ip.t22 avss_ip.t23 avss_ip.t0 sky130_fd_pr__res_xhigh_po_0p35 l=75
X317 avss.t1 x3.in_b x3.out.t0 avss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X318 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X319 dvss_ip standby_b dvss.t56 dvss.t55 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X320 a_18371_n2247# ena_ip dvdd.t68 dvdd.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X321 a_2130_n21508# a_24530_n21674# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X322 a_18371_n2247# a_17747_n2241# a_18263_n1869# dvdd.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X323 vbreg vbreg avdd_ip.t16 avdd_ip.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X324 a_16620_n2791# a_15705_n2791# a_16273_n2549# dvss.t202 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X325 x7.x2.x4.Q a_21211_n2817# dvdd.t96 dvdd.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X326 dvdd.t111 a_16620_n2791# a_16795_n2817# dvdd.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X327 dvss_ip standby_b dvss.t54 dvss.t53 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X328 a_2130_n22172# a_24530_n22338# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X329 a_10620_n8338# a_24220_n8504# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X330 dvdd.t90 x7.x1.Qb1 a_17747_n2241# dvdd.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X331 dvdd.t152 standby_ip dvdd_ip dvdd.t151 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X332 inv_in.t8 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X333 a_2132_n16586# a_18932_n16752# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X334 a_17913_n2791# a_17747_n2791# dvss.t189 dvss.t188 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X335 a_16055_n1869# a_15539_n2241# a_15960_n1881# dvss.t39 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X336 x7.x2.x2.Q a_16795_n2817# dvss.t212 dvss.t211 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X337 avdd_ip.t32 avss_ip.t35 sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X338 x7.ena_done_b a_21775_n2247# dvss.t176 dvss.t175 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X339 avss_ip.t65 vg2.t2 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X340 avss_ip.t45 avss_ip.t43 avss_ip.t44 avss_ip.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X341 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X342 a_20689_n2549# a_20471_n2791# dvss.t100 dvss.t99 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X343 dvss.t52 standby_b dvss_ip dvss.t51 sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X344 dvdd.t30 a_19003_n1943# a_19567_n2247# dvdd.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X345 dvdd_ip a_9120_n9346.t1 a_9120_n9346.t2 dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X346 dvdd.t94 a_21211_n2817# a_21775_n2791# dvdd.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X347 a_20376_n1881# x7.ena_done_b dvdd.t20 dvdd.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X348 a_18937_n1869# a_17747_n2241# a_18828_n1869# dvss.t174 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X349 avss_ip.t7 xin.t21 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
**devattr s=257843176,88584 d=257843176,88584
X350 dvdd_ip vbp tail dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X351 a_21211_n2817# a_21036_n2791# a_21390_n2791# dvss.t157 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X352 tail vbp dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X353 a_17913_n2241# a_17747_n2241# dvss.t173 dvss.t172 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X354 dvdd.t3 a_20689_n2549# a_20579_n2425# dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X355 dvdd_ip standby_ip dvdd.t150 dvdd.t149 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X356 a_20567_n1869# a_20121_n2241# a_20471_n1869# dvss.t181 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X357 dvdd.t176 dvss.t114 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X358 dvss.t105 a_19003_n2817# a_19567_n2791# dvss.t104 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X359 a_18481_n2273# a_18263_n1869# dvss.t132 dvss.t131 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X360 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X361 dvss_ip vn vn dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X362 a_2130_n18852# a_24530_n19018# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X363 dvss.t130 x7.x2.Qb1 a_17747_n2791# dvss.t129 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X364 dvdd.t177 dvss.t115 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X365 avss.t28 avdd.t17 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X366 avss.t23 standby_ip x4.out_b.t1 avss.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X367 icnode vg2.t8 avss_ip.t18 avss_ip.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X368 avdd_ip.t15 vbreg xout.t14 avdd_ip.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X369 a_21211_n1943# a_21036_n1869# a_21390_n1881# dvss.t197 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X370 a_15960_n2791# x7.x2.Qb1 dvss.t128 dvss.t127 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X371 a_11526_n12394# icnode a_8268_n12482# avss_ip.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X372 avss_ip.t15 avss_ip.t16 avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X373 dvss.t28 a_19003_n1943# a_19567_n2247# dvss.t27 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X374 xout.t13 vbreg avdd_ip.t14 avdd_ip.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X375 dvss.t156 a_4857_n1521# standby_ip dvss.t155 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X376 a_14009_n2404# standby_ip dvss.t192 dvss.t21 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X377 inv_in.t9 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X378 dvdd_ip vbp vbp dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X379 a_2132_n14594# a_18932_n14760# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X380 a_16620_n2791# a_15539_n2791# a_16273_n2549# dvdd.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X381 dvss.t120 x7.x1.Qb1 a_17747_n2241# dvss.t119 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X382 a_18263_n2791# a_17913_n2791# a_18168_n2791# dvdd.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X383 dvdd.t172 a_16795_n2817# a_17359_n2791# dvdd.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X384 a_2971_n1521# ena.t1 dvss.t199 dvss.t198 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X385 dvss.t50 standby_b a_20733_n2791# dvss.t49 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X386 a_15960_n1881# x7.x1.Qb1 dvss.t118 dvss.t117 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X387 a_14035_n2281# x7.stby_done_b dvss.t141 dvss.t21 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X388 a_20579_n2425# a_19955_n2791# a_20471_n2791# dvdd.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X389 a_21145_n2791# a_19955_n2791# a_21036_n2791# dvss.t167 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X390 dvdd.t112 a_16273_n2549# a_16163_n2425# dvdd.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X391 a_16151_n1869# a_15705_n2241# a_16055_n1869# dvss.t3 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X392 a_2130_n18852# xout.t2 avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X393 dvdd.t136 a_18828_n2791# a_19003_n2817# dvdd.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X394 a_16782_n2247# a_15705_n2241# a_16620_n1869# dvdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X395 x3.out_b.t1 ena_ip avss.t11 avss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X396 dvss.t38 a_14009_n2404# x7.clk_disable dvss.t21 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X397 avss.t29 avdd.t16 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X398 dvdd.t148 standby_ip dvdd_ip dvdd.t147 sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X399 a_18481_n2549# a_18263_n2791# dvss.t201 dvss.t200 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X400 a_18359_n2791# a_17913_n2791# a_18263_n2791# dvss.t158 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X401 avdd_ip.t1 x3.out_b.t7 avdd.t3 avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X402 a_18263_n1869# a_17747_n2241# a_18168_n1881# dvss.t171 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X403 dvss.t88 ena_ip a_20733_n1881# dvss.t87 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X404 x7.x2.x3.Q a_19003_n2817# dvss.t103 dvss.t102 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X405 xout.t12 vbreg avdd_ip.t13 avdd_ip.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X406 avss_ip.t58 avss_ip.t59 avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X407 x7.x1.x3.Q a_19003_n1943# dvdd.t28 dvdd.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X408 a_21036_n2791# a_20121_n2791# a_20689_n2549# dvss.t183 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X409 dvss.t48 standby_b dvss_ip dvss.t47 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X410 avdd_ip.t33 icnode sky130_fd_pr__cap_mim_m3_1 l=20 w=20
X411 a_21211_n1943# ena_ip dvdd.t67 dvdd.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X412 inv_in.t10 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X413 inv_in.t11 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X414 a_10620_n8006# a_24220_n8172# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X415 avdd_ip.t12 vbreg xout.t11 avdd_ip.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X416 a_2130_n21840# a_24530_n21674# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X417 inv_in.t12 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X418 a_10620_n8006# a_24220_n7840# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X419 avdd.t12 x3.out_b.t8 avdd_ip.t4 avdd.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X420 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X421 avss.t9 ena_ip x3.out_b.t0 avss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X422 a_2132_n16254# a_18932_n16420# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X423 a_16163_n2425# a_15539_n2791# a_16055_n2791# dvdd.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X424 tail vbp dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X425 a_8268_n12482# a_8268_n12482# avss_ip.t54 avss_ip.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X426 x7.x2.x3.Q a_19003_n2817# dvdd.t78 dvdd.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X427 dvss.t187 a_14009_n2701# a_14035_n2743# dvss.t82 sky130_fd_pr__nfet_01v8 ad=0.07665 pd=0.785 as=0.0441 ps=0.63 w=0.42 l=0.15
X428 x7.x2.x2.CLK a_15000_n2791# dvdd.t22 dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X429 dvdd_ip vbp dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X430 a_21390_n2791# standby_b dvss.t46 dvss.t45 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X431 dvss.t122 a_21211_n2817# a_21145_n2791# dvss.t121 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X432 vg1.t8 xin.t2 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X433 dvss_ip standby_b dvss.t44 dvss.t43 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X434 inv_in.t13 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X435 a_16729_n2791# a_15539_n2791# a_16620_n2791# dvss.t34 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X436 a_9120_n9346.t4 a_9120_n9346.t3 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X437 a_2130_n21176# a_24530_n21010# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X438 a_2132_n17914# vg1.t0 avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X439 a_15960_n1881# x7.x1.Qb1 dvdd.t88 dvdd.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X440 a_20121_n2791# a_19955_n2791# dvdd.t126 dvdd.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X441 dvdd.t92 a_21211_n2817# a_21198_n2425# dvdd.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X442 a_14357_n2743# dout_ip dout_filt dvdd.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X443 a_2971_n1521# ena.t2 dvdd.t40 dvdd.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X444 a_21390_n1881# ena_ip dvss.t86 dvss.t85 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X445 standby_b standby_ip dvdd.t146 dvdd.t145 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X446 dvss_ip ibias_ip ibias_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X447 avss_ip.t32 x3.out.t7 avss.t21 avss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X448 a_18828_n2791# a_17747_n2791# a_18481_n2549# dvdd.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X449 a_18168_n1881# x7.x1.Qb2 dvdd.t59 dvdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X450 dvdd.t178 dvss.t116 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X451 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X452 dvss.t161 a_21211_n1943# a_21145_n1869# dvss.t160 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X453 a_14285_n2281# ena_ip a_14285_n2079# dvdd.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X454 avdd_ip.t11 vbreg avdd_ip.t10 avdd_ip.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X455 a_2132_n16254# a_18932_n16088# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X456 a_20689_n2549# a_20471_n2791# dvdd.t75 dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X457 dvdd.t18 x7.ena_done_b a_15000_n1881# dvdd.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X458 dvdd.t45 standby_b a_14285_n2281# dvdd.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X459 dvdd.t139 a_18481_n2549# a_18371_n2425# dvdd.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X460 dvdd_ip vbp tail dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X461 xout.t10 vbreg avdd_ip.t8 avdd_ip.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X462 a_18990_n2247# a_17913_n2241# a_18828_n1869# dvdd.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X463 a_20689_n2273# a_20471_n1869# dvdd.t7 dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X464 dvss_ip ibias_ip dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X465 vg1.t9 xin.t1 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X466 avss.t17 x3.out.t8 avss_ip.t24 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X467 avss_ip.t42 avss_ip.t40 avss_ip.t41 avss_ip.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X468 a_2132_n17914# a_18932_n17748# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X469 a_2132_n14262# a_18932_n14428# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X470 a_21198_n2425# a_20121_n2791# a_21036_n2791# dvdd.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X471 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X472 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X473 dvss.t210 a_16795_n2817# a_16729_n2791# dvss.t209 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X474 inv_in.t14 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X475 dvdd_ip vbp dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X476 dvdd_ip standby_ip dvdd.t144 dvdd.t143 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X477 avss_ip.t66 vg2.t1 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X478 a_2132_n15922# a_18932_n16088# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X479 a_18371_n2425# standby_b dvdd.t43 dvdd.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X480 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X481 a_18371_n2425# a_17747_n2791# a_18263_n2791# dvdd.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X482 ibias_ip ibias_ip dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X483 dvss.t10 a_16795_n1943# a_16729_n1869# dvss.t9 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X484 dout.t0 dout_filt dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X485 a_2132_n14262# vg2.t0 avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
X486 dvdd.t11 a_16795_n1943# a_16782_n2247# dvdd.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X487 avdd_ip.t7 vbreg avdd_ip.t6 avdd_ip.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X488 xout.t26 avdd_ip.t3 sky130_fd_pr__diode_pd2nw_05v5 perim=1.8e+06 area=2.025e+11
X489 a_20471_n2791# a_19955_n2791# a_20376_n2791# dvss.t166 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X490 x7.x1.Qb1 a_17359_n2247# dvss.t138 dvss.t137 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X491 a_20471_n1869# a_20121_n2241# a_20376_n1881# dvdd.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X492 dvdd.t142 standby_ip dvdd_ip dvdd.t141 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X493 a_2130_n21508# a_24530_n21342# avss_ip.t2 sky130_fd_pr__res_xhigh_po_0p35 l=110
X494 a_10620_n7674# inv_in.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X495 dvdd.t26 a_19003_n1943# a_18990_n2247# dvdd.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X496 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X497 a_18168_n2791# x7.x2.Qb2 dvss.t134 dvss.t133 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X498 vrb.t1 vg2.t9 vbreg avss_ip.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X499 a_2132_n15922# a_18932_n15756# avss_ip.t3 sky130_fd_pr__res_xhigh_po_0p35 l=82
R0 dvss.n623 dvss.n622 844724
R1 dvss.n146 dvss.n145 148018
R2 dvss.n650 dvss.n17 121073
R3 dvss.n144 dvss.n44 20785.4
R4 dvss.n145 dvss.n144 13161.6
R5 dvss.n43 dvss.n42 10590.5
R6 dvss.n142 dvss.n40 8607.23
R7 dvss.n562 dvss.n546 8366.71
R8 dvss.n546 dvss.n92 8366.71
R9 dvss.n544 dvss.n92 8366.71
R10 dvss.n562 dvss.n544 8366.71
R11 dvss.n613 dvss.n612 5881.35
R12 dvss.n88 dvss.n40 5784.65
R13 dvss.n624 dvss.n31 5227.07
R14 dvss.n32 dvss.n31 5083.5
R15 dvss.n612 dvss.n44 4954.5
R16 dvss.n229 dvss.n227 4604.94
R17 dvss.n603 dvss.n44 4392.82
R18 dvss.n101 dvss.n93 4247.09
R19 dvss.n541 dvss.n93 4247.09
R20 dvss.n101 dvss.n94 4247.09
R21 dvss.n541 dvss.n94 4247.09
R22 dvss.n213 dvss.n206 4247.09
R23 dvss.n218 dvss.n206 4247.09
R24 dvss.n213 dvss.n207 4247.09
R25 dvss.n218 dvss.n207 4247.09
R26 dvss.n623 dvss.n32 3898.89
R27 dvss.n622 dvss.n621 3764.56
R28 dvss.n625 dvss.n624 3697.38
R29 dvss.n227 dvss.n90 3234.36
R30 dvss.n29 dvss.n15 2798.56
R31 dvss.n653 dvss.n15 2798.56
R32 dvss.n29 dvss.n16 2798.56
R33 dvss.n653 dvss.n16 2798.56
R34 dvss.n589 dvss.n55 2798.56
R35 dvss.n56 dvss.n55 2798.56
R36 dvss.n589 dvss.n60 2798.56
R37 dvss.n60 dvss.n56 2798.56
R38 dvss.n543 dvss.n542 2575.49
R39 dvss.n624 dvss.n623 2562.64
R40 dvss.n613 dvss.n43 2543.9
R41 dvss.n233 dvss.n83 2397.52
R42 dvss.n303 dvss.n302 2387.64
R43 dvss.n436 dvss.n146 2316.35
R44 dvss.n143 dvss.n142 2162.81
R45 dvss.n566 dvss.n90 2000.34
R46 dvss.n649 dvss.n18 1686.66
R47 dvss.n304 dvss.n303 1680.95
R48 dvss.n630 dvss.n626 1407.97
R49 dvss.n636 dvss.n626 1407.97
R50 dvss.n636 dvss.n627 1407.97
R51 dvss.n586 dvss.n62 1407.97
R52 dvss.n70 dvss.n62 1407.97
R53 dvss.n586 dvss.n63 1407.97
R54 dvss.n70 dvss.n63 1407.97
R55 dvss.n34 dvss.n32 1313.59
R56 dvss.n681 dvss.n0 1212.38
R57 dvss.n588 dvss.n61 1202.51
R58 dvss.n220 dvss.n7 1198.25
R59 dvss.n302 dvss.n301 1198.25
R60 dvss.n289 dvss.n235 1198.25
R61 dvss.n518 dvss.n109 1198.25
R62 dvss.n478 dvss.n126 1198.25
R63 dvss.n438 dvss.n437 1198.25
R64 dvss.n435 dvss.n434 1198.25
R65 dvss.n209 dvss.n164 1198.25
R66 dvss.n210 dvss.n181 1198.25
R67 dvss.n315 dvss.n200 1198.25
R68 dvss.n305 dvss.n304 1198.25
R69 dvss.n639 dvss.n638 1198.25
R70 dvss.n73 dvss.n72 1198.25
R71 dvss.n651 dvss.n650 1184.03
R72 dvss.n681 dvss.n680 1175.19
R73 dvss.n615 dvss.n35 1127.15
R74 dvss.n42 dvss.n41 1064.88
R75 dvss.t17 dvss.t111 935.78
R76 dvss.t80 dvss.t172 935.78
R77 dvss.t117 dvss.t40 935.78
R78 dvss.n574 dvss.n85 927.908
R79 dvss.n145 dvss.n49 900.194
R80 dvss.n620 dvss.n35 884.347
R81 dvss.n554 dvss.n553 784.03
R82 dvss.n561 dvss.n560 783.962
R83 dvss.n553 dvss.n552 783.75
R84 dvss.n561 dvss.n551 783.683
R85 dvss.n235 dvss.t0 748.625
R86 dvss.n614 dvss.n613 720.655
R87 dvss.t168 dvss.t142 717.851
R88 dvss.t188 dvss.t133 717.851
R89 dvss.t162 dvss.t164 689.909
R90 dvss.t164 dvss.t197 689.909
R91 dvss.t27 dvss.t29 689.909
R92 dvss.t29 dvss.t150 689.909
R93 dvss.t13 dvss.t11 689.909
R94 dvss.t179 dvss.t13 689.909
R95 dvss.n211 dvss.t35 655.918
R96 dvss.n652 dvss.n651 639.12
R97 dvss.n598 dvss.n597 626.816
R98 dvss.n30 dvss.t89 618.75
R99 dvss.n652 dvss.t89 618.75
R100 dvss.t153 dvss.t181 609.174
R101 dvss.t33 dvss.t152 609.174
R102 dvss.t3 dvss.t101 609.174
R103 dvss.n84 dvss.n81 585
R104 dvss.n84 dvss.n61 585
R105 dvss.n605 dvss.n604 585
R106 dvss.n604 dvss.n603 585
R107 dvss.n229 dvss.n107 585
R108 dvss.n229 dvss.n228 585
R109 dvss.n230 dvss.n83 585
R110 dvss.n91 dvss.n83 585
R111 dvss.n571 dvss.n570 585
R112 dvss.n572 dvss.n571 585
R113 dvss.n569 dvss.n88 585
R114 dvss.n88 dvss.n86 585
R115 dvss.t23 dvss.n200 574.28
R116 dvss.n437 dvss.t175 554.129
R117 dvss.n126 dvss.t75 554.129
R118 dvss.t137 dvss.n109 554.129
R119 dvss.t85 dvss.t160 546.789
R120 dvss.t91 dvss.t31 546.789
R121 dvss.t9 dvss.t93 546.789
R122 dvss.t123 dvss.t125 529.24
R123 dvss.t157 dvss.t123 529.24
R124 dvss.t102 dvss.t104 529.24
R125 dvss.t180 dvss.t102 529.24
R126 dvss.t211 dvss.t213 529.24
R127 dvss.t146 dvss.t211 529.24
R128 dvss.t5 dvss.t87 484.404
R129 dvss.t131 dvss.t95 484.404
R130 dvss.t97 dvss.t139 484.404
R131 dvss.t184 dvss.t2 467.307
R132 dvss.t158 dvss.t186 467.307
R133 dvss.t203 dvss.t147 467.307
R134 dvss.n615 dvss.n39 467.033
R135 dvss.t0 dvss.t19 447.707
R136 dvss.n303 dvss.n220 426.382
R137 dvss.n435 dvss.t25 425.08
R138 dvss.t148 dvss.n209 425.08
R139 dvss.t177 dvss.n210 425.08
R140 dvss.t121 dvss.t45 419.45
R141 dvss.t106 dvss.t59 419.45
R142 dvss.t209 dvss.t61 419.45
R143 dvss.n638 dvss.n637 419.18
R144 dvss.n597 dvss.n50 404.022
R145 dvss.t113 dvss.t182 400
R146 dvss.t174 dvss.t151 400
R147 dvss.t4 dvss.t42 400
R148 dvss.n630 dvss.n629 390.825
R149 dvss.t49 dvss.t99 371.594
R150 dvss.t67 dvss.t200 371.594
R151 dvss.t71 dvss.t108 371.594
R152 dvss.n651 dvss.t204 366.435
R153 dvss.t182 dvss.t5 363.303
R154 dvss.t151 dvss.t131 363.303
R155 dvss.t139 dvss.t4 363.303
R156 dvss.t175 dvss.t162 355.964
R157 dvss.t75 dvss.t27 355.964
R158 dvss.t11 dvss.t137 355.964
R159 dvss.t160 dvss.t113 352.295
R160 dvss.t181 dvss.t110 352.295
R161 dvss.t31 dvss.t174 352.295
R162 dvss.t152 dvss.t171 352.295
R163 dvss.t42 dvss.t9 352.295
R164 dvss.t110 dvss.t17 348.625
R165 dvss.t171 dvss.t80 348.625
R166 dvss.t39 dvss.t117 348.625
R167 dvss.n637 dvss.n625 344.228
R168 dvss.t144 dvss.t23 343.442
R169 dvss.n233 dvss.n229 335.039
R170 dvss.t197 dvss.t85 333.945
R171 dvss.t150 dvss.t91 333.945
R172 dvss.t93 dvss.t179 333.945
R173 dvss.n85 dvss.n84 331.606
R174 dvss.n228 dvss.t39 326.606
R175 dvss.n615 dvss.n40 310.599
R176 dvss.n41 dvss.n35 308.933
R177 dvss.n437 dvss.n436 308.257
R178 dvss.t111 dvss.t78 308.257
R179 dvss.t172 dvss.t119 308.257
R180 dvss.n638 dvss 308.139
R181 dvss.n283 dvss.t118 307.536
R182 dvss.n512 dvss.t81 307.536
R183 dvss.n472 dvss.t18 307.536
R184 dvss.n161 dvss.t143 307.536
R185 dvss.n178 dvss.t134 307.536
R186 dvss.n321 dvss.t128 307.536
R187 dvss.t183 dvss.t167 306.846
R188 dvss.t159 dvss.t191 306.846
R189 dvss.t202 dvss.t34 306.846
R190 dvss.n70 dvss.n69 292.5
R191 dvss.n71 dvss.n70 292.5
R192 dvss.n68 dvss.n63 292.5
R193 dvss.t154 dvss.n63 292.5
R194 dvss.n586 dvss.n585 292.5
R195 dvss.n587 dvss.n586 292.5
R196 dvss.n64 dvss.n62 292.5
R197 dvss.t154 dvss.n62 292.5
R198 dvss.n633 dvss.n627 292.5
R199 dvss.n636 dvss.n635 292.5
R200 dvss.n637 dvss.n636 292.5
R201 dvss.n628 dvss.n626 292.5
R202 dvss.t185 dvss.n626 292.5
R203 dvss.n631 dvss.n630 292.5
R204 dvss.t83 dvss 289.909
R205 dvss.t99 dvss.t183 278.695
R206 dvss.t200 dvss.t159 278.695
R207 dvss.t108 dvss.t202 278.695
R208 dvss.n217 dvss.n215 276.286
R209 dvss dvss.n126 275.229
R210 dvss dvss.n109 275.229
R211 dvss.n235 dvss 275.229
R212 dvss.n302 dvss 275.229
R213 dvss.t193 dvss.n0 273.678
R214 dvss.n542 dvss.t193 273.678
R215 dvss.t125 dvss.t25 273.065
R216 dvss.t104 dvss.t148 273.065
R217 dvss.t213 dvss.t177 273.065
R218 dvss.t167 dvss.t121 270.25
R219 dvss.t166 dvss.t184 270.25
R220 dvss.t191 dvss.t106 270.25
R221 dvss.t190 dvss.t158 270.25
R222 dvss.t34 dvss.t209 270.25
R223 dvss.t142 dvss.t166 267.435
R224 dvss.t133 dvss.t190 267.435
R225 dvss.t37 dvss.t127 267.435
R226 dvss.t87 dvss.t153 264.221
R227 dvss.t95 dvss.t33 264.221
R228 dvss.t101 dvss.t97 264.221
R229 dvss.t19 dvss.t83 264.221
R230 dvss.n611 dvss.n45 258.5
R231 dvss.t45 dvss.t157 256.175
R232 dvss.t59 dvss.t180 256.175
R233 dvss.t61 dvss.t146 256.175
R234 dvss.n543 dvss.t51 255.168
R235 dvss.n256 dvss.t14 246.817
R236 dvss.n485 dvss.t30 246.817
R237 dvss.n445 dvss.t165 246.817
R238 dvss.n151 dvss.t124 246.817
R239 dvss.n386 dvss.t103 246.817
R240 dvss.n347 dvss.t212 246.817
R241 dvss.t198 dvss.t204 244.291
R242 dvss.t78 dvss 238.532
R243 dvss.t119 dvss 238.532
R244 dvss dvss.t15 238.532
R245 dvss.n436 dvss.n435 236.469
R246 dvss.t135 dvss.t168 236.469
R247 dvss.t129 dvss.t188 236.469
R248 dvss.t35 dvss.t7 236.469
R249 dvss.n61 dvss.n42 236.023
R250 dvss.n588 dvss.n587 230.855
R251 dvss.n325 dvss.t207 229.185
R252 dvss.n522 dvss.n521 227.357
R253 dvss.n97 dvss.t194 219.8
R254 dvss.n540 dvss.n95 217.329
R255 dvss.n215 dvss.n214 217.225
R256 dvss.n249 dvss.n248 214.742
R257 dvss.n123 dvss.n122 214.742
R258 dvss.n140 dvss.n139 214.742
R259 dvss.n150 dvss.n149 214.742
R260 dvss.n392 dvss.n166 214.742
R261 dvss.n353 dvss.n183 214.742
R262 dvss.n571 dvss.n87 213.325
R263 dvss.n209 dvss 211.132
R264 dvss.n210 dvss 211.132
R265 dvss dvss.n200 211.132
R266 dvss.n304 dvss 211.132
R267 dvss.n263 dvss.n245 209.254
R268 dvss.n492 dvss.n119 209.254
R269 dvss.n452 dvss.n136 209.254
R270 dvss.n154 dvss.n153 209.254
R271 dvss.n172 dvss.n171 209.254
R272 dvss.n189 dvss.n188 209.254
R273 dvss.t51 dvss.t55 208.894
R274 dvss.t55 dvss.t63 208.894
R275 dvss.t63 dvss.t43 208.894
R276 dvss.t43 dvss.t47 208.894
R277 dvss.t69 dvss.t73 208.894
R278 dvss.t73 dvss.t53 208.894
R279 dvss.t57 dvss.t65 208.894
R280 dvss.n526 dvss.n525 203.619
R281 dvss.t2 dvss.t49 202.688
R282 dvss.t186 dvss.t67 202.688
R283 dvss.t147 dvss.t71 202.688
R284 dvss.t84 dvss.t144 202.688
R285 dvss.n666 dvss.n6 202.067
R286 dvss.n604 dvss.n45 202.048
R287 dvss.n3 dvss.n2 200.516
R288 dvss.n237 dvss.n236 199.739
R289 dvss.n271 dvss.n270 199.739
R290 dvss.n111 dvss.n110 199.739
R291 dvss.n500 dvss.n499 199.739
R292 dvss.n128 dvss.n127 199.739
R293 dvss.n460 dvss.n459 199.739
R294 dvss.n412 dvss.n158 199.739
R295 dvss.n399 dvss.n163 199.739
R296 dvss.n373 dvss.n175 199.739
R297 dvss.n360 dvss.n180 199.739
R298 dvss.n334 dvss.n192 199.739
R299 dvss.n199 dvss.n198 199.739
R300 dvss.n24 dvss.n23 199.739
R301 dvss.n75 dvss.n74 199.739
R302 dvss.n540 dvss.n539 198.024
R303 dvss.n587 dvss.t195 187.785
R304 dvss.n295 dvss.n294 185
R305 dvss.n205 dvss.n204 185
R306 dvss.n679 dvss.n678 185
R307 dvss dvss.t135 182.982
R308 dvss dvss.t129 182.982
R309 dvss.n28 dvss.n12 181.835
R310 dvss.n28 dvss.n27 181.835
R311 dvss.n58 dvss.n57 181.835
R312 dvss.n59 dvss.n58 181.835
R313 dvss.n629 dvss.n627 174.962
R314 dvss.n212 dvss.t37 166.091
R315 dvss.n234 dvss.t40 161.469
R316 dvss.n31 dvss.n30 155.325
R317 dvss.n219 dvss.t84 154.831
R318 dvss.n95 dvss.n93 148.029
R319 dvss.t15 dvss.n234 146.79
R320 dvss.n218 dvss.n217 146.25
R321 dvss.n219 dvss.n218 146.25
R322 dvss.n214 dvss.n213 146.25
R323 dvss.n213 dvss.n212 146.25
R324 dvss.n96 dvss.n94 146.25
R325 dvss.n94 dvss.t193 146.25
R326 dvss.n93 dvss.t193 146.25
R327 dvss.n102 dvss.n95 143.809
R328 dvss.n577 dvss.n81 143.196
R329 dvss.t155 dvss 141.269
R330 dvss.t7 dvss.t206 140.756
R331 dvss dvss.t82 140.144
R332 dvss.n545 dvss.n86 129.567
R333 dvss.n574 dvss.n83 128.583
R334 dvss.n217 dvss.n216 127.487
R335 dvss.n72 dvss.n33 122.319
R336 dvss.t65 dvss.n572 120.312
R337 dvss.n58 dvss.n56 117.001
R338 dvss.n56 dvss.n33 117.001
R339 dvss.n60 dvss.n59 117.001
R340 dvss.t195 dvss.n60 117.001
R341 dvss.n590 dvss.n589 117.001
R342 dvss.n589 dvss.n588 117.001
R343 dvss.n57 dvss.n55 117.001
R344 dvss.t195 dvss.n55 117.001
R345 dvss.n654 dvss.n653 117.001
R346 dvss.n653 dvss.n652 117.001
R347 dvss.n16 dvss.n12 117.001
R348 dvss.t89 dvss.n16 117.001
R349 dvss.n29 dvss.n28 117.001
R350 dvss.n30 dvss.n29 117.001
R351 dvss.n27 dvss.n15 117.001
R352 dvss.t89 dvss.n15 117.001
R353 dvss.n573 dvss.t53 113.703
R354 dvss.n232 dvss.n231 108.201
R355 dvss.n622 dvss.n33 105.091
R356 dvss.n212 dvss.t203 104.159
R357 dvss.n654 dvss.n13 102.025
R358 dvss.n655 dvss.n654 102.025
R359 dvss.n590 dvss.n52 102.025
R360 dvss.n590 dvss.n54 102.025
R361 dvss.n648 dvss.n19 101.874
R362 dvss.t47 dvss.n91 101.803
R363 dvss.n245 dvss.t94 100.001
R364 dvss.n119 dvss.t92 100.001
R365 dvss.n136 dvss.t86 100.001
R366 dvss.n153 dvss.t46 100.001
R367 dvss.n171 dvss.t60 100.001
R368 dvss.n188 dvss.t62 100.001
R369 dvss.n599 dvss.n598 98.4337
R370 dvss.n573 dvss.t57 95.1928
R371 dvss.n631 dvss.n628 91.4829
R372 dvss.n69 dvss.n64 91.4829
R373 dvss.n545 dvss.n43 85.938
R374 dvss.n53 dvss.t196 83.7183
R375 dvss.n646 dvss.t90 83.7183
R376 dvss.n142 dvss.n45 81.509
R377 dvss.n629 dvss.t185 81.1932
R378 dvss dvss.t198 80.5052
R379 dvss.n655 dvss.n12 79.8123
R380 dvss.n27 dvss.n13 79.8123
R381 dvss.n59 dvss.n52 79.8123
R382 dvss.n57 dvss.n54 79.8123
R383 dvss.n617 dvss.n616 73.2369
R384 dvss.n616 dvss.n615 73.1255
R385 dvss.n615 dvss.n614 73.1255
R386 dvss.n294 dvss.t1 72.8576
R387 dvss.n270 dvss.t98 72.8576
R388 dvss.n499 dvss.t96 72.8576
R389 dvss.n459 dvss.t88 72.8576
R390 dvss.n204 dvss.t24 72.8576
R391 dvss.n158 dvss.t50 72.8576
R392 dvss.n175 dvss.t68 72.8576
R393 dvss.n192 dvss.t72 72.8576
R394 dvss.n41 dvss.n39 72.01
R395 dvss.n521 dvss.n107 71.4371
R396 dvss.n245 dvss.t10 70.0005
R397 dvss.n119 dvss.t32 70.0005
R398 dvss.n136 dvss.t161 70.0005
R399 dvss.n153 dvss.t122 70.0005
R400 dvss.n171 dvss.t107 70.0005
R401 dvss.n188 dvss.t210 70.0005
R402 dvss.n69 dvss.n68 69.6045
R403 dvss.n635 dvss.n628 69.0306
R404 dvss dvss.t154 68.912
R405 dvss.n208 dvss.n196 68.8106
R406 dvss dvss.n219 67.5629
R407 dvss.n585 dvss.n64 66.3131
R408 dvss.n632 dvss.n631 65.475
R409 dvss.n527 dvss.n526 64.5768
R410 dvss.n564 dvss.t69 63.462
R411 dvss.t127 dvss.n211 61.9327
R412 dvss.n270 dvss.t140 60.5809
R413 dvss.n499 dvss.t132 60.5809
R414 dvss.n459 dvss.t6 60.5809
R415 dvss.n158 dvss.t100 60.5809
R416 dvss.n175 dvss.t201 60.5809
R417 dvss.n192 dvss.t109 60.5809
R418 dvss.n294 dvss.t20 58.5719
R419 dvss.n204 dvss.t145 58.5719
R420 dvss.n619 dvss.n617 57.4606
R421 dvss.n599 dvss.n49 57.2559
R422 dvss.n248 dvss.t12 57.1434
R423 dvss.n122 dvss.t28 57.1434
R424 dvss.n139 dvss.t163 57.1434
R425 dvss.n149 dvss.t126 57.1434
R426 dvss.n166 dvss.t105 57.1434
R427 dvss.n183 dvss.t214 57.1434
R428 dvss.n614 dvss.n42 54.0496
R429 dvss.n678 dvss.t187 52.8576
R430 dvss.n678 dvss.t208 51.4291
R431 dvss.n576 dvss.n575 45.2502
R432 dvss.n85 dvss.n39 44.978
R433 dvss.t206 dvss 42.227
R434 dvss.n216 dvss.n207 41.7862
R435 dvss.t206 dvss.n207 41.7862
R436 dvss.n215 dvss.n206 41.7862
R437 dvss.t206 dvss.n206 41.7862
R438 dvss.n541 dvss.n540 41.7862
R439 dvss.n542 dvss.n541 41.7862
R440 dvss.n102 dvss.n101 41.7862
R441 dvss.n101 dvss.n0 41.7862
R442 dvss.n554 dvss.n546 41.7862
R443 dvss.n546 dvss.n545 41.7862
R444 dvss.n552 dvss.n544 41.7862
R445 dvss.n544 dvss.n543 41.7862
R446 dvss.n231 dvss.n230 40.2432
R447 dvss.n677 dvss.n676 40.0735
R448 dvss.n236 dvss.t41 38.5719
R449 dvss.n236 dvss.t16 38.5719
R450 dvss.n110 dvss.t173 38.5719
R451 dvss.n110 dvss.t120 38.5719
R452 dvss.n127 dvss.t112 38.5719
R453 dvss.n127 dvss.t79 38.5719
R454 dvss.n163 dvss.t169 38.5719
R455 dvss.n163 dvss.t136 38.5719
R456 dvss.n180 dvss.t189 38.5719
R457 dvss.n180 dvss.t130 38.5719
R458 dvss.n198 dvss.t36 38.5719
R459 dvss.n198 dvss.t8 38.5719
R460 dvss.n634 dvss.n633 37.6894
R461 dvss.n584 dvss.n65 37.4862
R462 dvss.n611 dvss.n40 36.1883
R463 dvss.t154 dvss.t195 36.179
R464 dvss.n72 dvss.n71 36.179
R465 dvss.n6 dvss.t22 36.0005
R466 dvss.n565 dvss.n563 35.6976
R467 dvss.n537 dvss.n536 35.5421
R468 dvss.n670 dvss.n5 34.6358
R469 dvss.n671 dvss.n670 34.6358
R470 dvss.n672 dvss.n671 34.6358
R471 dvss.n300 dvss.n225 34.6358
R472 dvss.n293 dvss.n226 34.6358
R473 dvss.n276 dvss.n241 34.6358
R474 dvss.n277 dvss.n276 34.6358
R475 dvss.n278 dvss.n277 34.6358
R476 dvss.n278 dvss.n239 34.6358
R477 dvss.n282 dvss.n239 34.6358
R478 dvss.n264 dvss.n243 34.6358
R479 dvss.n268 dvss.n243 34.6358
R480 dvss.n269 dvss.n268 34.6358
R481 dvss.n272 dvss.n269 34.6358
R482 dvss.n251 dvss.n108 34.6358
R483 dvss.n255 dvss.n254 34.6358
R484 dvss.n257 dvss.n255 34.6358
R485 dvss.n261 dvss.n246 34.6358
R486 dvss.n262 dvss.n261 34.6358
R487 dvss.n505 dvss.n115 34.6358
R488 dvss.n506 dvss.n505 34.6358
R489 dvss.n507 dvss.n506 34.6358
R490 dvss.n507 dvss.n113 34.6358
R491 dvss.n511 dvss.n113 34.6358
R492 dvss.n493 dvss.n117 34.6358
R493 dvss.n497 dvss.n117 34.6358
R494 dvss.n498 dvss.n497 34.6358
R495 dvss.n501 dvss.n498 34.6358
R496 dvss.n480 dvss.n479 34.6358
R497 dvss.n484 dvss.n483 34.6358
R498 dvss.n486 dvss.n484 34.6358
R499 dvss.n490 dvss.n120 34.6358
R500 dvss.n491 dvss.n490 34.6358
R501 dvss.n465 dvss.n132 34.6358
R502 dvss.n466 dvss.n465 34.6358
R503 dvss.n467 dvss.n466 34.6358
R504 dvss.n467 dvss.n130 34.6358
R505 dvss.n471 dvss.n130 34.6358
R506 dvss.n453 dvss.n134 34.6358
R507 dvss.n457 dvss.n134 34.6358
R508 dvss.n458 dvss.n457 34.6358
R509 dvss.n461 dvss.n458 34.6358
R510 dvss.n440 dvss.n439 34.6358
R511 dvss.n444 dvss.n443 34.6358
R512 dvss.n446 dvss.n444 34.6358
R513 dvss.n450 dvss.n137 34.6358
R514 dvss.n451 dvss.n450 34.6358
R515 dvss.n433 dvss.n147 34.6358
R516 dvss.n429 dvss.n428 34.6358
R517 dvss.n428 dvss.n427 34.6358
R518 dvss.n424 dvss.n423 34.6358
R519 dvss.n423 dvss.n422 34.6358
R520 dvss.n419 dvss.n418 34.6358
R521 dvss.n418 dvss.n417 34.6358
R522 dvss.n417 dvss.n156 34.6358
R523 dvss.n413 dvss.n156 34.6358
R524 dvss.n411 dvss.n410 34.6358
R525 dvss.n410 dvss.n159 34.6358
R526 dvss.n406 dvss.n159 34.6358
R527 dvss.n406 dvss.n405 34.6358
R528 dvss.n405 dvss.n404 34.6358
R529 dvss.n394 dvss.n393 34.6358
R530 dvss.n391 dvss.n167 34.6358
R531 dvss.n387 dvss.n167 34.6358
R532 dvss.n385 dvss.n384 34.6358
R533 dvss.n384 dvss.n169 34.6358
R534 dvss.n380 dvss.n379 34.6358
R535 dvss.n379 dvss.n378 34.6358
R536 dvss.n378 dvss.n173 34.6358
R537 dvss.n374 dvss.n173 34.6358
R538 dvss.n372 dvss.n371 34.6358
R539 dvss.n371 dvss.n176 34.6358
R540 dvss.n367 dvss.n176 34.6358
R541 dvss.n367 dvss.n366 34.6358
R542 dvss.n366 dvss.n365 34.6358
R543 dvss.n355 dvss.n354 34.6358
R544 dvss.n352 dvss.n184 34.6358
R545 dvss.n348 dvss.n184 34.6358
R546 dvss.n346 dvss.n345 34.6358
R547 dvss.n345 dvss.n186 34.6358
R548 dvss.n341 dvss.n340 34.6358
R549 dvss.n340 dvss.n190 34.6358
R550 dvss.n336 dvss.n190 34.6358
R551 dvss.n336 dvss.n335 34.6358
R552 dvss.n333 dvss.n193 34.6358
R553 dvss.n329 dvss.n193 34.6358
R554 dvss.n329 dvss.n328 34.6358
R555 dvss.n328 dvss.n195 34.6358
R556 dvss.n322 dvss.n195 34.6358
R557 dvss.n314 dvss.n202 34.6358
R558 dvss.n309 dvss.n308 34.6358
R559 dvss.n23 dvss.t199 33.462
R560 dvss.n23 dvss.t205 33.462
R561 dvss.n74 dvss.t170 33.462
R562 dvss.n74 dvss.t156 33.462
R563 dvss.n2 dvss.t38 33.2313
R564 dvss.n24 dvss.n21 31.5123
R565 dvss.n254 dvss.n249 31.2476
R566 dvss.n483 dvss.n123 31.2476
R567 dvss.n443 dvss.n140 31.2476
R568 dvss.n429 dvss.n150 31.2476
R569 dvss.n392 dvss.n391 31.2476
R570 dvss.n353 dvss.n352 31.2476
R571 dvss.t21 dvss.t82 30.4092
R572 dvss dvss.n681 30.4092
R573 dvss.n616 dvss.n37 30.2484
R574 dvss.n284 dvss.n283 29.7417
R575 dvss.n513 dvss.n512 29.7417
R576 dvss.n473 dvss.n472 29.7417
R577 dvss.n400 dvss.n161 29.7417
R578 dvss.n361 dvss.n178 29.7417
R579 dvss.n321 dvss.n320 29.7417
R580 dvss.n80 dvss.n37 28.5338
R581 dvss.n538 dvss.n99 28.3255
R582 dvss.n527 dvss.n100 27.9866
R583 dvss.n256 dvss.n246 27.8593
R584 dvss.n485 dvss.n120 27.8593
R585 dvss.n445 dvss.n137 27.8593
R586 dvss.n424 dvss.n151 27.8593
R587 dvss.n386 dvss.n385 27.8593
R588 dvss.n347 dvss.n346 27.8593
R589 dvss.n676 dvss.n3 25.977
R590 dvss.n228 dvss.t3 25.6886
R591 dvss.n248 dvss.t138 25.4291
R592 dvss.n122 dvss.t76 25.4291
R593 dvss.n139 dvss.t176 25.4291
R594 dvss.n149 dvss.t26 25.4291
R595 dvss.n166 dvss.t149 25.4291
R596 dvss.n183 dvss.t178 25.4291
R597 dvss.n2 dvss.t141 24.9236
R598 dvss.n6 dvss.t192 24.9236
R599 dvss.n562 dvss.n561 24.3755
R600 dvss.n563 dvss.n562 24.3755
R601 dvss.n553 dvss.n92 24.3755
R602 dvss.n563 dvss.n92 24.3755
R603 dvss.n296 dvss.n225 23.7737
R604 dvss.n310 dvss.n309 23.7737
R605 dvss.n665 dvss.n7 23.7181
R606 dvss.n301 dvss.n300 23.7181
R607 dvss.n289 dvss.n226 23.7181
R608 dvss.n289 dvss.n288 23.7181
R609 dvss.n518 dvss.n108 23.7181
R610 dvss.n518 dvss.n517 23.7181
R611 dvss.n479 dvss.n478 23.7181
R612 dvss.n478 dvss.n477 23.7181
R613 dvss.n439 dvss.n438 23.7181
R614 dvss.n434 dvss.n433 23.7181
R615 dvss.n398 dvss.n164 23.7181
R616 dvss.n394 dvss.n164 23.7181
R617 dvss.n359 dvss.n181 23.7181
R618 dvss.n355 dvss.n181 23.7181
R619 dvss.n316 dvss.n315 23.7181
R620 dvss.n315 dvss.n314 23.7181
R621 dvss.n308 dvss.n305 23.7181
R622 dvss.n639 dvss.n26 23.7181
R623 dvss.n76 dvss.n73 23.7181
R624 dvss.n666 dvss.n5 22.9652
R625 dvss.n284 dvss.n237 22.9652
R626 dvss.n513 dvss.n111 22.9652
R627 dvss.n473 dvss.n128 22.9652
R628 dvss.n400 dvss.n399 22.9652
R629 dvss.n361 dvss.n360 22.9652
R630 dvss.n320 dvss.n199 22.9652
R631 dvss.n537 dvss.n533 22.1054
R632 dvss.n232 dvss.n107 21.7695
R633 dvss.n98 dvss.n97 21.753
R634 dvss.n666 dvss.n665 21.4593
R635 dvss.n288 dvss.n237 21.4593
R636 dvss.n517 dvss.n111 21.4593
R637 dvss.n477 dvss.n128 21.4593
R638 dvss.n399 dvss.n398 21.4593
R639 dvss.n360 dvss.n359 21.4593
R640 dvss.n316 dvss.n199 21.4593
R641 dvss.n680 dvss.n679 21.4265
R642 dvss.n552 dvss.t52 21.1687
R643 dvss.n554 dvss.t66 21.1687
R644 dvss.n220 dvss.t21 21.1543
R645 dvss.n295 dvss.n293 20.9718
R646 dvss.n205 dvss.n202 20.9718
R647 dvss.n576 dvss.n37 20.1009
R648 dvss.n617 dvss.n36 20.0732
R649 dvss.n528 dvss.n527 18.7867
R650 dvss.n559 dvss.n555 18.4515
R651 dvss.n558 dvss.n556 18.4515
R652 dvss.n549 dvss.n548 18.4515
R653 dvss.n550 dvss.n547 18.4515
R654 dvss.n672 dvss.n3 18.4476
R655 dvss.n263 dvss.n262 17.6946
R656 dvss.n492 dvss.n491 17.6946
R657 dvss.n452 dvss.n451 17.6946
R658 dvss.n422 dvss.n154 17.6946
R659 dvss.n172 dvss.n169 17.6946
R660 dvss.n189 dvss.n186 17.6946
R661 dvss.t185 dvss.n625 16.6567
R662 dvss dvss.n24 15.0593
R663 dvss dvss.n75 15.0593
R664 dvss.n283 dvss.n282 14.6829
R665 dvss.n512 dvss.n511 14.6829
R666 dvss.n472 dvss.n471 14.6829
R667 dvss.n404 dvss.n161 14.6829
R668 dvss.n365 dvss.n178 14.6829
R669 dvss.n322 dvss.n321 14.6829
R670 dvss.n594 dvss.n593 14.3573
R671 dvss.n570 dvss.n568 13.8612
R672 dvss.n71 dvss.t155 13.7828
R673 dvss.n99 dvss.n98 13.2836
R674 dvss.n606 dvss.n47 13.0628
R675 dvss.n610 dvss.n609 12.2414
R676 dvss.n97 dvss.n95 11.7338
R677 dvss.n581 dvss.n54 10.5081
R678 dvss.n597 dvss.n596 10.2484
R679 dvss.n592 dvss.n52 10.2179
R680 dvss.n656 dvss.n655 10.1264
R681 dvss.n649 dvss.n648 9.79535
R682 dvss.n582 dvss.n79 9.76662
R683 dvss.n596 dvss.n38 9.49353
R684 dvss.n80 dvss.n79 9.30109
R685 dvss.n306 dvss.n305 9.3005
R686 dvss.n324 dvss.n195 9.3005
R687 dvss.n323 dvss.n322 9.3005
R688 dvss.n321 dvss.n197 9.3005
R689 dvss.n320 dvss.n319 9.3005
R690 dvss.n318 dvss.n199 9.3005
R691 dvss.n317 dvss.n316 9.3005
R692 dvss.n315 dvss.n201 9.3005
R693 dvss.n314 dvss.n313 9.3005
R694 dvss.n312 dvss.n202 9.3005
R695 dvss.n311 dvss.n310 9.3005
R696 dvss.n309 dvss.n203 9.3005
R697 dvss.n308 dvss.n307 9.3005
R698 dvss.n434 dvss.n105 9.3005
R699 dvss.n433 dvss.n432 9.3005
R700 dvss.n431 dvss.n147 9.3005
R701 dvss.n430 dvss.n429 9.3005
R702 dvss.n428 dvss.n148 9.3005
R703 dvss.n427 dvss.n426 9.3005
R704 dvss.n425 dvss.n424 9.3005
R705 dvss.n423 dvss.n152 9.3005
R706 dvss.n422 dvss.n421 9.3005
R707 dvss.n420 dvss.n419 9.3005
R708 dvss.n418 dvss.n155 9.3005
R709 dvss.n417 dvss.n416 9.3005
R710 dvss.n415 dvss.n156 9.3005
R711 dvss.n414 dvss.n413 9.3005
R712 dvss.n411 dvss.n157 9.3005
R713 dvss.n410 dvss.n409 9.3005
R714 dvss.n408 dvss.n159 9.3005
R715 dvss.n407 dvss.n406 9.3005
R716 dvss.n405 dvss.n160 9.3005
R717 dvss.n404 dvss.n403 9.3005
R718 dvss.n402 dvss.n161 9.3005
R719 dvss.n401 dvss.n400 9.3005
R720 dvss.n399 dvss.n162 9.3005
R721 dvss.n398 dvss.n397 9.3005
R722 dvss.n396 dvss.n164 9.3005
R723 dvss.n395 dvss.n394 9.3005
R724 dvss.n393 dvss.n165 9.3005
R725 dvss.n391 dvss.n390 9.3005
R726 dvss.n389 dvss.n167 9.3005
R727 dvss.n388 dvss.n387 9.3005
R728 dvss.n385 dvss.n168 9.3005
R729 dvss.n384 dvss.n383 9.3005
R730 dvss.n382 dvss.n169 9.3005
R731 dvss.n381 dvss.n380 9.3005
R732 dvss.n379 dvss.n170 9.3005
R733 dvss.n378 dvss.n377 9.3005
R734 dvss.n376 dvss.n173 9.3005
R735 dvss.n375 dvss.n374 9.3005
R736 dvss.n372 dvss.n174 9.3005
R737 dvss.n371 dvss.n370 9.3005
R738 dvss.n369 dvss.n176 9.3005
R739 dvss.n368 dvss.n367 9.3005
R740 dvss.n366 dvss.n177 9.3005
R741 dvss.n365 dvss.n364 9.3005
R742 dvss.n363 dvss.n178 9.3005
R743 dvss.n362 dvss.n361 9.3005
R744 dvss.n360 dvss.n179 9.3005
R745 dvss.n359 dvss.n358 9.3005
R746 dvss.n357 dvss.n181 9.3005
R747 dvss.n356 dvss.n355 9.3005
R748 dvss.n354 dvss.n182 9.3005
R749 dvss.n352 dvss.n351 9.3005
R750 dvss.n350 dvss.n184 9.3005
R751 dvss.n349 dvss.n348 9.3005
R752 dvss.n346 dvss.n185 9.3005
R753 dvss.n345 dvss.n344 9.3005
R754 dvss.n343 dvss.n186 9.3005
R755 dvss.n342 dvss.n341 9.3005
R756 dvss.n340 dvss.n339 9.3005
R757 dvss.n338 dvss.n190 9.3005
R758 dvss.n337 dvss.n336 9.3005
R759 dvss.n335 dvss.n191 9.3005
R760 dvss.n333 dvss.n332 9.3005
R761 dvss.n331 dvss.n193 9.3005
R762 dvss.n330 dvss.n329 9.3005
R763 dvss.n328 dvss.n327 9.3005
R764 dvss.n438 dvss.n106 9.3005
R765 dvss.n439 dvss.n141 9.3005
R766 dvss.n441 dvss.n440 9.3005
R767 dvss.n443 dvss.n442 9.3005
R768 dvss.n444 dvss.n138 9.3005
R769 dvss.n447 dvss.n446 9.3005
R770 dvss.n448 dvss.n137 9.3005
R771 dvss.n450 dvss.n449 9.3005
R772 dvss.n451 dvss.n135 9.3005
R773 dvss.n454 dvss.n453 9.3005
R774 dvss.n455 dvss.n134 9.3005
R775 dvss.n457 dvss.n456 9.3005
R776 dvss.n458 dvss.n133 9.3005
R777 dvss.n462 dvss.n461 9.3005
R778 dvss.n463 dvss.n132 9.3005
R779 dvss.n465 dvss.n464 9.3005
R780 dvss.n466 dvss.n131 9.3005
R781 dvss.n468 dvss.n467 9.3005
R782 dvss.n469 dvss.n130 9.3005
R783 dvss.n471 dvss.n470 9.3005
R784 dvss.n472 dvss.n129 9.3005
R785 dvss.n474 dvss.n473 9.3005
R786 dvss.n475 dvss.n128 9.3005
R787 dvss.n477 dvss.n476 9.3005
R788 dvss.n478 dvss.n125 9.3005
R789 dvss.n479 dvss.n124 9.3005
R790 dvss.n481 dvss.n480 9.3005
R791 dvss.n483 dvss.n482 9.3005
R792 dvss.n484 dvss.n121 9.3005
R793 dvss.n487 dvss.n486 9.3005
R794 dvss.n488 dvss.n120 9.3005
R795 dvss.n490 dvss.n489 9.3005
R796 dvss.n491 dvss.n118 9.3005
R797 dvss.n494 dvss.n493 9.3005
R798 dvss.n495 dvss.n117 9.3005
R799 dvss.n497 dvss.n496 9.3005
R800 dvss.n498 dvss.n116 9.3005
R801 dvss.n502 dvss.n501 9.3005
R802 dvss.n503 dvss.n115 9.3005
R803 dvss.n505 dvss.n504 9.3005
R804 dvss.n506 dvss.n114 9.3005
R805 dvss.n508 dvss.n507 9.3005
R806 dvss.n509 dvss.n113 9.3005
R807 dvss.n511 dvss.n510 9.3005
R808 dvss.n512 dvss.n112 9.3005
R809 dvss.n514 dvss.n513 9.3005
R810 dvss.n515 dvss.n111 9.3005
R811 dvss.n517 dvss.n516 9.3005
R812 dvss.n519 dvss.n518 9.3005
R813 dvss.n250 dvss.n108 9.3005
R814 dvss.n252 dvss.n251 9.3005
R815 dvss.n254 dvss.n253 9.3005
R816 dvss.n255 dvss.n247 9.3005
R817 dvss.n258 dvss.n257 9.3005
R818 dvss.n259 dvss.n246 9.3005
R819 dvss.n261 dvss.n260 9.3005
R820 dvss.n262 dvss.n244 9.3005
R821 dvss.n265 dvss.n264 9.3005
R822 dvss.n266 dvss.n243 9.3005
R823 dvss.n268 dvss.n267 9.3005
R824 dvss.n269 dvss.n242 9.3005
R825 dvss.n273 dvss.n272 9.3005
R826 dvss.n274 dvss.n241 9.3005
R827 dvss.n276 dvss.n275 9.3005
R828 dvss.n277 dvss.n240 9.3005
R829 dvss.n279 dvss.n278 9.3005
R830 dvss.n280 dvss.n239 9.3005
R831 dvss.n282 dvss.n281 9.3005
R832 dvss.n283 dvss.n238 9.3005
R833 dvss.n285 dvss.n284 9.3005
R834 dvss.n286 dvss.n237 9.3005
R835 dvss.n288 dvss.n287 9.3005
R836 dvss.n290 dvss.n289 9.3005
R837 dvss.n291 dvss.n226 9.3005
R838 dvss.n293 dvss.n292 9.3005
R839 dvss.n297 dvss.n296 9.3005
R840 dvss.n298 dvss.n225 9.3005
R841 dvss.n300 dvss.n299 9.3005
R842 dvss.n301 dvss.n224 9.3005
R843 dvss.n662 dvss.n7 9.3005
R844 dvss.n667 dvss.n666 9.3005
R845 dvss.n673 dvss.n672 9.3005
R846 dvss.n671 dvss.n4 9.3005
R847 dvss.n670 dvss.n669 9.3005
R848 dvss.n668 dvss.n5 9.3005
R849 dvss.n665 dvss.n664 9.3005
R850 dvss.n674 dvss.n3 9.3005
R851 dvss.n676 dvss.n675 9.3005
R852 dvss.n640 dvss.n639 9.3005
R853 dvss.n24 dvss.n20 9.3005
R854 dvss.n26 dvss.n25 9.3005
R855 dvss.n644 dvss.n13 9.3005
R856 dvss.n77 dvss.n76 9.3005
R857 dvss.n73 dvss.n67 9.3005
R858 dvss.n635 dvss.n634 8.88939
R859 dvss.n68 dvss.n65 8.77764
R860 dvss.n528 dvss.n103 8.43597
R861 dvss.n271 dvss.n241 7.90638
R862 dvss.n500 dvss.n115 7.90638
R863 dvss.n460 dvss.n132 7.90638
R864 dvss.n412 dvss.n411 7.90638
R865 dvss.n373 dvss.n372 7.90638
R866 dvss.n334 dvss.n333 7.90638
R867 dvss.n620 dvss.n619 7.40556
R868 dvss.n621 dvss.n620 7.40556
R869 dvss.n603 dvss.n602 7.17831
R870 dvss.n75 dvss.n66 7.17078
R871 dvss.n26 dvss 7.15344
R872 dvss.n76 dvss 7.15344
R873 dvss.n569 dvss.n50 7.1196
R874 dvss.n257 dvss.n256 6.77697
R875 dvss.n486 dvss.n485 6.77697
R876 dvss.n446 dvss.n445 6.77697
R877 dvss.n427 dvss.n151 6.77697
R878 dvss.n387 dvss.n386 6.77697
R879 dvss.n348 dvss.n347 6.77697
R880 dvss.n538 dvss.n537 6.7205
R881 dvss.n216 dvss.n196 6.7005
R882 dvss.n679 dvss.n677 6.56103
R883 dvss.n525 dvss.n104 6.53261
R884 dvss.n230 dvss.n82 6.36591
R885 dvss.n602 dvss.n601 5.73579
R886 dvss.n621 dvss.n34 5.34031
R887 dvss.n598 dvss.n47 5.31835
R888 dvss.n565 dvss.n564 5.28896
R889 dvss.n572 dvss.n86 5.28896
R890 dvss.n609 dvss.n47 4.48642
R891 dvss.n555 dvss.t54 4.3505
R892 dvss.n555 dvss.t58 4.3505
R893 dvss.n556 dvss.t70 4.3505
R894 dvss.n556 dvss.t74 4.3505
R895 dvss.n548 dvss.t44 4.3505
R896 dvss.n548 dvss.t48 4.3505
R897 dvss.n547 dvss.t56 4.3505
R898 dvss.n547 dvss.t64 4.3505
R899 dvss.n529 dvss.n528 4.00961
R900 dvss.n577 dvss.n576 3.89404
R901 dvss.n583 dvss.n582 3.84425
R902 dvss.n602 dvss.n17 3.58941
R903 dvss.n579 dvss.n36 3.56414
R904 dvss.n584 dvss.n583 3.54405
R905 dvss.n251 dvss.n249 3.38874
R906 dvss.n480 dvss.n123 3.38874
R907 dvss.n440 dvss.n140 3.38874
R908 dvss.n150 dvss.n147 3.38874
R909 dvss.n393 dvss.n392 3.38874
R910 dvss.n354 dvss.n353 3.38874
R911 dvss.n666 dvss 3.29747
R912 dvss.n680 dvss.n1 3.21038
R913 dvss.n539 dvss.n96 3.01827
R914 dvss.n650 dvss.n649 2.88227
R915 dvss.n567 dvss.n566 2.75993
R916 dvss.n566 dvss.n565 2.75993
R917 dvss.n568 dvss.n87 2.75993
R918 dvss.n564 dvss.n87 2.75993
R919 dvss.n563 dvss.n91 2.64473
R920 dvss.n264 dvss.n263 2.63579
R921 dvss.n493 dvss.n492 2.63579
R922 dvss.n453 dvss.n452 2.63579
R923 dvss.n419 dvss.n154 2.63579
R924 dvss.n380 dvss.n172 2.63579
R925 dvss.n341 dvss.n189 2.63579
R926 dvss.n632 dvss.n22 2.47305
R927 dvss.n67 dvss.n65 2.41042
R928 dvss.n634 dvss.n22 2.33976
R929 dvss.n530 dvss.n96 2.3185
R930 dvss.n575 dvss.n82 1.98969
R931 dvss.n677 dvss.n1 1.93239
R932 dvss.n41 dvss.n36 1.92484
R933 dvss.n272 dvss.n271 1.88285
R934 dvss.n501 dvss.n500 1.88285
R935 dvss.n461 dvss.n460 1.88285
R936 dvss.n413 dvss.n412 1.88285
R937 dvss.n374 dvss.n373 1.88285
R938 dvss.n335 dvss.n334 1.88285
R939 dvss.n103 dvss.n102 1.85983
R940 dvss.n597 dvss.n46 1.80934
R941 dvss.n560 dvss.n559 1.57196
R942 dvss.n551 dvss.n550 1.57139
R943 dvss.n208 dvss.n194 1.5505
R944 dvss.n618 dvss.n18 1.48151
R945 dvss.n34 dvss.n18 1.48151
R946 dvss.n585 dvss.n584 1.46336
R947 dvss.n654 dvss.n14 1.32907
R948 dvss.n591 dvss.n590 1.32907
R949 dvss.n530 dvss.n529 1.21052
R950 dvss.n326 dvss.n196 1.11858
R951 dvss.n566 dvss.n87 1.10724
R952 dvss.n571 dvss.n88 1.10724
R953 dvss.n579 dvss.n37 1.01868
R954 dvss.n567 dvss.n89 0.899376
R955 dvss.n618 dvss.n19 0.804872
R956 dvss.n593 dvss.n38 0.778315
R957 dvss.n575 dvss.n574 0.774309
R958 dvss.n574 dvss.n573 0.774309
R959 dvss.n214 dvss.n208 0.649775
R960 dvss.n296 dvss.n295 0.630008
R961 dvss.n310 dvss.n205 0.630008
R962 dvss.n536 dvss.n89 0.629714
R963 dvss.n620 dvss.n18 0.538751
R964 dvss.n610 dvss.n46 0.533285
R965 dvss.n233 dvss.n232 0.519117
R966 dvss.n234 dvss.n233 0.519117
R967 dvss.n535 dvss.n533 0.482579
R968 dvss.t77 dvss.n657 0.474702
R969 dvss.n657 dvss.n656 0.447064
R970 dvss.n529 dvss.n100 0.443357
R971 dvss.n531 dvss.n530 0.443357
R972 dvss.n227 dvss.n104 0.428132
R973 dvss.n227 dvss.n146 0.428132
R974 dvss.n522 dvss.n104 0.411509
R975 dvss.n616 dvss.n38 0.362946
R976 dvss.n526 dvss.n90 0.355045
R977 dvss.n211 dvss.n90 0.355045
R978 dvss.n604 dvss.n601 0.336965
R979 dvss.n600 dvss.n17 0.328522
R980 dvss.n103 dvss 0.326572
R981 dvss.n605 dvss.n600 0.326101
R982 dvss.n592 dvss.n11 0.313726
R983 dvss.n557 dvss.n82 0.277008
R984 dvss.n662 dvss.n661 0.274194
R985 dvss.n534 dvss.n51 0.271039
R986 dvss.n583 dvss.n78 0.262597
R987 dvss.n611 dvss.n610 0.2605
R988 dvss.n612 dvss.n611 0.2605
R989 dvss.n539 dvss.n538 0.248336
R990 dvss.n81 dvss.n80 0.218682
R991 dvss.n608 dvss.n48 0.210906
R992 dvss.n642 dvss.n641 0.206439
R993 dvss.n595 dvss.n48 0.202526
R994 dvss.n187 dvss.t116 0.189075
R995 dvss.n525 dvss.n524 0.181217
R996 dvss.n633 dvss.n632 0.178278
R997 dvss.n582 dvss.n581 0.170143
R998 dvss.n607 dvss.n606 0.166164
R999 dvss.n601 dvss.n600 0.155797
R1000 dvss dvss.n660 0.150986
R1001 dvss.n51 dvss.n50 0.145813
R1002 dvss.n325 dvss 0.142307
R1003 dvss.n222 dvss 0.140841
R1004 dvss.n660 dvss.n659 0.13579
R1005 dvss.n607 dvss.n599 0.130165
R1006 dvss.n223 dvss 0.127978
R1007 dvss.n223 dvss.n222 0.123227
R1008 dvss.n532 dvss.n531 0.122311
R1009 dvss.n523 dvss.n106 0.121873
R1010 dvss.n324 dvss.n323 0.120292
R1011 dvss.n323 dvss.n197 0.120292
R1012 dvss.n319 dvss.n197 0.120292
R1013 dvss.n319 dvss.n318 0.120292
R1014 dvss.n318 dvss.n317 0.120292
R1015 dvss.n313 dvss.n312 0.120292
R1016 dvss.n311 dvss.n203 0.120292
R1017 dvss.n307 dvss.n203 0.120292
R1018 dvss.n668 dvss.n667 0.120292
R1019 dvss.n669 dvss.n668 0.120292
R1020 dvss.n669 dvss.n4 0.120292
R1021 dvss.n673 dvss.n4 0.120292
R1022 dvss.n674 dvss.n673 0.120292
R1023 dvss.n675 dvss.n674 0.120292
R1024 dvss.n144 dvss.n143 0.104964
R1025 dvss.n312 dvss 0.104667
R1026 dvss.n594 dvss.n51 0.103194
R1027 dvss.n326 dvss 0.0999624
R1028 dvss.n667 dvss 0.0968542
R1029 dvss.n643 dvss 0.0941255
R1030 dvss.n606 dvss.n605 0.0879466
R1031 dvss.n648 dvss.n647 0.0850455
R1032 dvss.n66 dvss 0.080434
R1033 dvss.n221 dvss 0.0781256
R1034 dvss.n77 dvss.n66 0.0777204
R1035 dvss.n645 dvss 0.0770968
R1036 dvss.n578 dvss.n577 0.0749
R1037 dvss.n524 dvss.n523 0.0737044
R1038 dvss.n568 dvss.n567 0.0724101
R1039 dvss.n570 dvss.n569 0.0724101
R1040 dvss.t115 dvss.t114 0.070611
R1041 dvss.n560 dvss.n554 0.0678684
R1042 dvss.n658 dvss.t77 0.0675999
R1043 dvss.n552 dvss.n551 0.0671667
R1044 dvss.n595 dvss.n594 0.06684
R1045 dvss.n222 dvss.n221 0.0638562
R1046 dvss.n557 dvss 0.0633141
R1047 dvss.n581 dvss.n580 0.0614929
R1048 dvss.n659 dvss.t116 0.060491
R1049 dvss.n201 dvss 0.0603958
R1050 dvss.n313 dvss 0.0603958
R1051 dvss dvss.n306 0.0603958
R1052 dvss.n664 dvss 0.0603958
R1053 dvss.n657 dvss.n11 0.0595861
R1054 dvss.n221 dvss.n8 0.0586797
R1055 dvss.n98 dvss.n9 0.0559625
R1056 dvss.n143 dvss.n49 0.0535781
R1057 dvss.n608 dvss.n607 0.0533794
R1058 dvss.n1 dvss 0.0525833
R1059 dvss.n14 dvss 0.0515042
R1060 dvss.n25 dvss.n20 0.0480207
R1061 dvss.n643 dvss.n642 0.0476863
R1062 dvss.n524 dvss.n105 0.0461989
R1063 dvss.n550 dvss.n549 0.0457733
R1064 dvss.n325 dvss.n324 0.0447708
R1065 dvss.n658 dvss.n10 0.0405094
R1066 dvss.n642 dvss.n21 0.0402727
R1067 dvss.n593 dvss.n592 0.0393298
R1068 dvss.n531 dvss.n100 0.0374705
R1069 dvss.n619 dvss.n618 0.0354727
R1070 dvss dvss.n591 0.0347199
R1071 dvss.n559 dvss 0.0346686
R1072 dvss.n580 dvss.n579 0.0341957
R1073 dvss dvss.n201 0.0330521
R1074 dvss.n306 dvss 0.0330521
R1075 dvss.n19 dvss.n11 0.0323493
R1076 dvss.n656 dvss 0.0323446
R1077 dvss.n534 dvss.n89 0.0321327
R1078 dvss.n48 dvss.n46 0.0315
R1079 dvss.n581 dvss.n578 0.0306418
R1080 dvss.n532 dvss.n99 0.0284126
R1081 dvss dvss.n662 0.0271393
R1082 dvss.n592 dvss 0.0255
R1083 dvss.n641 dvss.n22 0.0247851
R1084 dvss.n641 dvss.n640 0.0242603
R1085 dvss.n25 dvss 0.0242603
R1086 dvss.n21 dvss 0.0242603
R1087 dvss.n536 dvss.n535 0.0239848
R1088 dvss.n664 dvss 0.0239375
R1089 dvss.n647 dvss.n645 0.0230951
R1090 dvss.n549 dvss.n10 0.0228519
R1091 dvss.n317 dvss 0.0226354
R1092 dvss.n307 dvss 0.0226354
R1093 dvss.n78 dvss 0.0215598
R1094 dvss.n8 dvss 0.0206613
R1095 dvss.n231 dvss.n9 0.0206307
R1096 dvss.n663 dvss 0.0199672
R1097 dvss.n523 dvss.n522 0.0192879
R1098 dvss.n521 dvss.n520 0.0189524
R1099 dvss.n596 dvss.n595 0.0189524
R1100 dvss.n558 dvss.n557 0.0184385
R1101 dvss.n67 dvss 0.0174837
R1102 dvss.n578 dvss.n79 0.0174213
R1103 dvss.n609 dvss.n608 0.0166458
R1104 dvss dvss.n311 0.016125
R1105 dvss.n432 dvss.n431 0.015957
R1106 dvss.n431 dvss.n430 0.015957
R1107 dvss.n430 dvss.n148 0.015957
R1108 dvss.n426 dvss.n148 0.015957
R1109 dvss.n426 dvss.n425 0.015957
R1110 dvss.n425 dvss.n152 0.015957
R1111 dvss.n421 dvss.n152 0.015957
R1112 dvss.n421 dvss.n420 0.015957
R1113 dvss.n420 dvss.n155 0.015957
R1114 dvss.n416 dvss.n155 0.015957
R1115 dvss.n416 dvss.n415 0.015957
R1116 dvss.n415 dvss.n414 0.015957
R1117 dvss.n414 dvss.n157 0.015957
R1118 dvss.n409 dvss.n157 0.015957
R1119 dvss.n409 dvss.n408 0.015957
R1120 dvss.n408 dvss.n407 0.015957
R1121 dvss.n407 dvss.n160 0.015957
R1122 dvss.n403 dvss.n160 0.015957
R1123 dvss.n403 dvss.n402 0.015957
R1124 dvss.n402 dvss.n401 0.015957
R1125 dvss.n401 dvss.n162 0.015957
R1126 dvss.n397 dvss.n162 0.015957
R1127 dvss.n395 dvss.n165 0.015957
R1128 dvss.n390 dvss.n165 0.015957
R1129 dvss.n390 dvss.n389 0.015957
R1130 dvss.n389 dvss.n388 0.015957
R1131 dvss.n388 dvss.n168 0.015957
R1132 dvss.n383 dvss.n168 0.015957
R1133 dvss.n383 dvss.n382 0.015957
R1134 dvss.n382 dvss.n381 0.015957
R1135 dvss.n381 dvss.n170 0.015957
R1136 dvss.n377 dvss.n170 0.015957
R1137 dvss.n377 dvss.n376 0.015957
R1138 dvss.n376 dvss.n375 0.015957
R1139 dvss.n375 dvss.n174 0.015957
R1140 dvss.n370 dvss.n174 0.015957
R1141 dvss.n370 dvss.n369 0.015957
R1142 dvss.n369 dvss.n368 0.015957
R1143 dvss.n368 dvss.n177 0.015957
R1144 dvss.n364 dvss.n177 0.015957
R1145 dvss.n364 dvss.n363 0.015957
R1146 dvss.n363 dvss.n362 0.015957
R1147 dvss.n362 dvss.n179 0.015957
R1148 dvss.n358 dvss.n179 0.015957
R1149 dvss.n356 dvss.n182 0.015957
R1150 dvss.n351 dvss.n182 0.015957
R1151 dvss.n351 dvss.n350 0.015957
R1152 dvss.n350 dvss.n349 0.015957
R1153 dvss.n349 dvss.n185 0.015957
R1154 dvss.n344 dvss.n185 0.015957
R1155 dvss.n344 dvss.n343 0.015957
R1156 dvss.n343 dvss.n342 0.015957
R1157 dvss.n339 dvss.n338 0.015957
R1158 dvss.n338 dvss.n337 0.015957
R1159 dvss.n337 dvss.n191 0.015957
R1160 dvss.n332 dvss.n191 0.015957
R1161 dvss.n332 dvss.n331 0.015957
R1162 dvss.n331 dvss.n330 0.015957
R1163 dvss.n326 dvss.n325 0.0141555
R1164 dvss.n644 dvss.n643 0.0140978
R1165 dvss.n640 dvss 0.0139298
R1166 dvss.n441 dvss.n141 0.0125293
R1167 dvss.n442 dvss.n441 0.0125293
R1168 dvss.n442 dvss.n138 0.0125293
R1169 dvss.n447 dvss.n138 0.0125293
R1170 dvss.n448 dvss.n447 0.0125293
R1171 dvss.n449 dvss.n448 0.0125293
R1172 dvss.n449 dvss.n135 0.0125293
R1173 dvss.n454 dvss.n135 0.0125293
R1174 dvss.n455 dvss.n454 0.0125293
R1175 dvss.n456 dvss.n455 0.0125293
R1176 dvss.n456 dvss.n133 0.0125293
R1177 dvss.n462 dvss.n133 0.0125293
R1178 dvss.n463 dvss.n462 0.0125293
R1179 dvss.n464 dvss.n463 0.0125293
R1180 dvss.n464 dvss.n131 0.0125293
R1181 dvss.n468 dvss.n131 0.0125293
R1182 dvss.n469 dvss.n468 0.0125293
R1183 dvss.n470 dvss.n469 0.0125293
R1184 dvss.n470 dvss.n129 0.0125293
R1185 dvss.n474 dvss.n129 0.0125293
R1186 dvss.n475 dvss.n474 0.0125293
R1187 dvss.n476 dvss.n475 0.0125293
R1188 dvss.n481 dvss.n124 0.0125293
R1189 dvss.n482 dvss.n481 0.0125293
R1190 dvss.n482 dvss.n121 0.0125293
R1191 dvss.n487 dvss.n121 0.0125293
R1192 dvss.n488 dvss.n487 0.0125293
R1193 dvss.n489 dvss.n488 0.0125293
R1194 dvss.n489 dvss.n118 0.0125293
R1195 dvss.n494 dvss.n118 0.0125293
R1196 dvss.n495 dvss.n494 0.0125293
R1197 dvss.n496 dvss.n495 0.0125293
R1198 dvss.n496 dvss.n116 0.0125293
R1199 dvss.n502 dvss.n116 0.0125293
R1200 dvss.n503 dvss.n502 0.0125293
R1201 dvss.n504 dvss.n503 0.0125293
R1202 dvss.n504 dvss.n114 0.0125293
R1203 dvss.n508 dvss.n114 0.0125293
R1204 dvss.n509 dvss.n508 0.0125293
R1205 dvss.n510 dvss.n509 0.0125293
R1206 dvss.n510 dvss.n112 0.0125293
R1207 dvss.n514 dvss.n112 0.0125293
R1208 dvss.n515 dvss.n514 0.0125293
R1209 dvss.n516 dvss.n515 0.0125293
R1210 dvss.n252 dvss.n250 0.0125293
R1211 dvss.n253 dvss.n252 0.0125293
R1212 dvss.n253 dvss.n247 0.0125293
R1213 dvss.n258 dvss.n247 0.0125293
R1214 dvss.n259 dvss.n258 0.0125293
R1215 dvss.n260 dvss.n259 0.0125293
R1216 dvss.n260 dvss.n244 0.0125293
R1217 dvss.n265 dvss.n244 0.0125293
R1218 dvss.n266 dvss.n265 0.0125293
R1219 dvss.n267 dvss.n266 0.0125293
R1220 dvss.n267 dvss.n242 0.0125293
R1221 dvss.n273 dvss.n242 0.0125293
R1222 dvss.n274 dvss.n273 0.0125293
R1223 dvss.n275 dvss.n274 0.0125293
R1224 dvss.n275 dvss.n240 0.0125293
R1225 dvss.n279 dvss.n240 0.0125293
R1226 dvss.n280 dvss.n279 0.0125293
R1227 dvss.n281 dvss.n280 0.0125293
R1228 dvss.n281 dvss.n238 0.0125293
R1229 dvss.n285 dvss.n238 0.0125293
R1230 dvss.n286 dvss.n285 0.0125293
R1231 dvss.n287 dvss.n286 0.0125293
R1232 dvss.n292 dvss.n291 0.0125293
R1233 dvss.n298 dvss.n297 0.0125293
R1234 dvss.n299 dvss.n298 0.0125293
R1235 dvss.n339 dvss.n187 0.0122608
R1236 dvss dvss.n558 0.0110353
R1237 dvss.n292 dvss 0.0109603
R1238 dvss.n78 dvss.n77 0.0106902
R1239 dvss.n659 dvss.t115 0.0106199
R1240 dvss.n580 dvss.n53 0.0101631
R1241 dvss.n327 dvss.n194 0.0099086
R1242 dvss.n661 dvss.n8 0.00990439
R1243 dvss.n660 dvss.n9 0.00933152
R1244 dvss.n675 dvss.n1 0.0083125
R1245 dvss.n642 dvss.n20 0.00824793
R1246 dvss.n535 dvss.n534 0.00822968
R1247 dvss.n432 dvss 0.00822849
R1248 dvss dvss.n396 0.00822849
R1249 dvss dvss.n395 0.00822849
R1250 dvss dvss.n357 0.00822849
R1251 dvss dvss.n356 0.00822849
R1252 dvss.n647 dvss.n646 0.00789958
R1253 dvss.n330 dvss.n194 0.00654839
R1254 dvss.n141 dvss 0.00651464
R1255 dvss dvss.n125 0.00651464
R1256 dvss dvss.n124 0.00651464
R1257 dvss.n250 dvss 0.00651464
R1258 dvss.n290 dvss 0.00651464
R1259 dvss.n291 dvss 0.00651464
R1260 dvss dvss.n224 0.00651464
R1261 dvss.n520 dvss.n519 0.00573013
R1262 dvss dvss.n1 0.00570833
R1263 dvss.n557 dvss.n10 0.00519818
R1264 dvss.n661 dvss 0.00481034
R1265 dvss dvss.n105 0.00470027
R1266 dvss.n396 dvss 0.00470027
R1267 dvss.n357 dvss 0.00470027
R1268 dvss.n342 dvss.n187 0.00419624
R1269 dvss.n645 dvss.n644 0.00411776
R1270 dvss dvss.n106 0.00376883
R1271 dvss.n125 dvss 0.00376883
R1272 dvss.n519 dvss 0.00376883
R1273 dvss dvss.n290 0.00376883
R1274 dvss.n224 dvss 0.00376883
R1275 dvss.t114 dvss.n658 0.00351108
R1276 dvss.n397 dvss 0.00335618
R1277 dvss.n358 dvss 0.00335618
R1278 dvss.n476 dvss 0.0027228
R1279 dvss.n516 dvss 0.0027228
R1280 dvss.n287 dvss 0.0027228
R1281 dvss.n299 dvss 0.0027228
R1282 dvss.n297 dvss 0.00206904
R1283 dvss dvss.n663 0.00180208
R1284 dvss.n533 dvss.n532 0.00156293
R1285 dvss.n663 dvss 0.00152459
R1286 dvss.n327 dvss.n326 0.00150806
R1287 dvss.n520 dvss 0.00128452
R1288 dvss dvss.n223 0.00077533
R1289 dvss.n646 dvss.n14 0.000632135
R1290 dvss.n591 dvss.n53 0.000588652
R1291 dvdd.n295 dvdd.n286 5128.23
R1292 dvdd.n295 dvdd.n287 5128.23
R1293 dvdd.n293 dvdd.n287 5128.23
R1294 dvdd.n293 dvdd.n286 5128.23
R1295 dvdd.n42 dvdd.n5 1736.47
R1296 dvdd.n45 dvdd.n4 1736.47
R1297 dvdd.n30 dvdd.n27 1736.47
R1298 dvdd.n33 dvdd.n29 1736.47
R1299 dvdd.n255 dvdd.t45 838.817
R1300 dvdd.n69 dvdd.t105 806.511
R1301 dvdd.n69 dvdd.t82 806.511
R1302 dvdd.n90 dvdd.t100 806.511
R1303 dvdd.n90 dvdd.t165 806.511
R1304 dvdd.n111 dvdd.t7 806.511
R1305 dvdd.n111 dvdd.t75 806.511
R1306 dvdd.n292 dvdd.n284 787.447
R1307 dvdd.n292 dvdd.n285 786.827
R1308 dvdd.n56 dvdd.t65 668.683
R1309 dvdd.n56 dvdd.t64 668.683
R1310 dvdd.n227 dvdd.t88 667.778
R1311 dvdd.n227 dvdd.t98 667.778
R1312 dvdd.n189 dvdd.t59 667.778
R1313 dvdd.n189 dvdd.t102 667.778
R1314 dvdd.n151 dvdd.t20 667.778
R1315 dvdd.n151 dvdd.t109 667.778
R1316 dvdd.n296 dvdd.n284 604.574
R1317 dvdd.n73 dvdd.n71 604.457
R1318 dvdd.n73 dvdd.n72 604.457
R1319 dvdd.n94 dvdd.n92 604.457
R1320 dvdd.n94 dvdd.n93 604.457
R1321 dvdd.n115 dvdd.n113 604.457
R1322 dvdd.n115 dvdd.n114 604.457
R1323 dvdd.n232 dvdd.n61 604.394
R1324 dvdd.n232 dvdd.n62 604.394
R1325 dvdd.n194 dvdd.n82 604.394
R1326 dvdd.n194 dvdd.n83 604.394
R1327 dvdd.n156 dvdd.n103 604.394
R1328 dvdd.n156 dvdd.n104 604.394
R1329 dvdd.n220 dvdd.n67 601.679
R1330 dvdd.n220 dvdd.n68 601.679
R1331 dvdd.n182 dvdd.n88 601.679
R1332 dvdd.n182 dvdd.n89 601.679
R1333 dvdd.n144 dvdd.n109 601.679
R1334 dvdd.n144 dvdd.n110 601.679
R1335 dvdd.n260 dvdd.n259 585
R1336 dvdd.t66 dvdd.t44 556.386
R1337 dvdd.n246 dvdd 538.664
R1338 dvdd.n18 dvdd 535.705
R1339 dvdd.n11 dvdd 535.705
R1340 dvdd.t37 dvdd 473.521
R1341 dvdd.t19 dvdd.t84 448.146
R1342 dvdd.t58 dvdd.t128 448.146
R1343 dvdd.t87 dvdd.t35 448.146
R1344 dvdd.n296 dvdd.n285 423.062
R1345 dvdd.t93 dvdd.t95 367.579
R1346 dvdd.t29 dvdd.t27 367.579
R1347 dvdd.t14 dvdd.t12 367.579
R1348 dvdd.n274 dvdd.t23 360.005
R1349 dvdd.t6 dvdd.t52 330.654
R1350 dvdd.t99 dvdd.t42 330.654
R1351 dvdd.t81 dvdd.t48 330.654
R1352 dvdd.n43 dvdd.n4 314.781
R1353 dvdd.n44 dvdd.n5 314.781
R1354 dvdd.n31 dvdd.n29 314.781
R1355 dvdd.n32 dvdd.n27 314.781
R1356 dvdd.n23 dvdd.n17 312.053
R1357 dvdd.n9 dvdd.n8 312.051
R1358 dvdd.n266 dvdd.n256 312.051
R1359 dvdd.t168 dvdd.t170 304.829
R1360 dvdd.t44 dvdd.t106 284.113
R1361 dvdd.t95 dvdd.t121 275.265
R1362 dvdd.t27 dvdd.t114 275.265
R1363 dvdd.t12 dvdd.t110 275.265
R1364 dvdd.t106 dvdd.t37 275.235
R1365 dvdd.n271 dvdd.t0 261.837
R1366 dvdd.t131 dvdd.t119 260.437
R1367 dvdd.t39 dvdd.t166 260.437
R1368 dvdd.n207 dvdd.n76 259.707
R1369 dvdd.n207 dvdd.n75 259.707
R1370 dvdd.n169 dvdd.n97 259.707
R1371 dvdd.n169 dvdd.n96 259.707
R1372 dvdd.n131 dvdd.n118 259.707
R1373 dvdd.n131 dvdd.n117 259.707
R1374 dvdd.t0 dvdd.t17 258.481
R1375 dvdd.n273 dvdd.t56 253.446
R1376 dvdd.n272 dvdd.t103 253.446
R1377 dvdd.t163 dvdd.t21 248.599
R1378 dvdd.t21 dvdd.t66 248.599
R1379 dvdd.n201 dvdd.n80 242.607
R1380 dvdd.n163 dvdd.n101 242.607
R1381 dvdd.n125 dvdd.n123 242.607
R1382 dvdd.n201 dvdd.n79 242.607
R1383 dvdd.n163 dvdd.n100 242.607
R1384 dvdd.n125 dvdd.n122 242.607
R1385 dvdd.t2 dvdd.t83 234.982
R1386 dvdd.t31 dvdd.t127 234.982
R1387 dvdd.t76 dvdd.t33 234.982
R1388 dvdd dvdd.n270 232.445
R1389 dvdd.n0 dvdd.t146 228.215
R1390 dvdd.n0 dvdd.t74 228.215
R1391 dvdd.n239 dvdd.n59 215.123
R1392 dvdd.n239 dvdd.n238 215.123
R1393 dvdd.t170 dvdd.t62 213.084
R1394 dvdd.n41 dvdd.n3 185.225
R1395 dvdd.n46 dvdd.n3 185.225
R1396 dvdd.n34 dvdd.n28 185.225
R1397 dvdd.n28 dvdd.n26 185.225
R1398 dvdd.t54 dvdd.t91 181.273
R1399 dvdd.t46 dvdd.t25 181.273
R1400 dvdd.t50 dvdd.t10 181.273
R1401 dvdd.t86 dvdd.t6 166.167
R1402 dvdd.t83 dvdd.t137 166.167
R1403 dvdd.t130 dvdd.t99 166.167
R1404 dvdd.t127 dvdd.t117 166.167
R1405 dvdd.t34 dvdd.t81 166.167
R1406 dvdd.t33 dvdd.t5 166.167
R1407 dvdd.t23 dvdd.t93 162.81
R1408 dvdd.t52 dvdd.t2 162.81
R1409 dvdd.t56 dvdd.t29 162.81
R1410 dvdd.t42 dvdd.t31 162.81
R1411 dvdd.t103 dvdd.t14 162.81
R1412 dvdd.t48 dvdd.t76 162.81
R1413 dvdd.t147 dvdd.n293 161.316
R1414 dvdd.n295 dvdd.t161 161.316
R1415 dvdd.t137 dvdd.t19 154.417
R1416 dvdd.t117 dvdd.t58 154.417
R1417 dvdd.t5 dvdd.t87 154.417
R1418 dvdd.t17 dvdd.t63 147.703
R1419 dvdd.n75 dvdd.t135 147.111
R1420 dvdd.n76 dvdd.t111 147.111
R1421 dvdd.n96 dvdd.t115 147.111
R1422 dvdd.n97 dvdd.t136 147.111
R1423 dvdd.n117 dvdd.t164 147.111
R1424 dvdd.n118 dvdd.t122 147.111
R1425 dvdd.t138 dvdd.t86 144.346
R1426 dvdd.t116 dvdd.t130 144.346
R1427 dvdd.t4 dvdd.t34 144.346
R1428 dvdd.t121 dvdd.t54 140.989
R1429 dvdd.t91 dvdd.t138 140.989
R1430 dvdd.t84 dvdd.t60 140.989
R1431 dvdd.t114 dvdd.t46 140.989
R1432 dvdd.t25 dvdd.t116 140.989
R1433 dvdd.t128 dvdd.t89 140.989
R1434 dvdd.t110 dvdd.t50 140.989
R1435 dvdd.t10 dvdd.t4 140.989
R1436 dvdd.t35 dvdd.t8 140.989
R1437 dvdd.t63 dvdd 132.597
R1438 dvdd dvdd.n273 125.883
R1439 dvdd dvdd.n272 125.883
R1440 dvdd dvdd.n271 125.883
R1441 dvdd.t153 dvdd.t147 121.245
R1442 dvdd.t155 dvdd.t153 121.245
R1443 dvdd.t149 dvdd.t155 121.245
R1444 dvdd.t151 dvdd.t149 121.245
R1445 dvdd.t141 dvdd.t159 121.245
R1446 dvdd.t143 dvdd.t141 121.245
R1447 dvdd.t157 dvdd.t143 121.245
R1448 dvdd.t161 dvdd.t157 121.245
R1449 dvdd.n71 dvdd.t11 119.608
R1450 dvdd.n72 dvdd.t174 119.608
R1451 dvdd.n92 dvdd.t26 119.608
R1452 dvdd.n93 dvdd.t79 119.608
R1453 dvdd.n113 dvdd.t124 119.608
R1454 dvdd.n114 dvdd.t92 119.608
R1455 dvdd.t60 dvdd 109.1
R1456 dvdd.t89 dvdd 109.1
R1457 dvdd.t8 dvdd 109.1
R1458 dvdd.n75 dvdd.t13 108.413
R1459 dvdd.n76 dvdd.t173 108.413
R1460 dvdd.n96 dvdd.t28 108.413
R1461 dvdd.n97 dvdd.t78 108.413
R1462 dvdd.n117 dvdd.t123 108.413
R1463 dvdd.n118 dvdd.t96 108.413
R1464 dvdd.n271 dvdd.n55 106.559
R1465 dvdd.n272 dvdd.n54 106.559
R1466 dvdd.n273 dvdd.n53 106.559
R1467 dvdd.n47 dvdd.n2 105.412
R1468 dvdd.n40 dvdd.n2 105.412
R1469 dvdd.n37 dvdd.n36 105.412
R1470 dvdd.n36 dvdd.n35 105.412
R1471 dvdd dvdd.t168 100.624
R1472 dvdd.n67 dvdd.t77 93.81
R1473 dvdd.n68 dvdd.t112 93.81
R1474 dvdd.n88 dvdd.t32 93.81
R1475 dvdd.n89 dvdd.t139 93.81
R1476 dvdd.n109 dvdd.t118 93.81
R1477 dvdd.n110 dvdd.t3 93.81
R1478 dvdd dvdd.t131 91.745
R1479 dvdd dvdd.t39 91.745
R1480 dvdd dvdd.t163 88.7855
R1481 dvdd.n259 dvdd.t169 86.7743
R1482 dvdd.n47 dvdd.n46 79.8123
R1483 dvdd.n41 dvdd.n40 79.8123
R1484 dvdd.n35 dvdd.n34 79.8123
R1485 dvdd.n37 dvdd.n26 79.8123
R1486 dvdd.n59 dvdd.t18 74.7554
R1487 dvdd.n238 dvdd.t108 74.7554
R1488 dvdd.n67 dvdd.t70 63.3219
R1489 dvdd.n68 dvdd.t49 63.3219
R1490 dvdd.n71 dvdd.t71 63.3219
R1491 dvdd.n72 dvdd.t51 63.3219
R1492 dvdd.n88 dvdd.t68 63.3219
R1493 dvdd.n89 dvdd.t43 63.3219
R1494 dvdd.n92 dvdd.t69 63.3219
R1495 dvdd.n93 dvdd.t47 63.3219
R1496 dvdd.n109 dvdd.t72 63.3219
R1497 dvdd.n110 dvdd.t53 63.3219
R1498 dvdd.n113 dvdd.t67 63.3219
R1499 dvdd.n114 dvdd.t55 63.3219
R1500 dvdd.n79 dvdd.t15 61.9829
R1501 dvdd.n100 dvdd.t30 61.9829
R1502 dvdd.n122 dvdd.t125 61.9829
R1503 dvdd.n80 dvdd.t172 61.9826
R1504 dvdd.n101 dvdd.t80 61.9826
R1505 dvdd.n123 dvdd.t94 61.9826
R1506 dvdd.n259 dvdd.t171 61.05
R1507 dvdd.n294 dvdd.t151 60.6225
R1508 dvdd.t159 dvdd.n294 60.6225
R1509 dvdd.n292 dvdd.t148 60.3236
R1510 dvdd.n296 dvdd.t162 60.3236
R1511 dvdd.n297 dvdd.n283 54.7085
R1512 dvdd.n298 dvdd.n282 54.7085
R1513 dvdd.n290 dvdd.n289 54.7085
R1514 dvdd.n291 dvdd.n288 54.7085
R1515 dvdd.n61 dvdd.t41 41.5552
R1516 dvdd.n61 dvdd.t16 41.5552
R1517 dvdd.n62 dvdd.t36 41.5552
R1518 dvdd.n62 dvdd.t9 41.5552
R1519 dvdd.n82 dvdd.t129 41.5552
R1520 dvdd.n82 dvdd.t90 41.5552
R1521 dvdd.n83 dvdd.t140 41.5552
R1522 dvdd.n83 dvdd.t97 41.5552
R1523 dvdd.n103 dvdd.t85 41.5552
R1524 dvdd.n103 dvdd.t61 41.5552
R1525 dvdd.n104 dvdd.t126 41.5552
R1526 dvdd.n104 dvdd.t101 41.5552
R1527 dvdd.n46 dvdd.n45 37.0005
R1528 dvdd.n42 dvdd.n41 37.0005
R1529 dvdd.n34 dvdd.n33 37.0005
R1530 dvdd.n30 dvdd.n26 37.0005
R1531 dvdd.n17 dvdd.t132 36.1587
R1532 dvdd.n17 dvdd.t120 36.1587
R1533 dvdd.n8 dvdd.t40 36.1587
R1534 dvdd.n8 dvdd.t167 36.1587
R1535 dvdd.n256 dvdd.t107 35.4605
R1536 dvdd.n250 dvdd.n249 34.6358
R1537 dvdd.n254 dvdd.n245 34.6358
R1538 dvdd.n265 dvdd.n257 34.6358
R1539 dvdd.n231 dvdd.n63 34.6358
R1540 dvdd.n221 dvdd.n65 34.6358
R1541 dvdd.n225 dvdd.n65 34.6358
R1542 dvdd.n226 dvdd.n225 34.6358
R1543 dvdd.n219 dvdd.n218 34.6358
R1544 dvdd.n213 dvdd.n212 34.6358
R1545 dvdd.n214 dvdd.n213 34.6358
R1546 dvdd.n200 dvdd.n199 34.6358
R1547 dvdd.n202 dvdd.n77 34.6358
R1548 dvdd.n206 dvdd.n77 34.6358
R1549 dvdd.n193 dvdd.n84 34.6358
R1550 dvdd.n183 dvdd.n86 34.6358
R1551 dvdd.n187 dvdd.n86 34.6358
R1552 dvdd.n188 dvdd.n187 34.6358
R1553 dvdd.n181 dvdd.n180 34.6358
R1554 dvdd.n175 dvdd.n174 34.6358
R1555 dvdd.n176 dvdd.n175 34.6358
R1556 dvdd.n162 dvdd.n161 34.6358
R1557 dvdd.n164 dvdd.n98 34.6358
R1558 dvdd.n168 dvdd.n98 34.6358
R1559 dvdd.n155 dvdd.n105 34.6358
R1560 dvdd.n145 dvdd.n107 34.6358
R1561 dvdd.n149 dvdd.n107 34.6358
R1562 dvdd.n150 dvdd.n149 34.6358
R1563 dvdd.n143 dvdd.n142 34.6358
R1564 dvdd.n137 dvdd.n136 34.6358
R1565 dvdd.n138 dvdd.n137 34.6358
R1566 dvdd.n124 dvdd.n52 34.6358
R1567 dvdd.n126 dvdd.n119 34.6358
R1568 dvdd.n130 dvdd.n119 34.6358
R1569 dvdd.n239 dvdd.n58 33.8829
R1570 dvdd.n227 dvdd.n226 32.377
R1571 dvdd.n189 dvdd.n188 32.377
R1572 dvdd.n151 dvdd.n150 32.377
R1573 dvdd.n214 dvdd.n69 32.0005
R1574 dvdd.n176 dvdd.n90 32.0005
R1575 dvdd.n138 dvdd.n111 32.0005
R1576 dvdd.n240 dvdd.n239 31.624
R1577 dvdd.n202 dvdd.n201 31.2476
R1578 dvdd.n164 dvdd.n163 31.2476
R1579 dvdd.n126 dvdd.n125 31.2476
R1580 dvdd.n5 dvdd.n3 30.8338
R1581 dvdd.n4 dvdd.n2 30.8338
R1582 dvdd.n36 dvdd.n27 30.8338
R1583 dvdd.n29 dvdd.n28 30.8338
R1584 dvdd.n79 dvdd.t104 30.1745
R1585 dvdd.n100 dvdd.t57 30.1745
R1586 dvdd.n122 dvdd.t133 30.1745
R1587 dvdd.n80 dvdd.t134 30.1738
R1588 dvdd.n101 dvdd.t113 30.1738
R1589 dvdd.n123 dvdd.t24 30.1738
R1590 dvdd.n208 dvdd.n73 30.1181
R1591 dvdd.n170 dvdd.n94 30.1181
R1592 dvdd.n132 dvdd.n115 30.1181
R1593 dvdd.n43 dvdd.n42 29.6618
R1594 dvdd.n45 dvdd.n44 29.6618
R1595 dvdd.n31 dvdd.n30 29.6618
R1596 dvdd.n33 dvdd.n32 29.6618
R1597 dvdd.n59 dvdd.t1 28.5349
R1598 dvdd.n238 dvdd.t22 28.5349
R1599 dvdd.n261 dvdd.n257 28.2952
R1600 dvdd dvdd.n245 27.8593
R1601 dvdd.n256 dvdd.t38 26.5955
R1602 dvdd.n260 dvdd.n258 25.2079
R1603 dvdd.n22 dvdd.n18 23.7181
R1604 dvdd.n11 dvdd.n10 23.7181
R1605 dvdd.n249 dvdd.n246 23.7181
R1606 dvdd.n233 dvdd.n55 23.7181
R1607 dvdd.n199 dvdd.n54 23.7181
R1608 dvdd.n195 dvdd.n54 23.7181
R1609 dvdd.n161 dvdd.n53 23.7181
R1610 dvdd.n157 dvdd.n53 23.7181
R1611 dvdd.n274 dvdd.n52 23.7181
R1612 dvdd.n58 dvdd.n55 23.7181
R1613 dvdd.n232 dvdd.n231 22.9652
R1614 dvdd.n194 dvdd.n193 22.9652
R1615 dvdd.n156 dvdd.n155 22.9652
R1616 dvdd.n267 dvdd.n255 22.5887
R1617 dvdd.n266 dvdd.n265 22.5887
R1618 dvdd.n267 dvdd.n266 21.8358
R1619 dvdd.n233 dvdd.n232 21.4593
R1620 dvdd.n195 dvdd.n194 21.4593
R1621 dvdd.n157 dvdd.n156 21.4593
R1622 dvdd.n212 dvdd.n73 20.3299
R1623 dvdd.n174 dvdd.n94 20.3299
R1624 dvdd.n136 dvdd.n115 20.3299
R1625 dvdd.n255 dvdd.n254 19.9534
R1626 dvdd.n240 dvdd.n56 19.577
R1627 dvdd.n270 dvdd.n56 18.4476
R1628 dvdd.n227 dvdd.n63 18.0711
R1629 dvdd.n189 dvdd.n84 18.0711
R1630 dvdd.n151 dvdd.n105 18.0711
R1631 dvdd.n23 dvdd 15.8123
R1632 dvdd dvdd.n9 15.8123
R1633 dvdd.n296 dvdd.n295 13.2148
R1634 dvdd.n293 dvdd.n292 13.2148
R1635 dvdd.n38 dvdd.n37 10.0436
R1636 dvdd.n35 dvdd.n1 9.59217
R1637 dvdd.n218 dvdd.n69 9.41227
R1638 dvdd.n180 dvdd.n90 9.41227
R1639 dvdd.n142 dvdd.n111 9.41227
R1640 dvdd.n19 dvdd.n18 9.3005
R1641 dvdd.n22 dvdd.n21 9.3005
R1642 dvdd.n10 dvdd.n6 9.3005
R1643 dvdd.n12 dvdd.n11 9.3005
R1644 dvdd.n40 dvdd.n39 9.3005
R1645 dvdd.n48 dvdd.n47 9.3005
R1646 dvdd.n262 dvdd.n261 9.3005
R1647 dvdd.n263 dvdd.n257 9.3005
R1648 dvdd.n265 dvdd.n264 9.3005
R1649 dvdd.n266 dvdd.n243 9.3005
R1650 dvdd.n255 dvdd.n244 9.3005
R1651 dvdd.n254 dvdd.n253 9.3005
R1652 dvdd.n252 dvdd.n245 9.3005
R1653 dvdd.n251 dvdd.n250 9.3005
R1654 dvdd.n249 dvdd.n248 9.3005
R1655 dvdd.n247 dvdd.n246 9.3005
R1656 dvdd.n270 dvdd.n269 9.3005
R1657 dvdd.n275 dvdd.n274 9.3005
R1658 dvdd.n120 dvdd.n52 9.3005
R1659 dvdd.n124 dvdd.n121 9.3005
R1660 dvdd.n127 dvdd.n126 9.3005
R1661 dvdd.n128 dvdd.n119 9.3005
R1662 dvdd.n130 dvdd.n129 9.3005
R1663 dvdd.n131 dvdd.n116 9.3005
R1664 dvdd.n133 dvdd.n132 9.3005
R1665 dvdd.n134 dvdd.n115 9.3005
R1666 dvdd.n136 dvdd.n135 9.3005
R1667 dvdd.n137 dvdd.n112 9.3005
R1668 dvdd.n139 dvdd.n138 9.3005
R1669 dvdd.n140 dvdd.n111 9.3005
R1670 dvdd.n142 dvdd.n141 9.3005
R1671 dvdd.n143 dvdd.n108 9.3005
R1672 dvdd.n146 dvdd.n145 9.3005
R1673 dvdd.n147 dvdd.n107 9.3005
R1674 dvdd.n149 dvdd.n148 9.3005
R1675 dvdd.n150 dvdd.n106 9.3005
R1676 dvdd.n152 dvdd.n151 9.3005
R1677 dvdd.n153 dvdd.n105 9.3005
R1678 dvdd.n155 dvdd.n154 9.3005
R1679 dvdd.n156 dvdd.n102 9.3005
R1680 dvdd.n158 dvdd.n157 9.3005
R1681 dvdd.n159 dvdd.n53 9.3005
R1682 dvdd.n161 dvdd.n160 9.3005
R1683 dvdd.n162 dvdd.n99 9.3005
R1684 dvdd.n165 dvdd.n164 9.3005
R1685 dvdd.n166 dvdd.n98 9.3005
R1686 dvdd.n168 dvdd.n167 9.3005
R1687 dvdd.n169 dvdd.n95 9.3005
R1688 dvdd.n171 dvdd.n170 9.3005
R1689 dvdd.n172 dvdd.n94 9.3005
R1690 dvdd.n174 dvdd.n173 9.3005
R1691 dvdd.n175 dvdd.n91 9.3005
R1692 dvdd.n177 dvdd.n176 9.3005
R1693 dvdd.n178 dvdd.n90 9.3005
R1694 dvdd.n180 dvdd.n179 9.3005
R1695 dvdd.n181 dvdd.n87 9.3005
R1696 dvdd.n184 dvdd.n183 9.3005
R1697 dvdd.n185 dvdd.n86 9.3005
R1698 dvdd.n187 dvdd.n186 9.3005
R1699 dvdd.n188 dvdd.n85 9.3005
R1700 dvdd.n190 dvdd.n189 9.3005
R1701 dvdd.n191 dvdd.n84 9.3005
R1702 dvdd.n193 dvdd.n192 9.3005
R1703 dvdd.n194 dvdd.n81 9.3005
R1704 dvdd.n196 dvdd.n195 9.3005
R1705 dvdd.n197 dvdd.n54 9.3005
R1706 dvdd.n199 dvdd.n198 9.3005
R1707 dvdd.n200 dvdd.n78 9.3005
R1708 dvdd.n203 dvdd.n202 9.3005
R1709 dvdd.n204 dvdd.n77 9.3005
R1710 dvdd.n206 dvdd.n205 9.3005
R1711 dvdd.n207 dvdd.n74 9.3005
R1712 dvdd.n209 dvdd.n208 9.3005
R1713 dvdd.n210 dvdd.n73 9.3005
R1714 dvdd.n212 dvdd.n211 9.3005
R1715 dvdd.n213 dvdd.n70 9.3005
R1716 dvdd.n215 dvdd.n214 9.3005
R1717 dvdd.n216 dvdd.n69 9.3005
R1718 dvdd.n218 dvdd.n217 9.3005
R1719 dvdd.n219 dvdd.n66 9.3005
R1720 dvdd.n222 dvdd.n221 9.3005
R1721 dvdd.n223 dvdd.n65 9.3005
R1722 dvdd.n225 dvdd.n224 9.3005
R1723 dvdd.n226 dvdd.n64 9.3005
R1724 dvdd.n228 dvdd.n227 9.3005
R1725 dvdd.n229 dvdd.n63 9.3005
R1726 dvdd.n231 dvdd.n230 9.3005
R1727 dvdd.n232 dvdd.n60 9.3005
R1728 dvdd.n234 dvdd.n233 9.3005
R1729 dvdd.n235 dvdd.n55 9.3005
R1730 dvdd.n236 dvdd.n58 9.3005
R1731 dvdd.n239 dvdd.n237 9.3005
R1732 dvdd.n239 dvdd.n57 9.3005
R1733 dvdd.n241 dvdd.n240 9.3005
R1734 dvdd.n242 dvdd.n56 9.3005
R1735 dvdd.n268 dvdd.n267 9.3005
R1736 dvdd.n208 dvdd.n207 9.03579
R1737 dvdd.n170 dvdd.n169 9.03579
R1738 dvdd.n132 dvdd.n131 9.03579
R1739 dvdd.n286 dvdd.n284 7.70883
R1740 dvdd.n294 dvdd.n286 7.70883
R1741 dvdd.n287 dvdd.n285 7.70883
R1742 dvdd.n294 dvdd.n287 7.70883
R1743 dvdd.n24 dvdd.n23 7.17001
R1744 dvdd.n9 dvdd.n7 7.15376
R1745 dvdd.n283 dvdd.t144 7.14175
R1746 dvdd.n283 dvdd.t158 7.14175
R1747 dvdd.n282 dvdd.t160 7.14175
R1748 dvdd.n282 dvdd.t142 7.14175
R1749 dvdd.n289 dvdd.t150 7.14175
R1750 dvdd.n289 dvdd.t152 7.14175
R1751 dvdd.n288 dvdd.t154 7.14175
R1752 dvdd.n288 dvdd.t156 7.14175
R1753 dvdd.n250 dvdd 6.77697
R1754 dvdd.n44 dvdd.t73 6.70818
R1755 dvdd.t73 dvdd.n43 6.70818
R1756 dvdd.n32 dvdd.t145 6.70818
R1757 dvdd.t145 dvdd.n31 6.70818
R1758 dvdd dvdd.n22 6.4005
R1759 dvdd.n10 dvdd 6.4005
R1760 dvdd.n221 dvdd.n220 6.02403
R1761 dvdd.n207 dvdd.n206 6.02403
R1762 dvdd.n183 dvdd.n182 6.02403
R1763 dvdd.n169 dvdd.n168 6.02403
R1764 dvdd.n145 dvdd.n144 6.02403
R1765 dvdd.n131 dvdd.n130 6.02403
R1766 dvdd.n220 dvdd.n219 3.76521
R1767 dvdd.n182 dvdd.n181 3.76521
R1768 dvdd.n144 dvdd.n143 3.76521
R1769 dvdd.n201 dvdd.n200 3.38874
R1770 dvdd.n163 dvdd.n162 3.38874
R1771 dvdd.n125 dvdd.n124 3.38874
R1772 dvdd.n297 dvdd.n296 1.66909
R1773 dvdd.n292 dvdd.n291 1.57188
R1774 dvdd.n36 dvdd.n0 1.32907
R1775 dvdd.n2 dvdd.n0 1.32907
R1776 dvdd.n261 dvdd.n260 1.23559
R1777 dvdd.n276 dvdd.n275 0.637387
R1778 dvdd.n276 dvdd.n51 0.496845
R1779 dvdd dvdd.n268 0.438
R1780 dvdd.n50 dvdd.n49 0.432317
R1781 dvdd.n16 dvdd 0.42713
R1782 dvdd dvdd.n16 0.32387
R1783 dvdd.n268 dvdd 0.313
R1784 dvdd.n247 dvdd.n51 0.280448
R1785 dvdd.n51 dvdd 0.232271
R1786 dvdd.n7 dvdd 0.203706
R1787 dvdd.n13 dvdd 0.167167
R1788 dvdd.n19 dvdd 0.164848
R1789 dvdd.n258 dvdd 0.159538
R1790 dvdd.n38 dvdd.n15 0.141704
R1791 dvdd.n262 dvdd.n258 0.141672
R1792 dvdd.n38 dvdd.n25 0.139389
R1793 dvdd.n14 dvdd.n6 0.127236
R1794 dvdd.n264 dvdd.n243 0.120292
R1795 dvdd.n252 dvdd.n251 0.120292
R1796 dvdd.n253 dvdd.n252 0.120292
R1797 dvdd.n253 dvdd.n244 0.120292
R1798 dvdd.n121 dvdd.n120 0.120292
R1799 dvdd.n127 dvdd.n121 0.120292
R1800 dvdd.n128 dvdd.n127 0.120292
R1801 dvdd.n129 dvdd.n128 0.120292
R1802 dvdd.n129 dvdd.n116 0.120292
R1803 dvdd.n133 dvdd.n116 0.120292
R1804 dvdd.n134 dvdd.n133 0.120292
R1805 dvdd.n135 dvdd.n134 0.120292
R1806 dvdd.n135 dvdd.n112 0.120292
R1807 dvdd.n139 dvdd.n112 0.120292
R1808 dvdd.n140 dvdd.n139 0.120292
R1809 dvdd.n141 dvdd.n140 0.120292
R1810 dvdd.n141 dvdd.n108 0.120292
R1811 dvdd.n146 dvdd.n108 0.120292
R1812 dvdd.n147 dvdd.n146 0.120292
R1813 dvdd.n148 dvdd.n147 0.120292
R1814 dvdd.n148 dvdd.n106 0.120292
R1815 dvdd.n152 dvdd.n106 0.120292
R1816 dvdd.n153 dvdd.n152 0.120292
R1817 dvdd.n154 dvdd.n153 0.120292
R1818 dvdd.n154 dvdd.n102 0.120292
R1819 dvdd.n158 dvdd.n102 0.120292
R1820 dvdd.n160 dvdd.n99 0.120292
R1821 dvdd.n165 dvdd.n99 0.120292
R1822 dvdd.n166 dvdd.n165 0.120292
R1823 dvdd.n167 dvdd.n166 0.120292
R1824 dvdd.n167 dvdd.n95 0.120292
R1825 dvdd.n171 dvdd.n95 0.120292
R1826 dvdd.n172 dvdd.n171 0.120292
R1827 dvdd.n173 dvdd.n172 0.120292
R1828 dvdd.n173 dvdd.n91 0.120292
R1829 dvdd.n177 dvdd.n91 0.120292
R1830 dvdd.n178 dvdd.n177 0.120292
R1831 dvdd.n179 dvdd.n178 0.120292
R1832 dvdd.n179 dvdd.n87 0.120292
R1833 dvdd.n184 dvdd.n87 0.120292
R1834 dvdd.n185 dvdd.n184 0.120292
R1835 dvdd.n186 dvdd.n185 0.120292
R1836 dvdd.n186 dvdd.n85 0.120292
R1837 dvdd.n190 dvdd.n85 0.120292
R1838 dvdd.n191 dvdd.n190 0.120292
R1839 dvdd.n192 dvdd.n191 0.120292
R1840 dvdd.n192 dvdd.n81 0.120292
R1841 dvdd.n196 dvdd.n81 0.120292
R1842 dvdd.n198 dvdd.n78 0.120292
R1843 dvdd.n203 dvdd.n78 0.120292
R1844 dvdd.n204 dvdd.n203 0.120292
R1845 dvdd.n205 dvdd.n204 0.120292
R1846 dvdd.n205 dvdd.n74 0.120292
R1847 dvdd.n209 dvdd.n74 0.120292
R1848 dvdd.n210 dvdd.n209 0.120292
R1849 dvdd.n211 dvdd.n210 0.120292
R1850 dvdd.n211 dvdd.n70 0.120292
R1851 dvdd.n215 dvdd.n70 0.120292
R1852 dvdd.n216 dvdd.n215 0.120292
R1853 dvdd.n217 dvdd.n216 0.120292
R1854 dvdd.n217 dvdd.n66 0.120292
R1855 dvdd.n222 dvdd.n66 0.120292
R1856 dvdd.n223 dvdd.n222 0.120292
R1857 dvdd.n224 dvdd.n223 0.120292
R1858 dvdd.n224 dvdd.n64 0.120292
R1859 dvdd.n228 dvdd.n64 0.120292
R1860 dvdd.n229 dvdd.n228 0.120292
R1861 dvdd.n230 dvdd.n229 0.120292
R1862 dvdd.n230 dvdd.n60 0.120292
R1863 dvdd.n234 dvdd.n60 0.120292
R1864 dvdd.n237 dvdd.n236 0.120292
R1865 dvdd.n241 dvdd.n57 0.120292
R1866 dvdd.n242 dvdd.n241 0.120292
R1867 dvdd.n277 dvdd.n276 0.109494
R1868 dvdd.n15 dvdd.n14 0.109053
R1869 dvdd.n268 dvdd.n244 0.107271
R1870 dvdd.n14 dvdd 0.0983618
R1871 dvdd dvdd.n262 0.0981562
R1872 dvdd.n251 dvdd 0.0968542
R1873 dvdd.n281 dvdd.n280 0.0944312
R1874 dvdd.n278 dvdd.n277 0.0856755
R1875 dvdd.n279 dvdd.n278 0.0856755
R1876 dvdd.n237 dvdd 0.0812292
R1877 dvdd dvdd.n6 0.0803611
R1878 dvdd.n280 dvdd.n279 0.0777774
R1879 dvdd.n14 dvdd.n7 0.070241
R1880 dvdd.n25 dvdd.n24 0.0685285
R1881 dvdd.n268 dvdd 0.063
R1882 dvdd.n264 dvdd 0.0603958
R1883 dvdd dvdd.n263 0.0603958
R1884 dvdd.n248 dvdd 0.0603958
R1885 dvdd.n120 dvdd 0.0603958
R1886 dvdd.n159 dvdd 0.0603958
R1887 dvdd.n160 dvdd 0.0603958
R1888 dvdd.n197 dvdd 0.0603958
R1889 dvdd.n198 dvdd 0.0603958
R1890 dvdd.n235 dvdd 0.0603958
R1891 dvdd.n236 dvdd 0.0603958
R1892 dvdd.n269 dvdd 0.0603958
R1893 dvdd dvdd.n13 0.0595278
R1894 dvdd.n21 dvdd.n16 0.0535523
R1895 dvdd.n12 dvdd 0.0508472
R1896 dvdd.n291 dvdd.n290 0.0456945
R1897 dvdd.n39 dvdd.n38 0.0456858
R1898 dvdd.n20 dvdd 0.0405
R1899 dvdd dvdd.n57 0.0395625
R1900 dvdd dvdd.n297 0.0385435
R1901 dvdd dvdd.n247 0.0382604
R1902 dvdd.n39 dvdd.n0 0.0379437
R1903 dvdd.n21 dvdd 0.0339302
R1904 dvdd.n13 dvdd.n12 0.0334861
R1905 dvdd.n275 dvdd 0.03175
R1906 dvdd dvdd.n159 0.03175
R1907 dvdd dvdd.n197 0.03175
R1908 dvdd dvdd.n235 0.03175
R1909 dvdd.n269 dvdd 0.03175
R1910 dvdd.n24 dvdd.n16 0.0300191
R1911 dvdd.n248 dvdd 0.0239375
R1912 dvdd.n49 dvdd.n0 0.0233041
R1913 dvdd.n263 dvdd 0.0226354
R1914 dvdd dvdd.n158 0.0226354
R1915 dvdd dvdd.n196 0.0226354
R1916 dvdd dvdd.n234 0.0226354
R1917 dvdd dvdd.n242 0.0226354
R1918 dvdd.n299 dvdd.n298 0.0219531
R1919 dvdd.n15 dvdd 0.0210592
R1920 dvdd.n20 dvdd.n19 0.0205
R1921 dvdd.n48 dvdd.n1 0.0182365
R1922 dvdd.n25 dvdd 0.0179419
R1923 dvdd.n49 dvdd.n48 0.0151396
R1924 dvdd.n290 dvdd.n281 0.0150881
R1925 dvdd dvdd.n20 0.0121279
R1926 dvdd.n299 dvdd.n281 0.00936728
R1927 dvdd.n268 dvdd.n243 0.0083125
R1928 dvdd.n277 dvdd.t178 0.0083125
R1929 dvdd.n278 dvdd.t177 0.0083125
R1930 dvdd.n279 dvdd.t176 0.0083125
R1931 dvdd.n50 dvdd.t175 0.0083125
R1932 dvdd.n298 dvdd 0.00765103
R1933 dvdd.n280 dvdd.n50 0.00754239
R1934 dvdd.n1 dvdd 0.00176689
R1935 dvdd.n299 dvdd 0.001125
R1936 avss_ip.n264 avss_ip.n33 79101.3
R1937 avss_ip.n264 avss_ip.n34 79101.3
R1938 avss_ip.n181 avss_ip.n34 79101.3
R1939 avss_ip.n260 avss_ip.n51 63358.7
R1940 avss_ip.n260 avss_ip.n52 63358.7
R1941 avss_ip.n261 avss_ip.n52 63358.7
R1942 avss_ip.n261 avss_ip.n51 63358.7
R1943 avss_ip.t2 avss_ip.t19 58137.7
R1944 avss_ip.n221 avss_ip.n77 48722.7
R1945 avss_ip.n224 avss_ip.n77 48722.7
R1946 avss_ip.n224 avss_ip.n222 48722.7
R1947 avss_ip.n222 avss_ip.n221 48722.7
R1948 avss_ip.n111 avss_ip.n110 9309.6
R1949 avss_ip.n124 avss_ip.n111 9309.6
R1950 avss_ip.n125 avss_ip.n124 9309.6
R1951 avss_ip.n125 avss_ip.n110 9309.6
R1952 avss_ip.n280 avss_ip.n16 8357.9
R1953 avss_ip.n280 avss_ip.n17 8357.9
R1954 avss_ip.n28 avss_ip.n17 8357.9
R1955 avss_ip.n28 avss_ip.n16 8357.9
R1956 avss_ip.n166 avss_ip.n139 5804.93
R1957 avss_ip.n266 avss_ip.n13 5420.45
R1958 avss_ip.n283 avss_ip.n12 5420.45
R1959 avss_ip.n283 avss_ip.n13 5420.45
R1960 avss_ip.n157 avss_ip.n139 3720.29
R1961 avss_ip.n170 avss_ip.n168 3694.37
R1962 avss_ip.n170 avss_ip.n169 3096.92
R1963 avss_ip.n158 avss_ip.n157 3017.95
R1964 avss_ip.n156 avss_ip.n149 3007.15
R1965 avss_ip.n156 avss_ip.n150 3007.15
R1966 avss_ip.n149 avss_ip.n140 3007.15
R1967 avss_ip.n150 avss_ip.n140 3007.15
R1968 avss_ip.n138 avss_ip.n137 3007.15
R1969 avss_ip.n171 avss_ip.n138 3007.15
R1970 avss_ip.n172 avss_ip.n137 3007.15
R1971 avss_ip.n172 avss_ip.n171 3007.15
R1972 avss_ip.n165 avss_ip.n164 2708.56
R1973 avss_ip.n167 avss_ip.n166 2670.93
R1974 avss_ip.t4 avss_ip.t2 2371.94
R1975 avss_ip.t2 avss_ip.n27 2099.81
R1976 avss_ip.n168 avss_ip.n167 2073.48
R1977 avss_ip.n227 avss_ip.n74 1735.47
R1978 avss_ip.n227 avss_ip.n75 1735.47
R1979 avss_ip.n118 avss_ip.n75 1735.47
R1980 avss_ip.n118 avss_ip.n74 1735.47
R1981 avss_ip.n226 avss_ip.n225 1571.92
R1982 avss_ip.n163 avss_ip.n141 1407.97
R1983 avss_ip.n159 avss_ip.n141 1407.97
R1984 avss_ip.n163 avss_ip.n142 1407.97
R1985 avss_ip.n159 avss_ip.n142 1407.97
R1986 avss_ip.n133 avss_ip.n132 1407.97
R1987 avss_ip.n179 avss_ip.n132 1407.97
R1988 avss_ip.n178 avss_ip.n133 1407.97
R1989 avss_ip.n179 avss_ip.n178 1407.97
R1990 avss_ip.n250 avss_ip.n249 1229.9
R1991 avss_ip.n165 avss_ip.n140 1206.87
R1992 avss_ip.t2 avss_ip.n29 930.019
R1993 avss_ip.n164 avss_ip.t25 916.668
R1994 avss_ip.n158 avss_ip.t25 916.668
R1995 avss_ip.n145 avss_ip.n144 800.33
R1996 avss_ip.n144 avss_ip.n143 754.842
R1997 avss_ip.t53 avss_ip.t55 629.222
R1998 avss_ip.t0 avss_ip.t56 506.262
R1999 avss_ip.n225 avss_ip.n76 380.267
R2000 avss_ip.t56 avss_ip.n31 365.466
R2001 avss_ip.n116 avss_ip.t53 365.466
R2002 avss_ip.t2 avss_ip.n30 354.363
R2003 avss_ip.n167 avss_ip.n29 332.149
R2004 avss_ip.n180 avss_ip.n179 292.5
R2005 avss_ip.n179 avss_ip.n14 292.5
R2006 avss_ip.n178 avss_ip.n176 292.5
R2007 avss_ip.n178 avss_ip.t7 292.5
R2008 avss_ip.n175 avss_ip.n133 292.5
R2009 avss_ip.n177 avss_ip.n133 292.5
R2010 avss_ip.n134 avss_ip.n132 292.5
R2011 avss_ip.t7 avss_ip.n132 292.5
R2012 avss_ip.n160 avss_ip.n159 292.5
R2013 avss_ip.n159 avss_ip.n158 292.5
R2014 avss_ip.n161 avss_ip.n142 292.5
R2015 avss_ip.n142 avss_ip.t25 292.5
R2016 avss_ip.n163 avss_ip.n162 292.5
R2017 avss_ip.n164 avss_ip.n163 292.5
R2018 avss_ip.n147 avss_ip.n141 292.5
R2019 avss_ip.n141 avss_ip.t25 292.5
R2020 avss_ip.n173 avss_ip.n136 285.072
R2021 avss_ip.n120 avss_ip.t54 225.291
R2022 avss_ip.n174 avss_ip.n135 206.174
R2023 avss_ip.n250 avss_ip.n50 193.964
R2024 avss_ip.n155 avss_ip.n151 193.506
R2025 avss_ip.n153 avss_ip.n151 193.506
R2026 avss_ip.n152 avss_ip.n136 192.754
R2027 avss_ip.n215 avss_ip.n53 190.071
R2028 avss_ip.n258 avss_ip.n54 185.68
R2029 avss_ip.n282 avss_ip.n281 176.851
R2030 avss_ip.n266 avss_ip.n265 167.284
R2031 avss_ip.n117 avss_ip.n116 157.875
R2032 avss_ip.n27 avss_ip.n15 151.044
R2033 avss_ip.n246 avss_ip.n245 150.476
R2034 avss_ip.n247 avss_ip.n246 145.577
R2035 avss_ip.n183 avss_ip.n61 142.894
R2036 avss_ip.n263 avss_ip.n49 142.772
R2037 avss_ip.n248 avss_ip.n61 141.448
R2038 avss_ip.t4 avss_ip.n25 139.263
R2039 avss_ip.n281 avss_ip.n15 124.478
R2040 avss_ip.n166 avss_ip.n30 124.028
R2041 avss_ip.n126 avss_ip.n125 117.001
R2042 avss_ip.n125 avss_ip.n31 117.001
R2043 avss_ip.n120 avss_ip.n111 117.001
R2044 avss_ip.n116 avss_ip.n111 117.001
R2045 avss_ip.n113 avss_ip.n74 117.001
R2046 avss_ip.t17 avss_ip.n74 117.001
R2047 avss_ip.n121 avss_ip.n75 117.001
R2048 avss_ip.t17 avss_ip.n75 117.001
R2049 avss_ip.n270 avss_ip.n22 116.959
R2050 avss_ip.n184 avss_ip.n183 115.465
R2051 avss_ip.n143 avss_ip.n23 115.07
R2052 avss_ip.t3 avss_ip.t0 114.612
R2053 avss_ip.n117 avss_ip.t17 99.8107
R2054 avss_ip.n226 avss_ip.t17 99.8107
R2055 avss_ip.n119 avss_ip.n118 97.5005
R2056 avss_ip.n118 avss_ip.n117 97.5005
R2057 avss_ip.n228 avss_ip.n227 97.5005
R2058 avss_ip.n227 avss_ip.n226 97.5005
R2059 avss_ip.n151 avss_ip.n150 97.5005
R2060 avss_ip.n150 avss_ip.n139 97.5005
R2061 avss_ip.n171 avss_ip.n136 97.5005
R2062 avss_ip.n171 avss_ip.n170 97.5005
R2063 avss_ip.n173 avss_ip.n172 97.5005
R2064 avss_ip.n172 avss_ip.n24 97.5005
R2065 avss_ip.n137 avss_ip.n135 97.5005
R2066 avss_ip.n137 avss_ip.n29 97.5005
R2067 avss_ip.n153 avss_ip.n140 97.5005
R2068 avss_ip.n152 avss_ip.n138 97.5005
R2069 avss_ip.n168 avss_ip.n138 97.5005
R2070 avss_ip.n154 avss_ip.n149 97.5005
R2071 avss_ip.n149 avss_ip.n30 97.5005
R2072 avss_ip.n156 avss_ip.n155 97.5005
R2073 avss_ip.n157 avss_ip.n156 97.5005
R2074 avss_ip.n146 avss_ip.n145 96.1303
R2075 avss_ip.n161 avss_ip.n160 91.4829
R2076 avss_ip.n162 avss_ip.n161 91.4829
R2077 avss_ip.n182 avss_ip.n180 90.3013
R2078 avss_ip.n114 avss_ip.n109 88.1783
R2079 avss_ip.t4 avss_ip.n24 86.9075
R2080 avss_ip.n245 avss_ip.n62 85.4613
R2081 avss_ip.n73 avss_ip.t18 85.3972
R2082 avss_ip.n93 avss_ip.t40 85.228
R2083 avss_ip.n98 avss_ip.t46 85.228
R2084 avss_ip.t49 avss_ip.n270 85.228
R2085 avss_ip.n278 avss_ip.t43 85.228
R2086 avss_ip.n115 avss_ip.n114 84.4534
R2087 avss_ip.n102 avss_ip.n88 83.7836
R2088 avss_ip.n177 avss_ip.n26 82.7329
R2089 avss_ip.n93 avss_ip.n91 79.642
R2090 avss_ip.n123 avss_ip.n122 76.3718
R2091 avss_ip.t2 avss_ip.n31 75.5223
R2092 avss_ip.n263 avss_ip.n262 71.3439
R2093 avss_ip.n112 avss_ip.n109 69.8187
R2094 avss_ip.n247 avss_ip.n60 67.2421
R2095 avss_ip.n224 avss_ip.n223 65.2949
R2096 avss_ip.n221 avss_ip.n220 65.0005
R2097 avss_ip.n221 avss_ip.n27 65.0005
R2098 avss_ip.n225 avss_ip.n224 65.0005
R2099 avss_ip.n174 avss_ip.n173 61.1561
R2100 avss_ip.n218 avss_ip.n79 55.5405
R2101 avss_ip.n97 avss_ip.t40 54.828
R2102 avss_ip.t46 avss_ip.n97 54.828
R2103 avss_ip.n271 avss_ip.t49 54.828
R2104 avss_ip.n271 avss_ip.t43 54.828
R2105 avss_ip.n107 avss_ip.n86 52.5148
R2106 avss_ip.n48 avss_ip.n36 50.85
R2107 avss_ip.t7 avss_ip.n177 49.3364
R2108 avss_ip.t19 avss_ip.n25 46.6753
R2109 avss_ip.n183 avss_ip.t10 41.915
R2110 avss_ip.n54 avss_ip.t12 41.0016
R2111 avss_ip.n245 avss_ip.t16 41.0016
R2112 avss_ip.n249 avss_ip.t61 41.0016
R2113 avss_ip.n252 avss_ip.t59 41.0016
R2114 avss_ip.n232 avss_ip.t23 41.0016
R2115 avss_ip.n145 avss_ip.t9 40.9915
R2116 avss_ip.n143 avss_ip.t60 40.954
R2117 avss_ip.n81 avss_ip.t15 40.8142
R2118 avss_ip.n79 avss_ip.t11 40.8142
R2119 avss_ip.n103 avss_ip.t22 40.8142
R2120 avss_ip.n87 avss_ip.t1 40.8142
R2121 avss_ip.t7 avss_ip.t8 40.6077
R2122 avss_ip.n282 avss_ip.n14 39.4692
R2123 avss_ip.n36 avss_ip.t58 39.3148
R2124 avss_ip.n105 avss_ip.n104 39.3148
R2125 avss_ip.n38 avss_ip.n13 39.0005
R2126 avss_ip.t4 avss_ip.n13 39.0005
R2127 avss_ip.n12 avss_ip.n4 39.0005
R2128 avss_ip.n265 avss_ip.n12 37.5274
R2129 avss_ip.n268 avss_ip.n4 37.3029
R2130 avss_ip.n91 avss_ip.n22 35.8089
R2131 avss_ip.n274 avss_ip.n273 34.0856
R2132 avss_ip.n279 avss_ip.n278 33.8591
R2133 avss_ip.n184 avss_ip.n182 32.622
R2134 avss_ip.n251 avss_ip.n250 32.583
R2135 avss_ip.n169 avss_ip.n24 32.2586
R2136 avss_ip.n272 avss_ip.n271 30.4005
R2137 avss_ip.n97 avss_ip.n96 30.4005
R2138 avss_ip.n229 avss_ip.n228 27.3252
R2139 avss_ip.n267 avss_ip.n23 27.0857
R2140 avss_ip.n82 avss_ip.n80 27.0817
R2141 avss_ip.n268 avss_ip.n267 25.4655
R2142 avss_ip.n91 avss_ip.t57 25.2421
R2143 avss_ip.n153 avss_ip.n152 24.5522
R2144 avss_ip.n69 avss_ip.t32 23.0489
R2145 avss_ip.n89 avss_ip.t47 20.9512
R2146 avss_ip.n92 avss_ip.t41 20.9512
R2147 avss_ip.n89 avss_ip.t48 20.9512
R2148 avss_ip.n92 avss_ip.t42 20.9512
R2149 avss_ip.n4 avss_ip.t26 20.9512
R2150 avss_ip.n38 avss_ip.t30 20.9512
R2151 avss_ip.n19 avss_ip.t44 20.9512
R2152 avss_ip.n21 avss_ip.t50 20.9512
R2153 avss_ip.n19 avss_ip.t45 20.9512
R2154 avss_ip.n21 avss_ip.t51 20.9512
R2155 avss_ip.n209 avss_ip.n208 20.2706
R2156 avss_ip.n96 avss_ip.n16 20.1729
R2157 avss_ip.n26 avss_ip.n16 20.1729
R2158 avss_ip.n272 avss_ip.n17 20.1729
R2159 avss_ip.n26 avss_ip.n17 20.1729
R2160 avss_ip.n267 avss_ip.n266 19.5005
R2161 avss_ip.n284 avss_ip.n283 19.5005
R2162 avss_ip.n283 avss_ip.n282 19.5005
R2163 avss_ip.n69 avss_ip.n68 18.9164
R2164 avss_ip.n69 avss_ip.n67 18.6458
R2165 avss_ip.n41 avss_ip.n40 18.4564
R2166 avss_ip.n289 avss_ip.n5 18.4545
R2167 avss_ip.n288 avss_ip.n6 18.4545
R2168 avss_ip.n42 avss_ip.n39 18.4545
R2169 avss_ip.n38 avss_ip.n23 17.0186
R2170 avss_ip.n215 avss_ip.n80 16.8541
R2171 avss_ip.n4 avss_ip.n3 16.8187
R2172 avss_ip.n38 avss_ip.n37 16.8187
R2173 avss_ip.n284 avss_ip.n11 16.2478
R2174 avss_ip.n217 avss_ip.n80 16.1777
R2175 avss_ip.n152 avss_ip.n135 16.0656
R2176 avss_ip.n285 avss_ip.n10 16.016
R2177 avss_ip.n154 avss_ip.n153 15.9156
R2178 avss_ip.n155 avss_ip.n154 15.9156
R2179 avss_ip.n105 avss_ip.n102 15.4672
R2180 avss_ip.n279 avss_ip.n18 14.7511
R2181 avss_ip.n262 avss_ip.n50 14.7129
R2182 avss_ip.n28 avss_ip.n22 14.3687
R2183 avss_ip.n280 avss_ip.n279 13.9291
R2184 avss_ip.n281 avss_ip.n280 13.9291
R2185 avss_ip.t19 avss_ip.n28 13.9291
R2186 avss_ip.n81 avss_ip.n18 12.0635
R2187 avss_ip.n176 avss_ip.n175 12.0186
R2188 avss_ip.n155 avss_ip.n148 11.8074
R2189 avss_ip.n162 avss_ip.n146 11.6811
R2190 avss_ip.n223 avss_ip.n54 11.6159
R2191 avss_ip.n106 avss_ip.n88 11.0473
R2192 avss_ip.n45 avss_ip.n44 10.9678
R2193 avss_ip.n115 avss_ip.n113 10.5881
R2194 avss_ip.n249 avss_ip.n248 10.4547
R2195 avss_ip.n76 avss_ip.n34 10.3497
R2196 avss_ip.n229 avss_ip.n64 10.0473
R2197 avss_ip.n123 avss_ip.n112 9.92203
R2198 avss_ip.n113 avss_ip.n73 9.90239
R2199 avss_ip.n122 avss_ip.n120 9.7605
R2200 avss_ip.n61 avss_ip.n34 9.59066
R2201 avss_ip.n144 avss_ip.n33 9.59066
R2202 avss_ip.n33 avss_ip.n32 9.58979
R2203 avss_ip.n122 avss_ip.n121 9.33884
R2204 avss_ip.n270 avss_ip.n21 9.33383
R2205 avss_ip.n272 avss_ip.n21 9.33383
R2206 avss_ip.n278 avss_ip.n19 9.33383
R2207 avss_ip.n174 avss_ip.n134 9.32519
R2208 avss_ip.n48 avss_ip.n47 9.28796
R2209 avss_ip.n51 avss_ip.n10 9.28621
R2210 avss_ip.n51 avss_ip.n15 9.28621
R2211 avss_ip.n246 avss_ip.n52 9.28621
R2212 avss_ip.n76 avss_ip.n52 9.28621
R2213 avss_ip.n119 avss_ip.n115 9.25764
R2214 avss_ip.n232 avss_ip.n64 9.21481
R2215 avss_ip.n208 avss_ip.n197 9.12258
R2216 avss_ip.n108 avss_ip.n107 8.98751
R2217 avss_ip.n209 avss_ip.n108 8.93556
R2218 avss_ip.t8 avss_ip.n14 8.72915
R2219 avss_ip.n121 avss_ip.n73 8.69884
R2220 avss_ip.t3 avss_ip.t55 8.34965
R2221 avss_ip.n216 avss_ip.n214 7.9153
R2222 avss_ip.n114 avss_ip.n110 7.8005
R2223 avss_ip.n110 avss_ip.t55 7.8005
R2224 avss_ip.n124 avss_ip.n123 7.8005
R2225 avss_ip.n124 avss_ip.t55 7.8005
R2226 avss_ip.n259 avss_ip.n53 7.67034
R2227 avss_ip.n244 avss_ip.n64 7.2005
R2228 avss_ip.n275 avss_ip.n4 6.94429
R2229 avss_ip.n220 avss_ip.n219 6.85764
R2230 avss_ip.n147 avss_ip.n146 6.76005
R2231 avss_ip.n274 avss_ip.n19 5.92871
R2232 avss_ip.n130 avss_ip.n129 5.2694
R2233 avss_ip.n127 avss_ip.n126 4.63427
R2234 avss_ip.n243 avss_ip.n62 4.58032
R2235 avss_ip.n148 avss_ip.n147 4.53239
R2236 avss_ip.n98 avss_ip.n78 4.24039
R2237 avss_ip.n129 avss_ip.n63 4.17857
R2238 avss_ip.t4 avss_ip.n26 4.17507
R2239 avss_ip.n3 avss_ip.t27 4.133
R2240 avss_ip.n3 avss_ip.t39 4.133
R2241 avss_ip.n5 avss_ip.t6 4.133
R2242 avss_ip.n5 avss_ip.t28 4.133
R2243 avss_ip.n6 avss_ip.t36 4.133
R2244 avss_ip.n6 avss_ip.t21 4.133
R2245 avss_ip.n40 avss_ip.t20 4.133
R2246 avss_ip.n40 avss_ip.t37 4.133
R2247 avss_ip.n39 avss_ip.t38 4.133
R2248 avss_ip.n39 avss_ip.t5 4.133
R2249 avss_ip.n37 avss_ip.t62 4.133
R2250 avss_ip.n37 avss_ip.t29 4.133
R2251 avss_ip.n67 avss_ip.t13 4.133
R2252 avss_ip.n67 avss_ip.t14 4.133
R2253 avss_ip.n68 avss_ip.t24 4.133
R2254 avss_ip.n68 avss_ip.t31 4.133
R2255 avss_ip.n134 avss_ip.n131 4.08638
R2256 avss_ip.n93 avss_ip.n92 4.06187
R2257 avss_ip.n96 avss_ip.n89 4.06187
R2258 avss_ip.n98 avss_ip.n89 4.06187
R2259 avss_ip.n176 avss_ip.n131 3.72833
R2260 avss_ip.n96 avss_ip.n90 3.66019
R2261 avss_ip.n219 avss_ip.n18 3.45272
R2262 avss_ip.n274 avss_ip.n272 3.40563
R2263 avss_ip.n102 avss_ip.n101 3.36563
R2264 avss_ip.n45 avss_ip.n11 3.15412
R2265 avss_ip.n218 avss_ip.n217 3.09777
R2266 avss_ip.n223 avss_ip.n62 2.80936
R2267 avss_ip.n175 avss_ip.n174 2.59291
R2268 avss_ip.n112 avss_ip.n77 2.5005
R2269 avss_ip.n77 avss_ip.t0 2.5005
R2270 avss_ip.n222 avss_ip.n53 2.5005
R2271 avss_ip.n222 avss_ip.t0 2.5005
R2272 avss_ip.n94 avss_ip.n93 2.35984
R2273 avss_ip.n270 avss_ip.n269 2.33555
R2274 avss_ip.n278 avss_ip.n277 2.3255
R2275 avss_ip.n272 avss_ip.n20 2.3255
R2276 avss_ip.n96 avss_ip.n95 2.3255
R2277 avss_ip.n99 avss_ip.n98 2.3255
R2278 avss_ip.n262 avss_ip.n261 2.30365
R2279 avss_ip.n261 avss_ip.t3 2.30365
R2280 avss_ip.n260 avss_ip.n259 2.30365
R2281 avss_ip.t3 avss_ip.n260 2.30365
R2282 avss_ip.n259 avss_ip.n258 2.18463
R2283 avss_ip.n169 avss_ip.n25 1.99449
R2284 avss_ip.n160 avss_ip.n148 1.88285
R2285 avss_ip.n190 avss_ip.n128 1.864
R2286 avss_ip.n128 avss_ip.n9 1.79647
R2287 avss_ip.n197 avss_ip.n127 1.77712
R2288 avss_ip.n181 avss_ip.n32 1.73666
R2289 avss_ip.n182 avss_ip.n181 1.73641
R2290 avss_ip.n264 avss_ip.n263 1.73641
R2291 avss_ip.t2 avss_ip.n264 1.73641
R2292 avss_ip.n213 avss_ip.n82 1.68005
R2293 avss_ip.n46 avss_ip.n35 1.66407
R2294 avss_ip.n86 avss_ip.n84 1.55377
R2295 avss_ip.n245 avss_ip.n63 1.55139
R2296 avss_ip.n233 avss_ip.n232 1.5505
R2297 avss_ip.n36 avss_ip.n35 1.5505
R2298 avss_ip.n253 avss_ip.n252 1.5505
R2299 avss_ip.n249 avss_ip.n59 1.5505
R2300 avss_ip.n65 avss_ip.n54 1.5505
R2301 avss_ip.n214 avss_ip.n213 1.5505
R2302 avss_ip.n104 avss_ip.n84 1.5505
R2303 avss_ip.n254 avss_ip.n253 1.38009
R2304 avss_ip.n245 avss_ip.n244 1.36564
R2305 avss_ip.n130 avss_ip.n58 1.308
R2306 avss_ip.n189 avss_ip.n186 1.308
R2307 avss_ip.n191 avss_ip.n190 1.298
R2308 avss_ip.n188 avss_ip.n55 1.298
R2309 avss_ip.n255 avss_ip.n254 1.298
R2310 avss_ip.n207 avss_ip.n72 1.26349
R2311 avss_ip.n219 avss_ip.n218 1.23599
R2312 avss_ip.n265 avss_ip.t4 1.2046
R2313 avss_ip.n292 avss_ip.n291 0.96015
R2314 avss_ip.n216 avss_ip.n215 0.890856
R2315 avss_ip.n256 avss_ip.n56 0.705502
R2316 avss_ip.n244 avss_ip.n243 0.705087
R2317 avss_ip.n166 avss_ip.n165 0.611283
R2318 avss_ip.n186 avss_ip.n128 0.60099
R2319 avss_ip.n189 avss_ip.n188 0.573464
R2320 avss_ip.n44 avss_ip.n43 0.570043
R2321 avss_ip.n212 avss_ip.n83 0.565252
R2322 avss_ip.n256 avss_ip.n255 0.564213
R2323 avss_ip.n71 avss_ip.n57 0.563097
R2324 avss_ip.n193 avss_ip.n192 0.561311
R2325 avss_ip.n254 avss_ip.n58 0.56102
R2326 avss_ip.n190 avss_ip.n189 0.553102
R2327 avss_ip.n290 avss_ip.n4 0.542817
R2328 avss_ip.n194 avss_ip.n85 0.519771
R2329 avss_ip.n195 avss_ip.n56 0.469362
R2330 avss_ip.n273 avss_ip.n8 0.4655
R2331 avss_ip.n11 avss_ip.n9 0.4655
R2332 avss_ip.n275 avss_ip.n274 0.460631
R2333 avss_ip.n269 avss_ip.n268 0.424176
R2334 avss_ip.n204 avss_ip.n200 0.419057
R2335 avss_ip.n205 avss_ip.n198 0.402572
R2336 avss_ip.n92 avss_ip.n90 0.402174
R2337 avss_ip.n43 avss_ip.n2 0.365261
R2338 avss_ip.n211 avss_ip.n210 0.356091
R2339 avss_ip.n186 avss_ip.n185 0.331536
R2340 avss_ip.n273 avss_ip.n10 0.325138
R2341 avss_ip.n70 avss_ip.n69 0.32382
R2342 avss_ip avss_ip.n0 0.311796
R2343 avss_ip.n101 avss_ip.n100 0.3105
R2344 avss_ip.n206 avss_ip.n1 0.298814
R2345 avss_ip.n188 avss_ip.n187 0.295466
R2346 avss_ip.n185 avss_ip.n130 0.287418
R2347 avss_ip.n7 avss_ip.n2 0.284875
R2348 avss_ip.n255 avss_ip.n57 0.284284
R2349 avss_ip.n191 avss_ip.n83 0.284284
R2350 avss_ip.n192 avss_ip.n55 0.282595
R2351 avss_ip.n193 avss_ip.n191 0.27809
R2352 avss_ip.n291 avss_ip.n290 0.273938
R2353 avss_ip.n187 avss_ip.n58 0.273407
R2354 avss_ip.n101 avss_ip.n78 0.259356
R2355 avss_ip.n220 avss_ip.n78 0.252717
R2356 avss_ip.n71 avss_ip.n65 0.245995
R2357 avss_ip.n180 avss_ip.n131 0.225293
R2358 avss_ip.n192 avss_ip.n56 0.207375
R2359 avss_ip.n257 avss_ip.n256 0.203564
R2360 avss_ip.n103 avss_ip.n88 0.177831
R2361 avss_ip.n88 avss_ip.n87 0.177831
R2362 avss_ip.n228 avss_ip.n73 0.177123
R2363 avss_ip.n126 avss_ip.n109 0.177123
R2364 avss_ip.n286 avss_ip.n8 0.176218
R2365 avss_ip.n286 avss_ip.n9 0.169383
R2366 avss_ip.n242 avss_ip.n65 0.167129
R2367 avss_ip.n47 avss_ip.n46 0.162784
R2368 avss_ip.n0 avss_ip 0.160253
R2369 avss_ip.n49 avss_ip.n35 0.157831
R2370 avss_ip.n257 avss_ip.n55 0.155905
R2371 avss_ip.n99 avss_ip.n0 0.15494
R2372 avss_ip.n194 avss_ip.n193 0.154875
R2373 avss_ip.n85 avss_ip.n83 0.154875
R2374 avss_ip.n210 avss_ip.n85 0.154406
R2375 avss_ip.n231 avss_ip.n71 0.153625
R2376 avss_ip.n72 avss_ip.n57 0.153625
R2377 avss_ip.n213 avss_ip.n212 0.152809
R2378 avss_ip.n251 avss_ip.n60 0.151816
R2379 avss_ip.n217 avss_ip.n216 0.146497
R2380 avss_ip.n240 avss_ip.n239 0.141572
R2381 avss_ip.n100 avss_ip.n84 0.135688
R2382 avss_ip.n269 avss_ip.n20 0.133352
R2383 avss_ip.n204 avss_ip.n203 0.126796
R2384 avss_ip.n230 avss_ip.n72 0.126776
R2385 avss_ip.n129 avss_ip.n59 0.124652
R2386 avss_ip.n277 avss_ip.n276 0.119062
R2387 avss_ip.n107 avss_ip.n106 0.106958
R2388 avss_ip.n211 avss_ip.n84 0.106495
R2389 avss_ip.n212 avss_ip.n211 0.1055
R2390 avss_ip.n100 avss_ip.n99 0.0992461
R2391 avss_ip.n94 avss_ip.n90 0.0916765
R2392 avss_ip.n240 avss_ip.n236 0.0874565
R2393 avss_ip.n46 avss_ip.n9 0.0871299
R2394 avss_ip.n291 avss_ip.n2 0.0816897
R2395 avss_ip.n237 avss_ip.t64 0.0794225
R2396 avss_ip.n207 avss_ip.n206 0.0783908
R2397 avss_ip.n238 avss_ip.n237 0.0770981
R2398 avss_ip.n239 avss_ip.n238 0.0770981
R2399 avss_ip.n243 avss_ip.n242 0.0743095
R2400 avss_ip.n236 avss_ip.n70 0.072538
R2401 avss_ip.n290 avss_ip.n289 0.0725156
R2402 avss_ip.n43 avss_ip.n42 0.071218
R2403 avss_ip.n289 avss_ip.n288 0.0688391
R2404 avss_ip.n42 avss_ip.n41 0.0688391
R2405 avss_ip.n233 avss_ip.n231 0.0659262
R2406 avss_ip.n196 avss_ip.n194 0.0640417
R2407 avss_ip.n106 avss_ip.n105 0.0601701
R2408 avss_ip.n276 avss_ip.n275 0.058625
R2409 avss_ip.n203 avss_ip.n198 0.0560826
R2410 avss_ip.n197 avss_ip.n196 0.0545698
R2411 avss_ip.n234 avss_ip.n233 0.0519706
R2412 avss_ip.n210 avss_ip.n209 0.0505
R2413 avss_ip.n285 avss_ip.n284 0.0468768
R2414 avss_ip.n292 avss_ip.n1 0.0468062
R2415 avss_ip.n120 avss_ip.n119 0.0462143
R2416 avss_ip.n196 avss_ip.n195 0.0450312
R2417 avss_ip.n206 avss_ip.n205 0.0421667
R2418 avss_ip.n108 avss_ip.n1 0.0402436
R2419 avss_ip avss_ip.n292 0.0386424
R2420 avss_ip.n249 avss_ip.n60 0.0350946
R2421 avss_ip.n286 avss_ip.n285 0.0349444
R2422 avss_ip.n41 avss_ip.n7 0.0344533
R2423 avss_ip.n288 avss_ip.n287 0.0340208
R2424 avss_ip.n44 avss_ip.n38 0.0332283
R2425 avss_ip.n252 avss_ip.n251 0.0328933
R2426 avss_ip.n287 avss_ip.n286 0.0295323
R2427 avss_ip.n95 avss_ip.n94 0.0286593
R2428 avss_ip.n195 avss_ip.n127 0.0283443
R2429 avss_ip.n49 avss_ip.n48 0.0262964
R2430 avss_ip.n276 avss_ip.n20 0.0248405
R2431 avss_ip.n231 avss_ip.n230 0.0238343
R2432 avss_ip.n234 avss_ip.n70 0.023
R2433 avss_ip.n241 avss_ip.n240 0.0219286
R2434 avss_ip.n199 avss_ip.t52 0.0199669
R2435 avss_ip.n205 avss_ip.n204 0.0199236
R2436 avss_ip.n201 avss_ip.t33 0.0197446
R2437 avss_ip.n236 avss_ip.n235 0.0187186
R2438 avss_ip.n235 avss_ip.n66 0.0182821
R2439 avss_ip.n95 avss_ip.n0 0.0171896
R2440 avss_ip.n208 avss_ip.n207 0.0163974
R2441 avss_ip.n277 avss_ip.n8 0.016031
R2442 avss_ip.n47 avss_ip.n45 0.0159589
R2443 avss_ip.n202 avss_ip.n201 0.0128949
R2444 avss_ip.n201 avss_ip.t34 0.0124791
R2445 avss_ip.n199 avss_ip.t35 0.0121969
R2446 avss_ip.n187 avss_ip.n50 0.0107423
R2447 avss_ip.n202 avss_ip.n200 0.0106706
R2448 avss_ip.n66 avss_ip.n63 0.0105375
R2449 avss_ip.n258 avss_ip.n257 0.0101473
R2450 avss_ip.n230 avss_ip.n229 0.00985614
R2451 avss_ip.n241 avss_ip.n66 0.00826231
R2452 avss_ip.n104 avss_ip.n103 0.00639018
R2453 avss_ip.n214 avss_ip.n79 0.00639018
R2454 avss_ip.n82 avss_ip.n81 0.00639018
R2455 avss_ip.n87 avss_ip.n86 0.00639018
R2456 avss_ip.n248 avss_ip.n247 0.00637916
R2457 avss_ip.n185 avss_ip.n184 0.00414706
R2458 avss_ip.n237 avss_ip.t63 0.00282438
R2459 avss_ip.n238 avss_ip.t66 0.00282438
R2460 avss_ip.n239 avss_ip.t65 0.00282438
R2461 avss_ip.n242 avss_ip.n241 0.00157066
R2462 avss_ip.n287 avss_ip.n7 0.00136505
R2463 avss_ip.t2 avss_ip.n32 0.00121043
R2464 avss_ip.n253 avss_ip.n59 0.00106561
R2465 avss_ip.n200 avss_ip.n199 0.00103899
R2466 avss_ip.n235 avss_ip.n234 0.00080012
R2467 avss_ip.n201 avss_ip.n198 0.000704348
R2468 avss_ip.n203 avss_ip.n202 0.000704348
R2469 a_9120_n9346.n1 a_9120_n9346.t2 649.659
R2470 a_9120_n9346.n0 a_9120_n9346.t4 227.685
R2471 a_9120_n9346.t0 a_9120_n9346.n2 44.6806
R2472 a_9120_n9346.n1 a_9120_n9346.t1 5.45407
R2473 a_9120_n9346.n0 a_9120_n9346.t3 5.07473
R2474 a_9120_n9346.n2 a_9120_n9346.n0 0.639781
R2475 a_9120_n9346.n2 a_9120_n9346.n1 0.0621233
R2476 ibias.n7 ibias.n1 1544.9
R2477 ibias.n4 ibias.n3 1544.9
R2478 ibias.n2 ibias.n0 300.425
R2479 ibias.n8 ibias.n2 300.425
R2480 ibias.n9 ibias.n0 177.746
R2481 ibias.n9 ibias.n8 177.746
R2482 ibias.n5 ibias.n1 139.143
R2483 ibias.n6 ibias.n3 139.143
R2484 ibias.n9 ibias.t1 60.1061
R2485 ibias.n4 ibias.n0 46.2505
R2486 ibias.n8 ibias.n7 46.2505
R2487 ibias.n5 ibias.n4 40.8622
R2488 ibias.n7 ibias.n6 40.8622
R2489 ibias.n3 ibias.n2 12.3338
R2490 ibias.n9 ibias.n1 12.3338
R2491 ibias.n6 ibias.t0 4.16651
R2492 ibias.t0 ibias.n5 4.16651
R2493 ibias ibias.n9 1.58676
R2494 avdd_ip.n81 avdd_ip.n73 58547.9
R2495 avdd_ip.n81 avdd_ip.n80 58547.9
R2496 avdd_ip.n79 avdd_ip.n73 58547.9
R2497 avdd_ip.n80 avdd_ip.n79 58547.9
R2498 avdd_ip.n43 avdd_ip.n42 54381
R2499 avdd_ip.n82 avdd_ip.n71 28978.4
R2500 avdd_ip.n82 avdd_ip.n72 28978.4
R2501 avdd_ip.n78 avdd_ip.n71 28978.4
R2502 avdd_ip.n78 avdd_ip.n72 28978.4
R2503 avdd_ip.n93 avdd_ip.n26 7296
R2504 avdd_ip.n91 avdd_ip.n26 7296
R2505 avdd_ip.n93 avdd_ip.n27 7296
R2506 avdd_ip.n91 avdd_ip.n27 7296
R2507 avdd_ip.n77 avdd_ip.n75 5062.04
R2508 avdd_ip.n75 avdd_ip.n74 3209.98
R2509 avdd_ip.n76 avdd_ip.n62 1005.14
R2510 avdd_ip.n44 avdd_ip.n36 857.648
R2511 avdd_ip.n40 avdd_ip.n37 857.648
R2512 avdd_ip.n44 avdd_ip.n37 857.648
R2513 avdd_ip.n55 avdd_ip.n54 857.648
R2514 avdd_ip.n57 avdd_ip.n50 857.648
R2515 avdd_ip.n43 avdd_ip.t3 337.433
R2516 avdd_ip.n77 avdd_ip.n76 269.44
R2517 avdd_ip.n57 avdd_ip.n56 267.182
R2518 avdd_ip.n54 avdd_ip.n51 267.182
R2519 avdd_ip.n41 avdd_ip.n40 267.182
R2520 avdd_ip.n84 avdd_ip.n63 212.139
R2521 avdd_ip.n90 avdd_ip.n89 202.696
R2522 avdd_ip.n88 avdd_ip.n29 134.065
R2523 avdd_ip.n74 avdd_ip.n29 110.358
R2524 avdd_ip.t5 avdd_ip.n26 105.665
R2525 avdd_ip.t9 avdd_ip.n27 105.665
R2526 avdd_ip.n85 avdd_ip.n84 96.3051
R2527 avdd_ip.n58 avdd_ip.n57 92.5005
R2528 avdd_ip.n55 avdd_ip.n49 92.5005
R2529 avdd_ip.n54 avdd_ip.n53 92.5005
R2530 avdd_ip.n52 avdd_ip.n50 92.5005
R2531 avdd_ip.n45 avdd_ip.n44 92.5005
R2532 avdd_ip.n44 avdd_ip.n43 92.5005
R2533 avdd_ip.n38 avdd_ip.n37 92.5005
R2534 avdd_ip.t3 avdd_ip.n37 92.5005
R2535 avdd_ip.n40 avdd_ip.n39 92.5005
R2536 avdd_ip.n36 avdd_ip.n35 92.5005
R2537 avdd_ip.n39 avdd_ip.n35 91.4862
R2538 avdd_ip.n53 avdd_ip.n49 91.4829
R2539 avdd_ip.n92 avdd_ip.t5 79.5673
R2540 avdd_ip.n92 avdd_ip.t9 79.5673
R2541 avdd_ip.n85 avdd_ip.n62 73.3959
R2542 avdd_ip.n39 avdd_ip.n38 66.8321
R2543 avdd_ip.n53 avdd_ip.n52 66.3131
R2544 avdd_ip.n59 avdd_ip.n49 63.936
R2545 avdd_ip.n46 avdd_ip.n35 63.936
R2546 avdd_ip.n2 avdd_ip.t4 62.0945
R2547 avdd_ip.n17 avdd_ip.t20 61.1041
R2548 avdd_ip.n15 avdd_ip.t21 60.1061
R2549 avdd_ip.n14 avdd_ip.t25 60.1061
R2550 avdd_ip.n21 avdd_ip.t19 60.1061
R2551 avdd_ip.n24 avdd_ip.t24 60.1061
R2552 avdd_ip.n89 avdd_ip.t13 60.1061
R2553 avdd_ip.n89 avdd_ip.t10 60.1061
R2554 avdd_ip.n89 avdd_ip.t11 60.1061
R2555 avdd_ip.n63 avdd_ip.t8 60.1061
R2556 avdd_ip.n63 avdd_ip.t6 60.1061
R2557 avdd_ip.n63 avdd_ip.t7 60.1061
R2558 avdd_ip.n31 avdd_ip.t14 60.1061
R2559 avdd_ip.n31 avdd_ip.t12 60.1061
R2560 avdd_ip.n30 avdd_ip.t16 60.1061
R2561 avdd_ip.n30 avdd_ip.t15 60.1061
R2562 avdd_ip.n65 avdd_ip.t23 60.1061
R2563 avdd_ip.n65 avdd_ip.t17 60.1061
R2564 avdd_ip.n64 avdd_ip.t26 60.1061
R2565 avdd_ip.n64 avdd_ip.t18 60.1061
R2566 avdd_ip.n16 avdd_ip.t22 60.1061
R2567 avdd_ip.n41 avdd_ip.n36 57.4849
R2568 avdd_ip.n56 avdd_ip.n55 57.4849
R2569 avdd_ip.n51 avdd_ip.n50 57.4849
R2570 avdd_ip.n2 avdd_ip.n1 55.1707
R2571 avdd_ip.n2 avdd_ip.n0 54.9038
R2572 avdd_ip.n69 avdd_ip.n13 44.6614
R2573 avdd_ip.n58 avdd_ip.n48 43.3376
R2574 avdd_ip.n45 avdd_ip.n34 43.3376
R2575 avdd_ip.n83 avdd_ip.n70 30.1747
R2576 avdd_ip.n51 avdd_ip.t28 28.8172
R2577 avdd_ip.n56 avdd_ip.t28 28.8172
R2578 avdd_ip.t3 avdd_ip.n41 28.8172
R2579 avdd_ip.n90 avdd_ip.n28 10.6324
R2580 avdd_ip.n74 avdd_ip.n25 8.37369
R2581 avdd_ip.n16 avdd_ip.n15 7.25561
R2582 avdd_ip.n0 avdd_ip.t0 6.92425
R2583 avdd_ip.n0 avdd_ip.t2 6.92425
R2584 avdd_ip.n1 avdd_ip.t27 6.92425
R2585 avdd_ip.n1 avdd_ip.t1 6.92425
R2586 avdd_ip.n91 avdd_ip.n90 6.37981
R2587 avdd_ip.n92 avdd_ip.n91 6.37981
R2588 avdd_ip.n94 avdd_ip.n93 6.37981
R2589 avdd_ip.n93 avdd_ip.n92 6.37981
R2590 avdd_ip.n24 avdd_ip.n23 6.17839
R2591 avdd_ip.n78 avdd_ip.n77 6.15262
R2592 avdd_ip.n94 avdd_ip.n25 5.31953
R2593 avdd_ip.n52 avdd_ip.n48 4.38907
R2594 avdd_ip.n38 avdd_ip.n34 4.38907
R2595 avdd_ip.n95 avdd_ip.n94 3.87825
R2596 avdd_ip.n84 avdd_ip.n83 3.6009
R2597 avdd_ip.n60 avdd_ip.n48 2.4925
R2598 avdd_ip.n47 avdd_ip.n34 2.44611
R2599 avdd_ip.n29 avdd_ip.n27 2.43471
R2600 avdd_ip.n70 avdd_ip.n26 2.43471
R2601 avdd_ip.n59 avdd_ip.n58 2.37764
R2602 avdd_ip.n46 avdd_ip.n45 2.37764
R2603 avdd_ip.n60 avdd_ip.n59 2.3255
R2604 avdd_ip.n47 avdd_ip.n46 2.3255
R2605 avdd_ip.n22 avdd_ip.n21 1.87566
R2606 avdd_ip.n95 avdd_ip.n13 1.41891
R2607 avdd_ip.n4 avdd_ip.n3 1.18871
R2608 avdd_ip.n23 avdd_ip.n14 1.07773
R2609 avdd_ip.n79 avdd_ip.n78 1.05764
R2610 avdd_ip.n83 avdd_ip.n82 1.05764
R2611 avdd_ip.n82 avdd_ip.n81 1.05764
R2612 avdd_ip.n86 avdd_ip.n85 1.02375
R2613 avdd_ip.n21 avdd_ip.n20 0.982678
R2614 avdd_ip.n20 avdd_ip.n14 0.919312
R2615 avdd_ip.n17 avdd_ip.n16 0.90347
R2616 avdd_ip.n23 avdd_ip.n22 0.845955
R2617 avdd_ip.n11 avdd_ip.n4 0.827286
R2618 avdd_ip avdd_ip.n11 0.808179
R2619 avdd_ip.n66 avdd_ip.n64 0.65712
R2620 avdd_ip.n32 avdd_ip.n30 0.652725
R2621 avdd_ip.n88 avdd_ip.n87 0.613954
R2622 avdd_ip.n76 avdd_ip.n72 0.530586
R2623 avdd_ip.n80 avdd_ip.n72 0.530586
R2624 avdd_ip.n75 avdd_ip.n71 0.530586
R2625 avdd_ip.n73 avdd_ip.n71 0.530586
R2626 avdd_ip.n3 avdd_ip.n2 0.507794
R2627 avdd_ip.n70 avdd_ip.n69 0.448948
R2628 avdd_ip.n19 avdd_ip.n18 0.402976
R2629 avdd_ip.n33 avdd_ip.n32 0.319749
R2630 avdd_ip.n87 avdd_ip.n86 0.319015
R2631 avdd_ip.n67 avdd_ip.n66 0.319015
R2632 avdd_ip.n18 avdd_ip.n12 0.319015
R2633 avdd_ip.n20 avdd_ip.n19 0.282318
R2634 avdd_ip.n11 avdd_ip.n10 0.255087
R2635 avdd_ip.n32 avdd_ip.n31 0.25137
R2636 avdd_ip.n66 avdd_ip.n65 0.25137
R2637 avdd_ip.n96 avdd_ip.n12 0.243945
R2638 avdd_ip avdd_ip.n97 0.213307
R2639 avdd_ip.n87 avdd_ip.n28 0.211864
R2640 avdd_ip.n18 avdd_ip.n17 0.211864
R2641 avdd_ip.n97 avdd_ip 0.18211
R2642 avdd_ip.n25 avdd_ip.n24 0.174542
R2643 avdd_ip.n15 avdd_ip.n13 0.174542
R2644 avdd_ip.n62 avdd_ip.n61 0.166571
R2645 avdd_ip.n67 avdd_ip.n12 0.150396
R2646 avdd_ip.n86 avdd_ip.n33 0.150396
R2647 avdd_ip.n3 avdd_ip.t33 0.125045
R2648 avdd_ip.n7 avdd_ip.n4 0.123905
R2649 avdd_ip.n68 avdd_ip.n33 0.117461
R2650 avdd_ip.n10 avdd_ip.n9 0.111971
R2651 avdd_ip.n8 avdd_ip.n7 0.110265
R2652 avdd_ip.n68 avdd_ip.n67 0.108384
R2653 avdd_ip.n6 avdd_ip.n5 0.106696
R2654 avdd_ip.n9 avdd_ip.n8 0.106696
R2655 avdd_ip.n61 avdd_ip.n47 0.0839309
R2656 avdd_ip.n61 avdd_ip.n60 0.0812962
R2657 avdd_ip.n5 avdd_ip.t30 0.0180781
R2658 avdd_ip.n9 avdd_ip.t32 0.0180781
R2659 avdd_ip.n8 avdd_ip.t29 0.0180781
R2660 avdd_ip.n6 avdd_ip.t31 0.0180781
R2661 avdd_ip.n10 avdd_ip.n5 0.0174228
R2662 avdd_ip.n96 avdd_ip.n95 0.0173478
R2663 avdd_ip.n63 avdd_ip.n28 0.0154184
R2664 avdd_ip.n89 avdd_ip.n88 0.0154184
R2665 avdd_ip.n7 avdd_ip.n6 0.0150053
R2666 avdd_ip.n69 avdd_ip.n68 0.0108333
R2667 avdd_ip.n97 avdd_ip.n96 0.00292843
R2668 avdd_ip.n22 avdd_ip.n19 0.000885802
R2669 xout.n29 xout.t26 594.784
R2670 xout.n29 xout.t24 194.649
R2671 xout.n25 xout.t23 124.457
R2672 xout.n25 xout.t25 106.793
R2673 xout.t23 xout.n24 86.3125
R2674 xout.t25 xout.n23 86.3125
R2675 xout.n3 xout.t15 62.0071
R2676 xout.n4 xout.t13 62.0071
R2677 xout.n3 xout.t20 60.1061
R2678 xout.n4 xout.t21 60.1061
R2679 xout.n8 xout.t11 60.1061
R2680 xout.n8 xout.t10 60.1061
R2681 xout.n10 xout.t14 60.1061
R2682 xout.n10 xout.t12 60.1061
R2683 xout.n0 xout.t17 60.1061
R2684 xout.n0 xout.t19 60.1061
R2685 xout.n1 xout.t16 60.1061
R2686 xout.n1 xout.t18 60.1061
R2687 xout.n24 xout.n23 58.6245
R2688 xout.n22 xout.t2 43.5339
R2689 xout.n28 xout.n27 21.3269
R2690 xout.n16 xout.n15 18.5533
R2691 xout.n20 xout.n13 18.553
R2692 xout.n19 xout.n18 18.4723
R2693 xout.n19 xout.n17 18.4564
R2694 xout.n16 xout.n14 18.4564
R2695 xout.n27 xout.n23 12.2455
R2696 xout.n18 xout.t5 4.133
R2697 xout.n18 xout.t6 4.133
R2698 xout.n17 xout.t4 4.133
R2699 xout.n17 xout.t3 4.133
R2700 xout.n15 xout.t0 4.133
R2701 xout.n15 xout.t22 4.133
R2702 xout.n14 xout.t7 4.133
R2703 xout.n14 xout.t8 4.133
R2704 xout.n13 xout.t9 4.133
R2705 xout.n13 xout.t1 4.133
R2706 xout.n5 xout.n4 3.64406
R2707 xout.n5 xout.n3 3.61238
R2708 xout.n26 xout.n24 3.56553
R2709 xout.n22 xout.n21 2.24362
R2710 xout.n29 xout.n28 2.18092
R2711 xout.n28 xout.n22 1.03102
R2712 xout.n27 xout.n26 0.742745
R2713 xout.n26 xout.n25 0.715885
R2714 xout.n21 xout.n12 0.464586
R2715 xout.n2 xout.n0 0.424187
R2716 xout.n11 xout.n9 0.402558
R2717 xout xout.n29 0.377063
R2718 xout.n6 xout.n2 0.316998
R2719 xout.n2 xout.n1 0.310571
R2720 xout.n12 xout.n7 0.273717
R2721 xout.n7 xout.n6 0.261913
R2722 xout.n9 xout.n8 0.254998
R2723 xout.n11 xout.n10 0.25137
R2724 xout.n6 xout.n5 0.143668
R2725 xout.n9 xout.n7 0.126918
R2726 xout.n12 xout.n11 0.125886
R2727 xout.n21 xout.n20 0.0947164
R2728 xout.n20 xout.n16 0.0657574
R2729 xout.n20 xout.n19 0.0480746
R2730 inv_in.n19 inv_in.t0 47.4896
R2731 inv_in.n18 inv_in.t3 6.48745
R2732 inv_in.n19 inv_in.t1 6.24255
R2733 inv_in inv_in.n17 2.2182
R2734 inv_in.n18 inv_in 0.342687
R2735 inv_in inv_in.n18 0.217687
R2736 inv_in.n5 inv_in.n4 0.110198
R2737 inv_in.n7 inv_in.n6 0.110101
R2738 inv_in.n10 inv_in.n9 0.110101
R2739 inv_in.n8 inv_in.n2 0.110101
R2740 inv_in.n16 inv_in.n15 0.109734
R2741 inv_in.n14 inv_in.n0 0.109734
R2742 inv_in.n13 inv_in.n12 0.109709
R2743 inv_in.n11 inv_in.n1 0.109709
R2744 inv_in.n9 inv_in.n7 0.109325
R2745 inv_in.n9 inv_in.n8 0.109325
R2746 inv_in.n12 inv_in.n11 0.109325
R2747 inv_in.n11 inv_in.n3 0.109325
R2748 inv_in.n15 inv_in.n14 0.1086
R2749 inv_in.n16 inv_in.n0 0.1086
R2750 inv_in.n4 inv_in.n3 0.10222
R2751 inv_in.n7 inv_in.n5 0.101755
R2752 inv_in inv_in.n19 0.09425
R2753 inv_in.n18 inv_in 0.063
R2754 inv_in.n0 inv_in.t11 0.00880157
R2755 inv_in.n7 inv_in.t9 0.00848368
R2756 inv_in.n9 inv_in.t10 0.00848368
R2757 inv_in.n8 inv_in.t2 0.00848368
R2758 inv_in.n5 inv_in.t12 0.00838586
R2759 inv_in.n4 inv_in.t14 0.0083125
R2760 inv_in.n6 inv_in.t13 0.0083125
R2761 inv_in.n2 inv_in.t6 0.0083125
R2762 inv_in.n10 inv_in.t4 0.0083125
R2763 inv_in.n1 inv_in.t5 0.0083125
R2764 inv_in.n13 inv_in.t8 0.0083125
R2765 inv_in.n17 inv_in.t7 0.0083125
R2766 inv_in.n6 inv_in.n3 0.00106244
R2767 inv_in.n12 inv_in.n2 0.00106244
R2768 inv_in.n11 inv_in.n10 0.00106244
R2769 inv_in.n17 inv_in.n16 0.000989074
R2770 inv_in.n15 inv_in.n1 0.000548907
R2771 inv_in.n14 inv_in.n13 0.000548907
R2772 avss.n20 avss.n19 18580.7
R2773 avss.n38 avss.n37 15308.7
R2774 avss.n76 avss.n20 12246.6
R2775 avss.n40 avss.n35 3599.36
R2776 avss.n41 avss.n35 3599.36
R2777 avss.n41 avss.n34 3599.36
R2778 avss.n40 avss.n34 3599.36
R2779 avss.n67 avss.n25 2489.59
R2780 avss.n67 avss.n26 2489.59
R2781 avss.n69 avss.n26 2489.59
R2782 avss.n69 avss.n25 2489.59
R2783 avss.n28 avss.n21 2489.59
R2784 avss.n28 avss.n22 2489.59
R2785 avss.n74 avss.n22 2489.59
R2786 avss.n74 avss.n21 2489.59
R2787 avss.n78 avss.n13 2489.59
R2788 avss.n78 avss.n14 2489.59
R2789 avss.n16 avss.n14 2489.59
R2790 avss.n16 avss.n13 2489.59
R2791 avss.n88 avss.n6 2489.59
R2792 avss.n90 avss.n6 2489.59
R2793 avss.n90 avss.n5 2489.59
R2794 avss.n88 avss.n5 2489.59
R2795 avss.n36 avss.n20 2342.14
R2796 avss.n77 avss.n76 930.542
R2797 avss.n76 avss.n75 930.542
R2798 avss.n43 avss.n42 881.42
R2799 avss.n19 avss.t6 633.244
R2800 avss.n15 avss.t4 633.244
R2801 avss.t22 avss.n17 633.244
R2802 avss.n77 avss.t24 633.244
R2803 avss.n75 avss.t8 633.244
R2804 avss.n29 avss.t10 633.244
R2805 avss.t0 avss.n30 633.244
R2806 avss.n37 avss.t2 633.244
R2807 avss.t20 avss.n36 412.863
R2808 avss.t18 avss.n38 397.358
R2809 avss.n17 avss.n15 362.704
R2810 avss.n30 avss.n29 362.704
R2811 avss.t12 avss.t20 306.255
R2812 avss.t14 avss.t12 306.255
R2813 avss.t14 avss.t16 306.255
R2814 avss.t16 avss.t18 306.255
R2815 avss.n39 avss.n32 295.807
R2816 avss.n66 avss.n65 289.13
R2817 avss.n87 avss.n3 289.13
R2818 avss.n92 avss.n91 288.753
R2819 avss.n70 avss.n24 288.753
R2820 avss.n89 avss.t6 234.865
R2821 avss.n89 avss.t4 234.865
R2822 avss.n18 avss.t22 234.865
R2823 avss.t24 avss.n18 234.865
R2824 avss.n27 avss.t8 234.865
R2825 avss.t10 avss.n27 234.865
R2826 avss.n68 avss.t0 234.865
R2827 avss.n68 avss.t2 234.865
R2828 avss.n31 avss.n10 152.73
R2829 avss.n73 avss.n72 152.73
R2830 avss.n80 avss.n7 152.73
R2831 avss.n79 avss.n12 152.73
R2832 avss.n39 avss.n33 118.081
R2833 avss.n91 avss.n4 103.529
R2834 avss.n64 avss.n31 103.529
R2835 avss.n72 avss.n71 103.529
R2836 avss.n66 avss.n64 103.529
R2837 avss.n71 avss.n70 103.529
R2838 avss.n86 avss.n7 103.529
R2839 avss.n12 avss.n4 103.529
R2840 avss.n87 avss.n86 103.529
R2841 avss.n88 avss.n87 97.5005
R2842 avss.n89 avss.n88 97.5005
R2843 avss.n91 avss.n90 97.5005
R2844 avss.n90 avss.n89 97.5005
R2845 avss.n13 avss.n7 97.5005
R2846 avss.n18 avss.n13 97.5005
R2847 avss.n14 avss.n12 97.5005
R2848 avss.n18 avss.n14 97.5005
R2849 avss.n31 avss.n21 97.5005
R2850 avss.n27 avss.n21 97.5005
R2851 avss.n72 avss.n22 97.5005
R2852 avss.n27 avss.n22 97.5005
R2853 avss.n70 avss.n69 97.5005
R2854 avss.n69 avss.n68 97.5005
R2855 avss.n67 avss.n66 97.5005
R2856 avss.n68 avss.n67 97.5005
R2857 avss.n42 avss.n33 69.8003
R2858 avss.n38 avss.n35 54.5071
R2859 avss.n5 avss.n3 48.7505
R2860 avss.n19 avss.n5 48.7505
R2861 avss.n8 avss.n6 48.7505
R2862 avss.n15 avss.n6 48.7505
R2863 avss.n16 avss.n8 48.7505
R2864 avss.n17 avss.n16 48.7505
R2865 avss.n79 avss.n78 48.7505
R2866 avss.n78 avss.n77 48.7505
R2867 avss.n74 avss.n73 48.7505
R2868 avss.n75 avss.n74 48.7505
R2869 avss.n28 avss.n23 48.7505
R2870 avss.n29 avss.n28 48.7505
R2871 avss.n25 avss.n23 48.7505
R2872 avss.n30 avss.n25 48.7505
R2873 avss.n65 avss.n26 48.7505
R2874 avss.n37 avss.n26 48.7505
R2875 avss.n40 avss.n39 45.0005
R2876 avss.t14 avss.n40 45.0005
R2877 avss.n42 avss.n41 45.0005
R2878 avss.n41 avss.t14 45.0005
R2879 avss.n64 avss.n63 40.3697
R2880 avss.n71 avss.n23 40.3697
R2881 avss.n86 avss.n85 40.3697
R2882 avss.n8 avss.n4 40.3697
R2883 avss.n94 avss.n1 39.7977
R2884 avss.n34 avss.n33 39.0005
R2885 avss.n36 avss.n34 39.0005
R2886 avss.n35 avss.n32 39.0005
R2887 avss.n94 avss 33.7505
R2888 avss.n84 avss.t23 29.9199
R2889 avss.n62 avss.t1 29.9199
R2890 avss.n62 avss.t11 29.9199
R2891 avss.n84 avss.t5 29.9199
R2892 avss.n2 avss.t7 29.798
R2893 avss.n57 avss.t3 29.798
R2894 avss.n11 avss.t25 29.798
R2895 avss.n11 avss.t9 29.798
R2896 avss.n32 avss.t19 20.9512
R2897 avss.n46 avss.n45 18.8362
R2898 avss.n46 avss.n44 18.6458
R2899 avss.n44 avss.t15 4.133
R2900 avss.n44 avss.t17 4.133
R2901 avss.n45 avss.t21 4.133
R2902 avss.n45 avss.t13 4.133
R2903 avss.n47 avss.n43 1.61679
R2904 avss.n55 avss 1.33946
R2905 avss.n58 avss.n24 1.21803
R2906 avss.n93 avss.n92 1.21803
R2907 avss.n54 avss.n47 0.8655
R2908 avss.n63 avss.n62 0.664786
R2909 avss.n81 avss.n10 0.664786
R2910 avss.n81 avss.n80 0.664786
R2911 avss.n85 avss.n84 0.664786
R2912 avss.n55 avss.n54 0.53175
R2913 avss.n56 avss.n9 0.434977
R2914 avss.n95 avss.n0 0.433066
R2915 avss.n61 avss.n59 0.433066
R2916 avss.n61 avss.n60 0.433066
R2917 avss.n60 avss.n0 0.433066
R2918 avss.n65 avss.n24 0.376971
R2919 avss.n92 avss.n3 0.376971
R2920 avss.n84 avss.n0 0.299413
R2921 avss.n62 avss.n61 0.299413
R2922 avss.n62 avss.n9 0.247783
R2923 avss.n84 avss.n83 0.247783
R2924 avss.n83 avss 0.245943
R2925 avss.n59 avss.n58 0.231236
R2926 avss.n82 avss.n9 0.201672
R2927 avss.n83 avss.n82 0.201672
R2928 avss.n2 avss.n1 0.2005
R2929 avss.n95 avss.n94 0.2005
R2930 avss.n47 avss.n46 0.1855
R2931 avss.n49 avss.n48 0.122162
R2932 avss.n82 avss.n81 0.120904
R2933 avss.n50 avss.n49 0.105544
R2934 avss.n51 avss.n50 0.101695
R2935 avss.n73 avss.n10 0.1005
R2936 avss.n80 avss.n79 0.1005
R2937 avss.n60 avss.n11 0.0997647
R2938 avss.n53 avss.n48 0.0989292
R2939 avss.n56 avss.n55 0.096886
R2940 avss.n54 avss.n53 0.0847138
R2941 avss.n63 avss.n23 0.0825513
R2942 avss.n85 avss.n8 0.0825513
R2943 avss.n51 avss.n48 0.0586846
R2944 avss.n57 avss.n56 0.0480171
R2945 avss avss.n95 0.0332586
R2946 avss.n59 avss 0.0330342
R2947 avss.n94 avss.n93 0.0328276
R2948 avss.n43 avss.n32 0.0328232
R2949 avss.n53 avss.n52 0.0277801
R2950 avss.n50 avss.t28 0.0083125
R2951 avss.n49 avss.t29 0.0083125
R2952 avss.n48 avss.t26 0.0083125
R2953 avss.n52 avss.t27 0.0083125
R2954 avss avss.n1 0.00342969
R2955 avss.n93 avss.n2 0.000931034
R2956 avss.n58 avss.n57 0.000928082
R2957 avss.n81 avss.n11 0.000683824
R2958 avss.n52 avss.n51 0.000622332
R2959 avdd.n92 avdd.n91 15807.9
R2960 avdd.n93 avdd.n92 15807.9
R2961 avdd.n93 avdd.n28 15807.9
R2962 avdd.n91 avdd.n28 15807.9
R2963 avdd.n90 avdd.n27 8112.97
R2964 avdd.n94 avdd.n27 8112.97
R2965 avdd.n94 avdd.n26 8112.97
R2966 avdd.n90 avdd.n26 8112.97
R2967 avdd.n98 avdd.n6 2166
R2968 avdd.n97 avdd.n6 2166
R2969 avdd.n98 avdd.n7 2166
R2970 avdd.n97 avdd.n7 2166
R2971 avdd.n78 avdd.n77 1643.17
R2972 avdd.n77 avdd.n76 1643.17
R2973 avdd.n74 avdd.n69 1643.17
R2974 avdd.n80 avdd.n69 1643.17
R2975 avdd.n52 avdd.n37 1643.17
R2976 avdd.n60 avdd.n37 1643.17
R2977 avdd.n55 avdd.n54 1643.17
R2978 avdd.n58 avdd.n55 1643.17
R2979 avdd.n89 avdd.n88 1439.4
R2980 avdd.n89 avdd.n29 1352.37
R2981 avdd.n66 avdd.n25 1313.54
R2982 avdd.n71 avdd.n70 1106.59
R2983 avdd.n70 avdd.n68 1106.59
R2984 avdd.n40 avdd.n39 1106.59
R2985 avdd.n39 avdd.n36 1106.59
R2986 avdd.n78 avdd.n68 536.587
R2987 avdd.n76 avdd.n71 536.587
R2988 avdd.n74 avdd.n71 536.587
R2989 avdd.n80 avdd.n68 536.587
R2990 avdd.n52 avdd.n40 536.587
R2991 avdd.n54 avdd.n40 536.587
R2992 avdd.n58 avdd.n36 536.587
R2993 avdd.n60 avdd.n36 536.587
R2994 avdd.n75 avdd.t6 382.582
R2995 avdd.n79 avdd.t6 382.582
R2996 avdd.n53 avdd.t4 382.582
R2997 avdd.n59 avdd.t4 382.582
R2998 avdd.n73 avdd.n30 319.248
R2999 avdd.n57 avdd.n56 319.248
R3000 avdd.n88 avdd.n31 287.265
R3001 avdd.n38 avdd.n29 287.265
R3002 avdd.n88 avdd.n30 276.295
R3003 avdd.n56 avdd.n29 276.295
R3004 avdd.n86 avdd.t7 227.377
R3005 avdd.n1 avdd.t15 227.377
R3006 avdd.n34 avdd.t10 227.377
R3007 avdd.n43 avdd.t5 227.377
R3008 avdd.n66 avdd.n3 205.554
R3009 avdd.n72 avdd.n31 189.742
R3010 avdd.n38 avdd.n35 189.742
R3011 avdd.n101 avdd.n3 186.73
R3012 avdd.t13 avdd.n6 157.492
R3013 avdd.t11 avdd.n7 157.492
R3014 avdd.n25 avdd.n4 118.862
R3015 avdd.n100 avdd.n4 115.031
R3016 avdd.n73 avdd.n72 108.569
R3017 avdd.n57 avdd.n35 108.569
R3018 avdd.t2 avdd.t13 107.677
R3019 avdd.t0 avdd.t2 107.677
R3020 avdd.t0 avdd.t8 107.677
R3021 avdd.t8 avdd.t11 107.677
R3022 avdd.n62 avdd.n5 63.4672
R3023 avdd.n23 avdd.t14 60.1061
R3024 avdd.n21 avdd.n20 54.9038
R3025 avdd.n21 avdd.n19 54.9038
R3026 avdd.n72 avdd.n2 32.2138
R3027 avdd.n61 avdd.n35 32.2138
R3028 avdd.n101 avdd.n100 31.7005
R3029 avdd.n102 avdd.n101 30.3938
R3030 avdd.n76 avdd.n73 26.4291
R3031 avdd.n76 avdd.n75 26.4291
R3032 avdd.n74 avdd.n2 26.4291
R3033 avdd.n75 avdd.n74 26.4291
R3034 avdd.n78 avdd.n32 26.4291
R3035 avdd.n79 avdd.n78 26.4291
R3036 avdd.n81 avdd.n80 26.4291
R3037 avdd.n80 avdd.n79 26.4291
R3038 avdd.n58 avdd.n57 26.4291
R3039 avdd.n59 avdd.n58 26.4291
R3040 avdd.n61 avdd.n60 26.4291
R3041 avdd.n60 avdd.n59 26.4291
R3042 avdd.n54 avdd.n41 26.4291
R3043 avdd.n54 avdd.n53 26.4291
R3044 avdd.n52 avdd.n51 26.4291
R3045 avdd.n53 avdd.n52 26.4291
R3046 avdd.n96 avdd.n24 15.6997
R3047 avdd.n97 avdd.n96 14.2313
R3048 avdd.t0 avdd.n97 14.2313
R3049 avdd.n99 avdd.n98 14.2313
R3050 avdd.n98 avdd.t0 14.2313
R3051 avdd.n77 avdd.n30 13.2148
R3052 avdd.n77 avdd.t6 13.2148
R3053 avdd.n70 avdd.n31 13.2148
R3054 avdd.n70 avdd.t6 13.2148
R3055 avdd.n69 avdd.n3 13.2148
R3056 avdd.t6 avdd.n69 13.2148
R3057 avdd.n39 avdd.n38 13.2148
R3058 avdd.n39 avdd.t4 13.2148
R3059 avdd.n56 avdd.n55 13.2148
R3060 avdd.n55 avdd.t4 13.2148
R3061 avdd.n49 avdd.n37 13.2148
R3062 avdd.t4 avdd.n37 13.2148
R3063 avdd.n7 avdd.n4 12.3338
R3064 avdd.n47 avdd.n6 12.3338
R3065 avdd.n100 avdd.n99 8.13132
R3066 avdd.n95 avdd.n25 7.54184
R3067 avdd.n82 avdd.n32 7.30037
R3068 avdd.n46 avdd.n41 7.22016
R3069 avdd.n20 avdd.t3 6.92425
R3070 avdd.n20 avdd.t1 6.92425
R3071 avdd.n19 avdd.t9 6.92425
R3072 avdd.n19 avdd.t12 6.92425
R3073 avdd.n48 avdd.n47 6.88003
R3074 avdd.n99 avdd.n5 6.16704
R3075 avdd.n67 avdd.n66 3.51587
R3076 avdd.n50 avdd.n49 3.30818
R3077 avdd.n82 avdd.n81 2.8599
R3078 avdd.n90 avdd.n89 2.84665
R3079 avdd.n91 avdd.n90 2.84665
R3080 avdd.n95 avdd.n94 2.84665
R3081 avdd.n94 avdd.n93 2.84665
R3082 avdd.n51 avdd.n46 2.78239
R3083 avdd.n48 avdd.n5 2.51338
R3084 avdd.n49 avdd.n48 2.33395
R3085 avdd.n67 avdd.n27 2.28445
R3086 avdd.n92 avdd.n27 2.28445
R3087 avdd.n50 avdd.n26 2.28445
R3088 avdd.n28 avdd.n26 2.28445
R3089 avdd.n84 avdd 1.89829
R3090 avdd.n23 avdd.n22 1.87575
R3091 avdd.n102 avdd.n2 1.70717
R3092 avdd.n62 avdd.n61 1.70717
R3093 avdd.n81 avdd.n67 1.56476
R3094 avdd.n51 avdd.n50 1.54047
R3095 avdd.n85 avdd.n1 1.11161
R3096 avdd.n96 avdd.n95 1.03878
R3097 avdd.n65 avdd.n33 0.909856
R3098 avdd.n87 avdd.n65 0.871595
R3099 avdd.n42 avdd.n29 0.517167
R3100 avdd.n63 avdd.n62 0.517167
R3101 avdd.n103 avdd.n102 0.517167
R3102 avdd.n88 avdd.n87 0.517167
R3103 avdd.n83 avdd.n1 0.457832
R3104 avdd.n88 avdd.n32 0.30326
R3105 avdd.n41 avdd.n29 0.29856
R3106 avdd.n44 avdd.n34 0.277965
R3107 avdd.n44 avdd.n43 0.242141
R3108 avdd.n13 avdd.n12 0.221624
R3109 avdd.n45 avdd.n44 0.191202
R3110 avdd.n15 avdd.n8 0.171
R3111 avdd.n64 avdd 0.165618
R3112 avdd.n18 avdd.n8 0.158572
R3113 avdd.n45 avdd.n33 0.155105
R3114 avdd.n22 avdd.n18 0.129984
R3115 avdd.n65 avdd.n64 0.124867
R3116 avdd.n24 avdd.n23 0.0960224
R3117 avdd.n18 avdd.n17 0.0860931
R3118 avdd.n16 avdd.n15 0.0718577
R3119 avdd.n15 avdd.n14 0.0677409
R3120 avdd.n46 avdd.n45 0.058264
R3121 avdd.n83 avdd.n82 0.058264
R3122 avdd.n86 avdd.n85 0.0482015
R3123 avdd avdd.n63 0.0421667
R3124 avdd avdd.n0 0.035342
R3125 avdd.n12 avdd.n0 0.0293462
R3126 avdd.n22 avdd.n21 0.0285269
R3127 avdd.n17 avdd.n16 0.0255438
R3128 avdd.n14 avdd.n13 0.0253723
R3129 avdd.n12 avdd.n8 0.0246031
R3130 avdd.n85 avdd.n84 0.0240664
R3131 avdd.n11 avdd.t18 0.0122401
R3132 avdd avdd.n103 0.0122337
R3133 avdd.n17 avdd.t16 0.0122173
R3134 avdd.n10 avdd.t19 0.0113908
R3135 avdd.n9 avdd.t17 0.011362
R3136 avdd.n63 avdd.n34 0.0105575
R3137 avdd.n103 avdd.n1 0.0105575
R3138 avdd.n17 avdd.n9 0.00991802
R3139 avdd.n11 avdd.n10 0.00930403
R3140 avdd.n47 avdd.n24 0.00805162
R3141 avdd.n64 avdd 0.00600766
R3142 avdd.n43 avdd.n42 0.00573256
R3143 avdd.n42 avdd.n33 0.00515116
R3144 avdd.n87 avdd.n86 0.00333375
R3145 avdd.n14 avdd.n9 0.00220261
R3146 avdd.n16 avdd.n10 0.00176706
R3147 avdd.n84 avdd.n83 0.00111075
R3148 avdd.n64 avdd.n0 0.00109866
R3149 avdd.n13 avdd.n11 0.000671533
R3150 standby.n1 standby.t0 260.322
R3151 standby.n0 standby.t1 194.635
R3152 standby.n1 standby.t2 175.169
R3153 standby.n2 standby.n1 152
R3154 standby.n2 standby.n0 69.674
R3155 standby standby.n2 1.55726
R3156 standby.n0 standby 0.748625
R3157 x3.out_b.n5 x3.out_b.t8 397.163
R3158 x3.out_b.n3 x3.out_b.t4 397.163
R3159 x3.out_b.n6 x3.out_b.t8 396.286
R3160 x3.out_b.n4 x3.out_b.t4 396.286
R3161 x3.out_b.t3 x3.out_b.n5 375.649
R3162 x3.out_b.n6 x3.out_b.t3 375.649
R3163 x3.out_b.n0 x3.out_b.t6 375.649
R3164 x3.out_b.n7 x3.out_b.t6 375.649
R3165 x3.out_b.t7 x3.out_b.n3 375.649
R3166 x3.out_b.n4 x3.out_b.t7 375.649
R3167 x3.out_b.n2 x3.out_b.t2 227.887
R3168 x3.out_b.n2 x3.out_b.n8 25.0905
R3169 x3.out_b.n5 x3.out_b.n0 21.5154
R3170 x3.out_b.n3 x3.out_b.n0 21.1069
R3171 x3.out_b.n7 x3.out_b.n4 20.6372
R3172 x3.out_b.n7 x3.out_b.n6 20.6372
R3173 x3.out_b.n2 x3.out_b.t5 12.777
R3174 x3.out_b.n8 x3.out_b.t0 5.5105
R3175 x3.out_b.n8 x3.out_b.t1 5.5105
R3176 x3.out_b.n1 x3.out_b.n0 5.32901
R3177 x3.out_b.n1 x3.out_b.n7 2.74252
R3178 x3.out_b.n2 x3.out_b.n1 1.06508
R3179 ena.n0 ena.t2 260.322
R3180 ena.n2 ena.t0 194.63
R3181 ena.n0 ena.t1 175.169
R3182 ena.n1 ena.n0 152
R3183 ena.n3 ena.n2 51.6747
R3184 ena ena.n3 4.94983
R3185 ena.n3 ena.n1 3.45996
R3186 ena.n1 ena 1.55726
R3187 ena.n2 ena 0.746125
R3188 vg1.n10 vg1.t2 85.228
R3189 vg1.n0 vg1.t1 61.1305
R3190 vg1.n7 vg1.t5 54.828
R3191 vg1.n7 vg1.t2 54.828
R3192 vg1.n5 vg1.t0 42.6599
R3193 vg1.n8 vg1.n7 32.9015
R3194 vg1.n10 vg1.n9 30.9745
R3195 vg1.n9 vg1.t3 20.9512
R3196 vg1.n6 vg1.n5 3.63479
R3197 vg1.n11 vg1.n10 2.3255
R3198 vg1.n12 vg1.n0 0.471594
R3199 vg1.n5 vg1.n4 0.390524
R3200 vg1.n9 vg1.n8 0.238607
R3201 vg1.n11 vg1.n6 0.176742
R3202 vg1 vg1.n12 0.133236
R3203 vg1.n1 vg1.t9 0.0767969
R3204 vg1.n2 vg1.n1 0.0752537
R3205 vg1.n3 vg1.n2 0.0752537
R3206 vg1.n4 vg1.t8 0.0717511
R3207 vg1.n0 vg1 0.0387813
R3208 vg1.n12 vg1.n11 0.0257152
R3209 vg1.n8 vg1.n6 0.0123355
R3210 vg1.n4 vg1.n3 0.00554581
R3211 vg1.n1 vg1.t4 0.00204321
R3212 vg1.n2 vg1.t7 0.00204321
R3213 vg1.n3 vg1.t6 0.00204321
R3214 xin.n36 xin.t8 594.832
R3215 xin.t18 xin.n5 380.808
R3216 xin.n6 xin.t18 380.808
R3217 xin.n6 xin.t15 380.611
R3218 xin.t15 xin.n5 380.611
R3219 xin.t13 xin.n7 380.611
R3220 xin.n8 xin.t13 380.611
R3221 xin.t19 xin.n4 380.611
R3222 xin.n9 xin.t19 380.611
R3223 xin.n11 xin.t16 380.611
R3224 xin.t16 xin.n10 380.611
R3225 xin.n12 xin.t11 380.611
R3226 xin.t11 xin.n3 380.611
R3227 xin.t10 xin.n13 380.611
R3228 xin.n14 xin.t10 380.611
R3229 xin.t17 xin.n2 380.611
R3230 xin.n15 xin.t17 380.611
R3231 xin.n17 xin.t14 380.611
R3232 xin.t14 xin.n16 380.611
R3233 xin.n18 xin.t12 380.611
R3234 xin.t12 xin.n1 380.611
R3235 xin.t9 xin.n19 380.611
R3236 xin.n20 xin.t9 380.611
R3237 xin.n21 xin.t6 380.611
R3238 xin.t6 xin.n0 380.611
R3239 xin.n36 xin.t21 194.639
R3240 xin.n25 xin.t20 124.457
R3241 xin.n25 xin.t7 106.793
R3242 xin.t7 xin.n23 86.3125
R3243 xin.t20 xin.n24 86.3125
R3244 xin.n24 xin.n23 58.6245
R3245 xin.n30 xin.t0 45.927
R3246 xin.n28 xin.n27 20.1298
R3247 xin.n27 xin.n23 12.2455
R3248 xin.n35 xin.n34 4.04311
R3249 xin.n26 xin.n24 3.56553
R3250 xin.n34 xin.n29 3.51336
R3251 xin.n30 xin.n29 3.51061
R3252 xin.n28 xin.n22 1.95915
R3253 xin.n35 xin.n28 1.1106
R3254 xin.n22 xin.n21 0.8105
R3255 xin.n22 xin.n0 0.7905
R3256 xin.n27 xin.n26 0.741791
R3257 xin.n26 xin.n25 0.715885
R3258 xin.n36 xin.n35 0.4755
R3259 xin xin.n36 0.377063
R3260 xin.n8 xin.n5 0.198
R3261 xin.n9 xin.n8 0.198
R3262 xin.n10 xin.n9 0.198
R3263 xin.n10 xin.n3 0.198
R3264 xin.n14 xin.n3 0.198
R3265 xin.n15 xin.n14 0.198
R3266 xin.n16 xin.n15 0.198
R3267 xin.n16 xin.n1 0.198
R3268 xin.n20 xin.n1 0.198
R3269 xin.n21 xin.n20 0.198
R3270 xin.n7 xin.n6 0.198
R3271 xin.n7 xin.n4 0.198
R3272 xin.n11 xin.n4 0.198
R3273 xin.n12 xin.n11 0.198
R3274 xin.n13 xin.n12 0.198
R3275 xin.n13 xin.n2 0.198
R3276 xin.n17 xin.n2 0.198
R3277 xin.n18 xin.n17 0.198
R3278 xin.n19 xin.n18 0.198
R3279 xin.n19 xin.n0 0.198
R3280 xin.t4 xin.t2 0.0760058
R3281 xin.n31 xin.n30 0.0410952
R3282 xin.n32 xin.n29 0.0410952
R3283 xin.n34 xin.n33 0.0410952
R3284 xin.n32 xin.t5 0.0264927
R3285 xin.n31 xin.t1 0.0264885
R3286 xin.n33 xin.t4 0.0264703
R3287 xin.n33 xin.t3 0.0264296
R3288 xin.t3 xin.n32 0.0264114
R3289 xin.t5 xin.n31 0.0264072
R3290 vg2.n2 vg2.t9 87.8852
R3291 vg2.n9 vg2.t5 87.8852
R3292 vg2.n5 vg2.t6 85.228
R3293 vg2.n12 vg2.t7 85.228
R3294 vg2.n15 vg2.t8 67.0783
R3295 vg2.n4 vg2.t9 54.828
R3296 vg2.t6 vg2.n4 54.828
R3297 vg2.n11 vg2.t5 54.828
R3298 vg2.t7 vg2.n11 54.828
R3299 vg2.n16 vg2.t0 42.6015
R3300 vg2.n4 vg2.n3 30.4005
R3301 vg2.n11 vg2.n10 30.4005
R3302 vg2.n3 vg2.n1 29.1205
R3303 vg2.n5 vg2.n1 29.1205
R3304 vg2.n10 vg2.n8 29.1205
R3305 vg2.n12 vg2.n8 29.1205
R3306 vg2.n6 vg2.n5 2.3255
R3307 vg2.n13 vg2.n12 2.3255
R3308 vg2.n3 vg2.n2 2.13477
R3309 vg2.n10 vg2.n9 2.13477
R3310 vg2 vg2.n14 0.742464
R3311 vg2.n16 vg2.n15 0.714193
R3312 vg2.n14 vg2.n6 0.474719
R3313 vg2.n14 vg2.n13 0.474719
R3314 vg2.n1 vg2.n0 0.423227
R3315 vg2.n8 vg2.n7 0.423227
R3316 vg2.n2 vg2.n0 0.308459
R3317 vg2.n9 vg2.n7 0.308459
R3318 vg2.n6 vg2.n0 0.284875
R3319 vg2.n13 vg2.n7 0.284875
R3320 vg2.n15 vg2.t3 0.170134
R3321 vg2 vg2.n16 0.119455
R3322 vg2.t1 vg2.t2 0.0652716
R3323 vg2.t4 vg2.t1 0.0652716
R3324 vg2.t3 vg2.t4 0.0652716
R3325 vrb.n2 vrb.t0 43.1048
R3326 vrb.n0 vrb.t4 22.3777
R3327 vrb.n1 vrb.t1 22.1989
R3328 vrb.n1 vrb.t3 21.3671
R3329 vrb.n0 vrb.t2 21.3663
R3330 vrb.n3 vrb.n2 1.11856
R3331 vrb.n3 vrb.n0 0.759192
R3332 vrb.n2 vrb.n1 0.758408
R3333 vrb vrb.n3 0.0491111
R3334 x3.out.n3 x3.out.t6 393.144
R3335 x3.out.n5 x3.out.t7 393.144
R3336 x3.out.n4 x3.out.t6 391.815
R3337 x3.out.t7 x3.out.n2 391.815
R3338 x3.out.n5 x3.out.t4 371.31
R3339 x3.out.t4 x3.out.n2 371.31
R3340 x3.out.t3 x3.out.n1 371.31
R3341 x3.out.n6 x3.out.t3 371.31
R3342 x3.out.n4 x3.out.t8 371.31
R3343 x3.out.t8 x3.out.n3 371.31
R3344 x3.out.n0 x3.out.t2 227.886
R3345 x3.out.n0 x3.out.n9 25.0903
R3346 x3.out.n1 x3.out.n5 21.8335
R3347 x3.out.n3 x3.out.n1 21.6959
R3348 x3.out.n6 x3.out.n4 20.5053
R3349 x3.out.n7 x3.out.n2 19.6003
R3350 x3.out.n0 x3.out.t5 12.7763
R3351 x3.out.n9 x3.out.t0 5.5105
R3352 x3.out.n9 x3.out.t1 5.5105
R3353 x3.out.n8 x3.out.n1 5.0449
R3354 x3.out.n8 x3.out.n7 2.71826
R3355 x3.out.n7 x3.out.n6 0.90555
R3356 x3.out x3.out.n8 0.88175
R3357 x3.out x3.out.n0 0.794875
R3358 x4.out_b.n0 x4.out_b.t0 227.887
R3359 x4.out_b.n0 x4.out_b.n1 25.0905
R3360 x4.out_b.n0 x4.out_b.t3 12.777
R3361 x4.out_b.n1 x4.out_b.t1 5.5105
R3362 x4.out_b.n1 x4.out_b.t2 5.5105
R3363 x4.out_b x4.out_b.n0 0.83175
R3364 dout.n0 dout.t1 120.561
R3365 dout.n0 dout.t0 61.4115
R3366 dout dout.n0 3.88384
C0 avdd_ip inv_in 0.669037f
C1 dvss_ip xin_buf 27.955f
C2 dvdd_ip inv_m1 2.8465f
C3 x7.stby_done_b x7.clk_disable 0.724301f
C4 dvdd_ip ibias_ip 1.46921f
C5 x7.ena_done_b a_20376_n1881# 0.179696f
C6 standby_b a_19955_n2791# 0.613409f
C7 a_24530_n21674# xin 0.159429f
C8 a_19955_n2791# dvdd 0.843855f
C9 dvss_ip a_24220_n8836# 0.421193f
C10 vbp xin_buf 3.4756f
C11 vg2 vg1 1.36272f
C12 a_20121_n2241# a_20689_n2273# 0.174808f
C13 a_17913_n2241# dvdd 0.655351f
C14 a_19955_n2241# a_20471_n1869# 0.104035f
C15 a_17913_n2791# a_18828_n2791# 0.125324f
C16 a_4857_n1521# standby_ip 0.144556f
C17 a_24530_n19350# xin 0.159253f
C18 ena_ip a_21036_n1869# 0.254262f
C19 icnode a_11526_n12394# 0.136237f
C20 x3.out avss 5.85073f
C21 standby_b a_18263_n2791# 0.196932f
C22 a_18263_n2791# dvdd 0.23444f
C23 xin_buf a_10620_n9666# 0.140848f
C24 a_2130_n20844# a_2130_n21176# 0.306949f
C25 dvss_ip a_18932_n15092# 0.147461f
C26 x7.x2.Qb1 a_17747_n2791# 0.241144f
C27 vbreg xin 0.157652f
C28 x7.x2.x2.Q dvdd 0.11753f
C29 x7.x1.Qb1 a_15960_n1881# 0.171293f
C30 standby_b dvdd 6.03669f
C31 x7.clk_disable dout_filt 0.71038f
C32 a_14285_n2281# dvdd 0.170927f
C33 x7.stby_done_b a_20121_n2791# 0.953635f
C34 a_16055_n1869# dvdd 0.237126f
C35 a_17747_n2791# a_17913_n2791# 0.608363f
C36 a_15705_n2241# a_16620_n1869# 0.125324f
C37 a_16273_n2549# a_16055_n2791# 0.209641f
C38 a_2132_n15922# a_2132_n16254# 0.300147f
C39 a_17913_n2241# a_18263_n1869# 0.219472f
C40 a_16163_n2425# dvdd 0.147354f
C41 dvss_ip xin 1.63056f
C42 avdd_ip xout 7.21813f
C43 avss_ip a_2130_n21176# 0.242612f
C44 a_19003_n1943# x7.x1.x3.Q 0.119961f
C45 ena_ip x3.in_b 0.676051f
C46 standby_b a_20689_n2549# 0.183839f
C47 a_15539_n2241# a_15705_n2241# 0.608363f
C48 avss_ip vrb 6.48162f
C49 a_20689_n2549# dvdd 0.225901f
C50 dvss_ip inv_in 14.9291f
C51 dvdd_ip inv_m2 1.90217f
C52 avss_ip xin_buf 10.8147f
C53 avss_ip a_2132_n16254# 0.230757f
C54 a_19955_n2241# a_21036_n1869# 0.102355f
C55 a_24530_n22006# a_24530_n22338# 0.307023f
C56 dout_ip inv_m2 0.58891f
C57 a_18263_n1869# dvdd 0.234443f
C58 avss_ip a_2130_n18852# 0.557241f
C59 a_20689_n2273# a_20471_n1869# 0.209641f
C60 a_24220_n8504# a_24220_n8836# 0.309571f
C61 x7.stby_done_b dout_filt 0.19319f
C62 a_2971_n1521# dvdd 0.261493f
C63 standby_b a_18828_n2791# 0.25803f
C64 avss_ip a_24530_n22338# 0.488441f
C65 a_18828_n2791# dvdd 0.312702f
C66 vbp inv_in 0.265485f
C67 dvdd dout 0.550876f
C68 vn xin_buf 4.74796f
C69 avdd avss 0.110507p
C70 avss_ip a_18932_n17416# 0.56453f
C71 standby_b standby_33 0.96979f
C72 a_18932_n17084# a_18932_n17416# 0.299356f
C73 avss_ip a_24530_n20014# 0.193645f
C74 a_16620_n1869# dvdd 0.318883f
C75 a_20121_n2791# a_20471_n2791# 0.219472f
C76 dvdd_ip vg1 0.707385f
C77 a_17747_n2791# a_18263_n2791# 0.104035f
C78 a_16163_n2247# dvdd 0.146808f
C79 a_24530_n19682# a_24530_n20014# 0.307948f
C80 a_2130_n20844# xin 0.166057f
C81 dvdd_ip standby_ip 3.44007f
C82 dvss_ip a_10620_n8006# 0.203148f
C83 standby_b a_17747_n2791# 0.61356f
C84 avss_ip a_18932_n15092# 0.193668f
C85 vbreg xout 16.561699f
C86 vg2 a_2132_n17250# 0.155881f
C87 a_17913_n2241# a_18828_n1869# 0.125324f
C88 a_17747_n2791# dvdd 0.843691f
C89 standby_ip avdd 0.690112f
C90 a_19567_n2247# x7.x1.x3.Q 0.161495f
C91 x7.x2.x2.CLK a_15539_n2791# 0.240273f
C92 a_18932_n14760# a_18932_n15092# 0.299356f
C93 a_15539_n2241# dvdd 0.844577f
C94 standby_b a_21211_n2817# 0.305293f
C95 a_15539_n2241# a_16055_n1869# 0.104035f
C96 a_24530_n22006# xin 0.166657f
C97 a_21211_n2817# dvdd 0.467216f
C98 x7.x2.Qb1 a_15705_n2791# 0.756617f
C99 dvss_ip a_24220_n9168# 0.4382f
C100 dout_ip x7.ena_done_b 0.187514f
C101 a_18828_n1869# dvdd 0.312712f
C102 dvss_ip xout 14.2041f
C103 avss_ip xin 73.1079f
C104 a_17747_n2241# a_17913_n2241# 0.608363f
C105 a_19003_n2817# a_19567_n2791# 0.106826f
C106 ena_ip standby_b 3.80349f
C107 a_10620_n8670# a_10620_n9002# 0.307266f
C108 a_24530_n19682# xin 0.159253f
C109 ena_ip dvdd 7.78413f
C110 ena_ip a_16055_n1869# 0.196968f
C111 dvss_ip inv_m1 3.10099f
C112 dvdd_ip tail 3.21426f
C113 avss_ip inv_in 1.9489f
C114 a_2132_n17250# a_2132_n17582# 0.299692f
C115 x7.ena_done_b a_20121_n2241# 0.953602f
C116 dvss_ip ibias_ip 20.300303f
C117 vn xin 3.09633f
C118 a_20121_n2791# a_21036_n2791# 0.125324f
C119 dout_ip x7.clk_disable 0.150509f
C120 a_17747_n2241# dvdd 0.844319f
C121 a_16795_n1943# a_17359_n2247# 0.106826f
C122 avdd_ip avss 0.574893f
C123 a_17747_n2791# a_18828_n2791# 0.102355f
C124 xin_buf a_10620_n7674# 0.173169f
C125 standby_33 xin_buf 2.34818f
C126 a_16795_n2817# a_16620_n2791# 0.251137f
C127 a_2130_n19848# a_2130_n20180# 0.307023f
C128 a_16795_n1943# x7.x1.x2.Q 0.119961f
C129 vn inv_in 0.137437f
C130 standby_b a_14009_n2404# 0.139405f
C131 a_14009_n2404# dvdd 0.221473f
C132 a_14009_n2404# a_14285_n2281# 0.143754f
C133 ibias_ip vbp 1.36181f
C134 avdd_ip vg1 1.99589f
C135 x4.out_b avss 1.60462f
C136 ena_ip a_18263_n1869# 0.196932f
C137 avss_ip a_2130_n21508# 0.234275f
C138 inv_in dvdd 0.696511f
C139 a_2132_n14926# a_2132_n15258# 0.299356f
C140 a_15539_n2241# a_16620_n1869# 0.102355f
C141 a_21775_n2791# dvdd 0.235866f
C142 a_2971_n1521# ena_ip 0.142973f
C143 avss_ip a_2132_n16586# 0.229609f
C144 a_21211_n1943# a_21036_n1869# 0.251137f
C145 avss_ip a_2130_n19184# 0.234105f
C146 a_19955_n2241# dvdd 0.844484f
C147 a_17747_n2241# a_18263_n1869# 0.104035f
C148 standby_ip x4.out_b 0.931668f
C149 dout_ip x7.stby_done_b 0.251336f
C150 a_14009_n2701# dvdd 0.136733f
C151 ena_ip a_16620_n1869# 0.25803f
C152 avss_ip a_2132_n14262# 1.08299f
C153 a_24530_n21010# a_24530_n21342# 0.306038f
C154 a_15705_n2791# dvdd 0.631528f
C155 avss_ip a_18932_n17748# 0.633601f
C156 avss_ip xout 26.396301f
C157 x7.stby_done_b a_20376_n2791# 0.179696f
C158 avss_ip a_24530_n20346# 0.193441f
C159 x7.x2.Qb2 a_19567_n2791# 0.127083f
C160 a_2130_n21176# xin 0.159603f
C161 a_17359_n2247# x7.x1.x2.Q 0.161495f
C162 dvss_ip a_10620_n8338# 0.203056f
C163 dvss_ip inv_m2 1.69963f
C164 avss_ip a_18932_n15424# 0.222697f
C165 a_18932_n16088# a_18932_n16420# 0.299356f
C166 ena_ip a_15539_n2241# 0.611445f
C167 vbreg vg1 4.77853f
C168 vg2 a_2132_n17582# 0.155259f
C169 a_19003_n1943# a_19567_n2247# 0.106826f
C170 xin_buf xin 1.99369f
C171 ena_ip a_18828_n1869# 0.25803f
C172 dvdd_ip dout_filt 2.6369f
C173 vg2 a_2132_n15258# 0.154162f
C174 xin_buf inv_in 0.113575p
C175 x7.x1.Qb1 a_17359_n2247# 0.127083f
C176 a_24530_n22338# xin 0.168028f
C177 dout_ip dout_filt 3.64344f
C178 a_20579_n2425# dvdd 0.144018f
C179 dvss_ip a_24220_n9500# 0.412902f
C180 a_20689_n2273# dvdd 0.225909f
C181 dvss_ip vg1 6.37401f
C182 a_17747_n2241# a_18828_n1869# 0.102355f
C183 a_24530_n20014# xin 0.159204f
C184 ena_ip a_17747_n2241# 0.61356f
C185 vg2 icnode 0.421477f
C186 standby_b a_16055_n2791# 0.197065f
C187 a_2130_n21176# a_2130_n21508# 0.306949f
C188 standby_b ibias 0.299553f
C189 x3.in_b avss 1.85499f
C190 a_16055_n2791# dvdd 0.234f
C191 dvss_ip a_18932_n15756# 0.124217f
C192 a_15539_n2791# x7.x2.Qb1 0.630684f
C193 dvdd_ip vg2 0.10449f
C194 a_10620_n7674# a_10620_n8006# 0.306784f
C195 ena_ip a_14009_n2404# 0.156624f
C196 a_21211_n2817# a_21775_n2791# 0.106826f
C197 x7.x1.x4.Q dvdd 0.118427f
C198 xin_buf a_10620_n8006# 0.166951f
C199 dvss_ip x7.ena_done_b 1.48709f
C200 a_2132_n16254# a_2132_n16586# 0.299336f
C201 a_2130_n18852# a_2130_n19184# 0.307023f
C202 ena_ip a_19955_n2241# 0.613409f
C203 avss_ip a_2130_n21840# 0.234358f
C204 dvss_ip tail 0.416372f
C205 x3.out avdd 9.26841f
C206 avss_ip a_2132_n16918# 0.236584f
C207 xin_buf xout 3.51791f
C208 inv_in xin 0.302115f
C209 avss_ip a_2130_n19516# 0.234105f
C210 a_21211_n1943# dvdd 0.467188f
C211 avss_ip avss 7.31391f
C212 x7.x1.Qb2 a_19567_n2247# 0.127083f
C213 a_24220_n8836# a_24220_n9168# 0.309571f
C214 vbp tail 10.143401f
C215 avss_ip a_2132_n14594# 0.792432f
C216 standby_b a_16620_n2791# 0.25803f
C217 standby_33 ibias_ip 0.621612f
C218 a_16620_n2791# dvdd 0.320791f
C219 ibias_ip xin_buf 1.72895f
C220 standby_33 ibias 1.10533f
C221 x7.ena_done_b a_15000_n1881# 0.263497f
C222 avss_ip vg1 20.7774f
C223 a_18932_n17416# a_18932_n17748# 0.299356f
C224 x7.ena_done_b a_15705_n2241# 0.195776f
C225 avss_ip a_24530_n20678# 0.193645f
C226 a_24530_n20014# a_24530_n20346# 0.307948f
C227 a_2130_n21508# xin 0.167748f
C228 dvss_ip a_10620_n8670# 0.203056f
C229 standby_b avss 1.88627f
C230 avss_ip a_18932_n15756# 0.237057f
C231 dvdd avss 0.230567f
C232 avdd_ip vg2 0.488655f
C233 standby_b a_15539_n2791# 0.61161f
C234 vg2 a_2132_n17914# 0.154785f
C235 a_15539_n2791# dvdd 0.651082f
C236 a_17913_n2791# a_18481_n2549# 0.174808f
C237 dvss_ip x7.stby_done_b 1.50194f
C238 icnode avdd 0.342783f
C239 a_2130_n19184# xin 0.164971f
C240 ena_ip a_20689_n2273# 0.183839f
C241 x7.x1.Qb2 a_18168_n1881# 0.171293f
C242 dvdd_ip dout_ip 1.84294f
C243 a_18932_n15092# a_18932_n15424# 0.299356f
C244 vg2 a_2132_n15590# 0.156683f
C245 a_15000_n1881# x7.x1.x2.CLK 0.134958f
C246 dvss_ip a_24220_n9832# 0.676369f
C247 standby_ip standby_b 1.50129f
C248 x7.x2.Qb1 a_15960_n2791# 0.171293f
C249 standby_ip dvdd 10.280701f
C250 x7.ena_done_b a_17913_n2241# 0.193771f
C251 a_21775_n2247# dvdd 0.236037f
C252 vg1 a_22601_n15524# 0.440171f
C253 ena_ip ibias 0.171255f
C254 a_19003_n2817# x7.x2.x3.Q 0.119961f
C255 xin xout 12.4168f
C256 a_15705_n2241# a_16273_n2273# 0.174808f
C257 a_24530_n20346# xin 0.158905f
C258 a_10620_n9002# a_10620_n9334# 0.307266f
C259 x7.stby_done_b x7.x2.Qb1 0.111333f
C260 x7.stby_done_b a_15000_n2791# 0.263439f
C261 inv_in xout 1.1656f
C262 x7.stby_done_b a_17913_n2791# 0.193805f
C263 a_2132_n17582# a_2132_n17914# 0.299336f
C264 x7.ena_done_b dvdd 6.16668f
C265 dvss_ip dout_filt 7.440259f
C266 xin_buf a_10620_n8338# 0.166314f
C267 vn tail 0.670061f
C268 inv_in inv_m1 0.243271f
C269 vg2 a_18932_n14428# 0.5683f
C270 a_2130_n20180# a_2130_n20512# 0.308883f
C271 vg2 vbreg 4.29131f
C272 avss_ip a_3134_n13324# 1.13338f
C273 standby_33 avss 1.55853f
C274 a_18481_n2549# a_18263_n2791# 0.209641f
C275 ena_ip a_21211_n1943# 0.305293f
C276 x7.clk_disable dvdd 0.383458f
C277 icnode a_8268_n12482# 1.47989f
C278 x7.x1.x3.Q dvdd 0.112744f
C279 avss_ip a_2130_n22172# 0.237164f
C280 standby_b a_18481_n2549# 0.183839f
C281 a_2132_n15258# a_2132_n15590# 0.29969f
C282 a_4857_n1521# standby 0.18913f
C283 a_18481_n2549# dvdd 0.225643f
C284 vrb vg1 0.454276f
C285 x7.x2.x4.Q dvdd 0.118417f
C286 avdd_ip icnode 43.6422f
C287 dvss_ip vg2 3.9276f
C288 x7.x1.x2.CLK dvdd 0.406962f
C289 avss_ip a_2132_n17250# 0.236693f
C290 x7.stby_done_b a_19955_n2791# 0.648907f
C291 avss_ip a_2130_n19848# 0.234105f
C292 dvdd_ip avdd_ip 3.59467f
C293 a_16273_n2273# dvdd 0.230873f
C294 a_19955_n2791# a_20121_n2791# 0.608363f
C295 a_19567_n2791# x7.x2.x3.Q 0.161495f
C296 a_16273_n2273# a_16055_n1869# 0.209641f
C297 a_15705_n2791# a_16055_n2791# 0.219472f
C298 avdd_ip avdd 9.33419f
C299 avss_ip a_2132_n14926# 0.652798f
C300 a_24530_n21342# a_24530_n21674# 0.307869f
C301 a_17913_n2241# a_18481_n2273# 0.174808f
C302 a_24220_n7840# a_24220_n8172# 0.307266f
C303 ena_ip avss 1.87755f
C304 avss_ip a_24530_n21010# 0.193969f
C305 standby_b x7.stby_done_b 0.752988f
C306 a_2130_n21840# xin 0.172286f
C307 x4.out_b avdd 7.47205f
C308 x7.stby_done_b dvdd 5.41509f
C309 a_20121_n2791# dvdd 0.653362f
C310 dvss_ip a_10620_n9002# 0.19184f
C311 avss_ip a_18932_n16088# 0.544237f
C312 a_18932_n16420# a_18932_n16752# 0.299356f
C313 a_18481_n2273# dvdd 0.225651f
C314 a_20121_n2241# a_20471_n1869# 0.219472f
C315 a_24530_n19018# a_24530_n19350# 0.307948f
C316 a_2130_n19516# xin 0.164971f
C317 ena_ip standby_ip 4.63202f
C318 xin_buf tail 4.40803f
C319 standby_b a_19003_n2817# 0.357273f
C320 a_19003_n2817# dvdd 0.456345f
C321 vg2 a_2132_n15922# 0.154604f
C322 x3.in_b x3.out 0.933643f
C323 dvdd_ip vbreg 0.819111f
C324 inv_in avss 0.144174f
C325 a_20121_n2791# a_20689_n2549# 0.174808f
C326 a_16795_n1943# dvdd 0.461387f
C327 a_19955_n2791# a_20471_n2791# 0.104035f
C328 vg1 xin 0.215332p
C329 x7.x2.Qb2 a_17913_n2791# 0.756617f
C330 ibias_ip ibias 0.846688f
C331 a_24530_n20678# xin 0.159253f
C332 a_15705_n2791# a_16620_n2791# 0.125324f
C333 ena_ip x7.ena_done_b 0.702741f
C334 dvss_ip a_24220_n7840# 0.402598f
C335 avss_ip vg2 0.156017p
C336 a_2130_n21508# a_2130_n21840# 0.307948f
C337 dout_filt dvdd 1.76335f
C338 a_18481_n2273# a_18263_n1869# 0.209641f
C339 dvdd_ip dvss_ip 0.502455p
C340 a_10620_n8006# a_10620_n8338# 0.307266f
C341 x7.x1.x2.CLK a_15539_n2241# 0.240273f
C342 a_21211_n2817# x7.x2.x4.Q 0.119961f
C343 dvss_ip dout_ip 6.78359f
C344 xin_buf a_10620_n8670# 0.16582f
C345 standby_b a_20471_n2791# 0.196932f
C346 x7.x1.Qb1 a_15705_n2241# 0.756617f
C347 a_15539_n2791# a_15705_n2791# 0.608363f
C348 a_20471_n2791# dvdd 0.234572f
C349 a_2132_n16586# a_2132_n16918# 0.298902f
C350 a_14009_n2404# x7.ena_done_b 0.173521f
C351 a_19003_n1943# dvdd 0.456365f
C352 a_20121_n2241# a_21036_n1869# 0.125324f
C353 avss_ip x3.out 2.42141f
C354 dvdd_ip vbp 26.197498f
C355 a_19003_n2817# a_18828_n2791# 0.251137f
C356 a_2130_n19184# a_2130_n19516# 0.308883f
C357 x7.x2.Qb2 a_19955_n2791# 0.241144f
C358 a_4857_n1521# dvdd 0.264852f
C359 ena_ip a_16273_n2273# 0.183844f
C360 a_19567_n2791# dvdd 0.230807f
C361 tail xin 1.6128f
C362 avss_ip a_2132_n17582# 0.229847f
C363 x3.in_b avdd 1.00629f
C364 x7.ena_done_b a_19955_n2241# 0.648846f
C365 avss_ip a_2130_n20180# 0.234105f
C366 a_19955_n2791# a_21036_n2791# 0.102355f
C367 a_20689_n2549# a_20471_n2791# 0.209641f
C368 a_14009_n2404# x7.clk_disable 0.122842f
C369 dout_ip a_15000_n2791# 0.148426f
C370 a_17359_n2247# dvdd 0.234839f
C371 a_16795_n1943# a_16620_n1869# 0.251137f
C372 a_2132_n14262# a_2132_n14594# 0.299692f
C373 inv_m1 inv_m2 0.947856f
C374 inv_in tail 0.604094f
C375 a_21211_n1943# x7.x1.x4.Q 0.119961f
C376 x7.x1.x2.Q dvdd 0.116301f
C377 a_24220_n9168# a_24220_n9500# 0.30635f
C378 dout_filt dout 0.639323f
C379 standby_b x7.x2.Qb2 0.347451f
C380 avss_ip a_2132_n15258# 0.245921f
C381 dout_ip a_15000_n1881# 0.142224f
C382 avdd_ip vbreg 39.105396f
C383 x7.x2.Qb2 dvdd 1.2179f
C384 a_18932_n17748# vg1 0.408298f
C385 vg1 xout 0.637062f
C386 ena_ip a_18481_n2273# 0.183839f
C387 avss_ip a_24530_n21342# 0.187124f
C388 a_21775_n2791# x7.x2.x4.Q 0.161495f
C389 x7.x1.Qb1 dvdd 1.22948f
C390 standby_b a_21036_n2791# 0.254262f
C391 a_24530_n20346# a_24530_n20678# 0.307948f
C392 a_2130_n22172# xin 0.581116f
C393 avss_ip icnode 33.2949f
C394 a_15539_n2791# a_16055_n2791# 0.104035f
C395 a_21036_n2791# dvdd 0.31454f
C396 dvss_ip a_10620_n9334# 0.174627f
C397 x7.clk_disable a_14009_n2701# 0.419961f
C398 a_15000_n2791# x7.x2.x2.CLK 0.134958f
C399 avss_ip a_18932_n16420# 0.690377f
C400 a_18932_n15424# vg1 0.560332f
C401 a_19567_n2247# dvdd 0.230816f
C402 avss_ip a_24530_n19018# 0.187516f
C403 dvdd_ip avss_ip 2.2865f
C404 avdd_ip dvss_ip 20.735699f
C405 x7.x1.Qb2 a_17913_n2241# 0.756617f
C406 a_2130_n19848# xin 0.165429f
C407 a_14009_n2404# x7.stby_done_b 0.245503f
C408 avss_ip avdd 2.34938f
C409 vg2 vrb 4.64006f
C410 ena_ip a_16795_n1943# 0.357273f
C411 a_18932_n15424# a_18932_n15756# 0.299356f
C412 a_18371_n2425# dvdd 0.143768f
C413 vg2 a_2132_n16254# 0.155116f
C414 xin_buf vg2 3.5685f
C415 standby_ip ibias 0.288163f
C416 dvdd ena 0.377442f
C417 dvdd_ip vn 1.05192f
C418 x7.stby_done_b a_21775_n2791# 0.160191f
C419 x7.x1.Qb2 dvdd 1.22125f
C420 a_21775_n2247# x7.x1.x4.Q 0.161495f
C421 a_16795_n2817# a_17359_n2791# 0.106826f
C422 a_10620_n9334# a_10620_n9666# 0.310516f
C423 a_24530_n21010# xin 0.159641f
C424 dvss_ip a_24220_n8172# 0.412162f
C425 tail xout 1.23159f
C426 dvdd_ip dvdd 14.0307f
C427 standby_b dout_ip 0.325806f
C428 a_19003_n1943# a_18828_n1869# 0.251137f
C429 dout_ip dvdd 1.38045f
C430 dvss_ip a_18932_n16752# 0.11359f
C431 standby_b avdd 0.807362f
C432 avdd dvdd 0.106948f
C433 x7.stby_done_b a_15705_n2791# 0.20129f
C434 ena_ip a_19003_n1943# 0.357273f
C435 xin_buf a_10620_n9002# 0.156922f
C436 a_2130_n20512# a_2130_n20844# 0.307948f
C437 a_17747_n2791# x7.x2.Qb2 0.630684f
C438 dvss_ip a_18932_n14428# 0.117297f
C439 dvss_ip vbreg 7.841839f
C440 a_15539_n2791# a_16620_n2791# 0.102355f
C441 a_21211_n1943# a_21775_n2247# 0.106826f
C442 a_20121_n2241# dvdd 0.655086f
C443 a_2971_n1521# ena 0.188898f
C444 x7.x2.x2.CLK dvdd 0.367738f
C445 a_2132_n15590# a_2132_n15922# 0.298886f
C446 standby_b a_16273_n2549# 0.183867f
C447 avss_ip a_8268_n12482# 3.56481f
C448 a_16273_n2549# dvdd 0.232251f
C449 a_15539_n2241# x7.x1.Qb1 0.630684f
C450 vg2 xin 6.28706f
C451 avdd_ip avss_ip 0.856941p
C452 avss_ip a_2132_n17914# 0.528436f
C453 avss_ip a_2130_n20512# 0.234105f
C454 a_14009_n2701# dout_filt 0.140187f
C455 a_21211_n2817# a_21036_n2791# 0.251137f
C456 dvdd_ip dout 1.66314f
C457 x7.x2.Qb2 a_18168_n2791# 0.171293f
C458 a_20579_n2247# dvdd 0.144024f
C459 xin_buf icnode 3.62534f
C460 inv_in vg2 0.137694f
C461 standby_ip avss 1.86774f
C462 dvdd_ip a_10620_n7674# 0.100908f
C463 avss_ip a_2132_n15590# 0.241841f
C464 dvdd_ip standby_33 3.26892f
C465 ena_ip x7.x1.Qb1 0.347396f
C466 dvdd_ip vrb 0.182588f
C467 a_24530_n21674# a_24530_n22006# 0.306949f
C468 dvdd_ip xin_buf 19.1703f
C469 dvss_ip vbp 1.28877f
C470 standby_33 avdd 9.00234f
C471 a_24220_n8172# a_24220_n8504# 0.310516f
C472 dout_ip xin_buf 0.1539f
C473 avss_ip a_24530_n21674# 0.194498f
C474 xin_buf avdd 0.176178f
C475 x7.x1.Qb1 a_17747_n2241# 0.241144f
C476 dvss_ip a_10620_n9666# 0.193818f
C477 x7.x2.Qb1 a_17359_n2791# 0.127083f
C478 avss_ip a_18932_n16752# 0.452744f
C479 a_18932_n16752# a_18932_n17084# 0.299356f
C480 a_18932_n15756# vg1 0.267005f
C481 avss_ip a_24530_n19350# 0.193645f
C482 a_20471_n1869# dvdd 0.234574f
C483 a_24530_n19350# a_24530_n19682# 0.307948f
C484 a_2130_n20180# xin 0.1652f
C485 ena_ip x7.x1.Qb2 0.347451f
C486 a_16795_n2817# x7.x2.x2.Q 0.119961f
C487 avss_ip a_18932_n14428# 0.151712f
C488 standby_b a_16795_n2817# 0.357273f
C489 avss_ip vbreg 13.769401f
C490 vg2 a_2132_n16586# 0.154861f
C491 a_16795_n2817# dvdd 0.462729f
C492 standby_ip x7.ena_done_b 0.121215f
C493 x7.ena_done_b a_21775_n2247# 0.160065f
C494 ena_ip dout_ip 0.203453f
C495 a_18932_n14428# a_18932_n14760# 0.299356f
C496 a_17747_n2241# x7.x1.Qb2 0.630684f
C497 ena_ip avdd 0.711014f
C498 a_24530_n21342# xin 0.166712f
C499 dvss_ip a_24220_n8504# 0.435581f
C500 vg2 xout 0.938912f
C501 dvss_ip avss_ip 23.869501f
C502 a_2130_n21840# a_2130_n22172# 0.306949f
C503 a_10620_n8338# a_10620_n8670# 0.307266f
C504 a_24530_n19018# xin 0.126575f
C505 dvdd_ip xin 4.32555f
C506 inv_in a_24220_n7840# 0.423473f
C507 inv_in icnode 0.110238f
C508 xin_buf a_8268_n12482# 0.261082f
C509 xin_buf a_10620_n9334# 0.138691f
C510 dvss_ip a_18932_n14760# 0.144339f
C511 vbreg a_22601_n15524# 2.38713f
C512 dvss_ip vn 6.6789f
C513 avdd_ip xin_buf 9.05887f
C514 dvdd_ip inv_in 10.408401f
C515 a_2132_n16918# a_2132_n17250# 0.299677f
C516 a_21036_n1869# dvdd 0.31455f
C517 x7.x1.Qb2 a_19955_n2241# 0.241144f
C518 dvdd standby 0.386478f
C519 a_2130_n19516# a_2130_n19848# 0.307948f
C520 dvss_ip standby_b 3.55257f
C521 dvss_ip dvdd 20.2555f
C522 a_17359_n2791# x7.x2.x2.Q 0.161495f
C523 standby_33 x4.out_b 0.696369f
C524 x7.x2.x3.Q dvdd 0.112734f
C525 a_17359_n2791# dvdd 0.236098f
C526 dvss_ip a_22601_n15524# 0.147611f
C527 avss_ip a_2130_n20844# 0.234274f
C528 a_2132_n14594# a_2132_n14926# 0.298902f
C529 a_24220_n9500# a_24220_n9832# 0.307266f
C530 avss_ip a_2132_n15922# 0.231212f
C531 standby_b x7.x2.Qb1 0.347492f
C532 a_19955_n2241# a_20121_n2241# 0.608363f
C533 x7.x2.Qb1 dvdd 1.15446f
C534 x3.in_b dvdd 0.22553f
C535 a_17913_n2791# a_18263_n2791# 0.219472f
C536 vbreg vrb 0.239025f
C537 a_15000_n2791# dvdd 0.238886f
C538 ena_ip a_20471_n1869# 0.196932f
C539 a_18371_n2247# dvdd 0.143775f
C540 avss_ip a_24530_n22006# 0.186833f
C541 a_17913_n2791# dvdd 0.653627f
C542 x7.ena_done_b x7.stby_done_b 1.61077f
C543 a_24530_n20678# a_24530_n21010# 0.307948f
C544 a_15000_n1881# dvdd 0.25026f
C545 avss_ip a_18932_n17084# 0.726269f
C546 a_14285_n2079# dvdd 0.149051f
C547 avss_ip a_24530_n19682# 0.193645f
C548 a_24530_n19018# xout 0.377144f
C549 a_15705_n2241# dvdd 0.668389f
C550 dvdd_ip xout 4.80514f
C551 avdd_ip xin 6.74409f
C552 dvss_ip dout 6.66227f
C553 a_15705_n2241# a_16055_n1869# 0.219472f
C554 a_2130_n20512# xin 0.164971f
C555 a_15705_n2791# a_16273_n2549# 0.174808f
C556 dvss_ip a_10620_n7674# 0.359271f
C557 dvss_ip standby_33 3.27772f
C558 avss_ip a_18932_n14760# 0.178926f
C559 a_18932_n15756# a_18932_n16088# 0.299356f
C560 dvss_ip vrb 1.20334f
C561 vg2 a_2132_n16918# 0.156129f
C562 xout dvss 4.260475f
C563 xin dvss 11.878201f
C564 dout dvss 6.13496f
C565 standby dvss 1.31628f
C566 ena dvss 1.29685f
C567 avss dvss 11.55251f
C568 ibias dvss 6.38685f
C569 dvdd dvss 0.140297p
C570 avdd dvss 95.102425f
C571 a_24530_n22338# dvss 0.197063f
C572 a_2130_n22172# dvss 0.199586f
C573 a_24530_n22006# dvss 0.197123f
C574 a_2130_n21840# dvss 0.205689f
C575 a_24530_n21674# dvss 0.191047f
C576 a_2130_n21508# dvss 0.205669f
C577 a_24530_n21342# dvss 0.197488f
C578 a_2130_n21176# dvss 0.199691f
C579 a_24530_n21010# dvss 0.191047f
C580 a_2130_n20844# dvss 0.20567f
C581 a_24530_n20678# dvss 0.191047f
C582 a_2130_n20512# dvss 0.205512f
C583 a_24530_n20346# dvss 0.190888f
C584 a_2130_n20180# dvss 0.205515f
C585 a_24530_n20014# dvss 0.190952f
C586 a_2130_n19848# dvss 0.205518f
C587 a_24530_n19682# dvss 0.191047f
C588 a_2130_n19516# dvss 0.205512f
C589 a_24530_n19350# dvss 0.191047f
C590 a_2130_n19184# dvss 0.205515f
C591 a_24530_n19018# dvss 0.191047f
C592 a_2130_n18852# dvss 0.205518f
C593 vg1 dvss -0.243245f
C594 a_2132_n17914# dvss 0.204459f
C595 a_18932_n17748# dvss 0.183093f
C596 a_2132_n17582# dvss 0.204591f
C597 a_18932_n17416# dvss 0.183093f
C598 a_2132_n17250# dvss 0.199339f
C599 a_18932_n17084# dvss 0.183093f
C600 a_2132_n16918# dvss 0.199339f
C601 a_18932_n16752# dvss 0.183093f
C602 a_2132_n16586# dvss 0.204459f
C603 a_18932_n16420# dvss 0.183093f
C604 a_2132_n16254# dvss 0.204591f
C605 a_18932_n16088# dvss 0.183093f
C606 a_2132_n15922# dvss 0.204459f
C607 a_18932_n15756# dvss 0.182956f
C608 a_2132_n15590# dvss 0.199472f
C609 a_18932_n15424# dvss 0.182179f
C610 a_2132_n15258# dvss 0.204459f
C611 a_18932_n15092# dvss 0.207654f
C612 a_2132_n14926# dvss 0.204459f
C613 a_18932_n14760# dvss 0.204459f
C614 a_2132_n14594# dvss 0.205118f
C615 a_18932_n14428# dvss 0.179624f
C616 a_2132_n14262# dvss 0.204591f
C617 vrb dvss 0.16284f
C618 a_3134_n13324# dvss 0.190586f
C619 vbreg dvss 4.41296f
C620 a_8268_n12482# dvss 1.07843f
C621 icnode dvss 6.39639f
C622 vg2 dvss 4.397135f
C623 a_24220_n9832# dvss 0.206087f
C624 a_10620_n9666# dvss 0.186956f
C625 a_24220_n9500# dvss 0.206087f
C626 a_10620_n9334# dvss 0.205627f
C627 a_24220_n9168# dvss 0.187048f
C628 a_10620_n9002# dvss 0.205994f
C629 a_24220_n8836# dvss 0.186681f
C630 a_10620_n8670# dvss 0.205994f
C631 a_24220_n8504# dvss 0.186681f
C632 a_10620_n8338# dvss 0.205994f
C633 a_24220_n8172# dvss 0.20572f
C634 a_10620_n8006# dvss 0.205994f
C635 a_24220_n7840# dvss 0.206087f
C636 a_10620_n7674# dvss 0.200388f
C637 tail dvss 0.375177f
C638 inv_m2 dvss 0.562228f
C639 inv_m1 dvss 0.704134f
C640 inv_in dvss 6.596221f
C641 xin_buf dvss 7.43464f
C642 vn dvss 1.05209f
C643 vbp dvss 3.48575f
C644 x4.out_b dvss 1.061455f
C645 x3.out dvss 2.07027f
C646 a_21775_n2791# dvss 0.2255f
C647 a_21036_n2791# dvss 0.266719f
C648 a_21211_n2817# dvss 0.721269f
C649 a_20471_n2791# dvss 0.269124f
C650 a_20689_n2549# dvss 0.185767f
C651 a_20121_n2791# dvss 0.307225f
C652 a_19955_n2791# dvss 0.565683f
C653 a_19567_n2791# dvss 0.198301f
C654 a_18828_n2791# dvss 0.263274f
C655 a_19003_n2817# dvss 0.699257f
C656 a_18263_n2791# dvss 0.269103f
C657 a_18481_n2549# dvss 0.18572f
C658 a_17913_n2791# dvss 0.307195f
C659 x7.x2.Qb2 dvss 0.510929f
C660 a_17747_n2791# dvss 0.56557f
C661 dout_filt dvss 5.8975f
C662 a_17359_n2791# dvss 0.198798f
C663 a_16620_n2791# dvss 0.264546f
C664 a_16795_n2817# dvss 0.700156f
C665 a_16055_n2791# dvss 0.276301f
C666 a_16273_n2549# dvss 0.187951f
C667 a_15705_n2791# dvss 0.351701f
C668 x7.x2.Qb1 dvss 0.540099f
C669 a_15539_n2791# dvss 0.620802f
C670 x7.x2.x2.CLK dvss 0.389657f
C671 a_14009_n2701# dvss 0.233987f
C672 x7.clk_disable dvss 4.60726f
C673 a_15000_n2791# dvss 0.342356f
C674 x7.stby_done_b dvss 2.67735f
C675 ibias_ip dvss 4.3844f
C676 standby_33 dvss 5.81519f
C677 a_21775_n2247# dvss 0.225515f
C678 a_21036_n1869# dvss 0.266723f
C679 a_21211_n1943# dvss 0.721243f
C680 a_20471_n1869# dvss 0.269077f
C681 a_20689_n2273# dvss 0.185771f
C682 a_20121_n2241# dvss 0.307238f
C683 a_19955_n2241# dvss 0.56568f
C684 a_19567_n2247# dvss 0.198316f
C685 a_18828_n1869# dvss 0.263277f
C686 a_19003_n1943# dvss 0.699232f
C687 a_18263_n1869# dvss 0.269056f
C688 a_18481_n2273# dvss 0.185724f
C689 a_17913_n2241# dvss 0.307208f
C690 x7.x1.Qb2 dvss 0.510897f
C691 a_17747_n2241# dvss 0.565567f
C692 a_17359_n2247# dvss 0.198813f
C693 a_16620_n1869# dvss 0.264549f
C694 a_16795_n1943# dvss 0.70013f
C695 a_16055_n1869# dvss 0.271684f
C696 a_16273_n2273# dvss 0.187955f
C697 a_15705_n2241# dvss 0.341334f
C698 x7.x1.Qb1 dvss 0.528095f
C699 a_15539_n2241# dvss 0.580494f
C700 x7.x1.x2.CLK dvss 0.38222f
C701 a_15000_n1881# dvss 0.351108f
C702 x7.ena_done_b dvss 2.38862f
C703 dout_ip dvss 6.69846f
C704 a_14009_n2404# dvss 0.605583f
C705 standby_b dvss 25.5709f
C706 x3.in_b dvss 1.85375f
C707 standby_ip dvss 20.4485f
C708 ena_ip dvss 14.4202f
C709 a_4857_n1521# dvss 0.293752f
C710 a_2971_n1521# dvss 0.292633f
C711 avss_ip dvss 27.73396f
C712 dvss_ip dvss 41.9846f
C713 avdd_ip dvss 0.98484p
C714 dvdd_ip dvss 0.352295p
C715 dout.t0 dvss 0.223213f
C716 dout.n0 dvss 3.29562f
C717 x4.out_b.n0 dvss 5.53652f
C718 x4.out_b.t3 dvss 1.30743f
C719 x4.out_b.n1 dvss 0.140668f
C720 x3.out.n0 dvss 7.39524f
C721 x3.out.n1 dvss 0.893601f
C722 x3.out.n2 dvss 0.392503f
C723 x3.out.t6 dvss 0.479128f
C724 x3.out.n3 dvss 0.382459f
C725 x3.out.t8 dvss 0.458669f
C726 x3.out.n4 dvss 0.394877f
C727 x3.out.t7 dvss 0.479113f
C728 x3.out.t4 dvss 0.458669f
C729 x3.out.n5 dvss 0.382543f
C730 x3.out.t3 dvss 0.458669f
C731 x3.out.n6 dvss 0.161457f
C732 x3.out.n7 dvss 0.521199f
C733 x3.out.n8 dvss 1.69978f
C734 x3.out.t5 dvss 1.7568f
C735 x3.out.n9 dvss 0.188953f
C736 vrb.t2 dvss 0.274519f
C737 vrb.t4 dvss 0.33602f
C738 vrb.n0 dvss 3.02505f
C739 vrb.t3 dvss 0.274548f
C740 vrb.t1 dvss 0.333171f
C741 vrb.n1 dvss 3.02989f
C742 vrb.n2 dvss 2.40037f
C743 vrb.n3 dvss 1.30448f
C744 vg2.n0 dvss 0.282949f
C745 vg2.n1 dvss 0.261019f
C746 vg2.t9 dvss 0.640509f
C747 vg2.n2 dvss 1.17147f
C748 vg2.n3 dvss 0.244906f
C749 vg2.n4 dvss 0.522037f
C750 vg2.t6 dvss 0.628646f
C751 vg2.n5 dvss 0.314177f
C752 vg2.n6 dvss 0.32051f
C753 vg2.n7 dvss 0.282949f
C754 vg2.n8 dvss 0.261019f
C755 vg2.t5 dvss 0.640544f
C756 vg2.n9 dvss 1.17258f
C757 vg2.n10 dvss 0.244906f
C758 vg2.n11 dvss 0.522037f
C759 vg2.t7 dvss 0.628646f
C760 vg2.n12 dvss 0.313029f
C761 vg2.n13 dvss 0.32051f
C762 vg2.t8 dvss 0.505469f
C763 vg2.t2 dvss 39.125f
C764 vg2.t1 dvss 39.3426f
C765 vg2.t4 dvss 39.3426f
C766 vg2.t3 dvss 39.11f
C767 vg2.n15 dvss 9.00528f
C768 vg2.n16 dvss 2.91513f
C769 xin.n0 dvss 0.172822f
C770 xin.n5 dvss 0.184148f
C771 xin.t18 dvss 0.1922f
C772 xin.t15 dvss 0.19211f
C773 xin.n6 dvss 0.184148f
C774 xin.t13 dvss 0.19211f
C775 xin.t19 dvss 0.19211f
C776 xin.t16 dvss 0.19211f
C777 xin.t11 dvss 0.19211f
C778 xin.t10 dvss 0.19211f
C779 xin.t17 dvss 0.19211f
C780 xin.t14 dvss 0.19211f
C781 xin.t12 dvss 0.19211f
C782 xin.t9 dvss 0.19211f
C783 xin.t6 dvss 0.19211f
C784 xin.n21 dvss 0.175223f
C785 xin.n22 dvss 0.784969f
C786 xin.n23 dvss 0.308623f
C787 xin.n24 dvss 0.374761f
C788 xin.t20 dvss 0.828066f
C789 xin.t7 dvss 0.79628f
C790 xin.n25 dvss 0.514f
C791 xin.n26 dvss 0.386948f
C792 xin.n27 dvss 3.79487f
C793 xin.n28 dvss 4.5191f
C794 xin.n29 dvss 3.61279f
C795 xin.t2 dvss 57.0239f
C796 xin.t4 dvss 44.1862f
C797 xin.t1 dvss 44.012f
C798 xin.t0 dvss 0.124226f
C799 xin.n30 dvss 4.7746f
C800 xin.n31 dvss 27.2736f
C801 xin.t5 dvss 31.1925f
C802 xin.n32 dvss 27.266699f
C803 xin.t3 dvss 31.1614f
C804 xin.n33 dvss 27.270199f
C805 xin.n34 dvss 3.77704f
C806 xin.n35 dvss 1.85671f
C807 xin.n36 dvss 0.500575f
C808 vg1.n0 dvss 0.44953f
C809 vg1.t8 dvss 46.057503f
C810 vg1.t9 dvss 46.8352f
C811 vg1.t4 dvss 23.996801f
C812 vg1.n1 dvss 23.9575f
C813 vg1.t7 dvss 23.996801f
C814 vg1.n2 dvss 23.4861f
C815 vg1.t6 dvss 23.996801f
C816 vg1.n3 dvss 12.9859f
C817 vg1.n4 dvss 15.228601f
C818 vg1.n5 dvss 3.04049f
C819 vg1.n6 dvss 1.50262f
C820 vg1.t2 dvss 0.271659f
C821 vg1.t5 dvss 0.353472f
C822 vg1.n7 dvss 0.229145f
C823 vg1.n9 dvss 0.281876f
C824 vg1.n10 dvss 0.146945f
C825 vg1.n11 dvss 0.153437f
C826 vg1.n12 dvss 0.372304f
C827 x3.out_b.t6 dvss 0.402581f
C828 x3.out_b.n0 dvss 0.790285f
C829 x3.out_b.n1 dvss 1.5584f
C830 x3.out_b.n2 dvss 6.60541f
C831 x3.out_b.t4 dvss 0.420289f
C832 x3.out_b.n3 dvss 0.339622f
C833 x3.out_b.t7 dvss 0.402581f
C834 x3.out_b.n4 dvss 0.342378f
C835 x3.out_b.t8 dvss 0.420331f
C836 x3.out_b.n5 dvss 0.338349f
C837 x3.out_b.t3 dvss 0.402581f
C838 x3.out_b.n6 dvss 0.345348f
C839 x3.out_b.n7 dvss 0.58218f
C840 x3.out_b.t5 dvss 1.5189f
C841 x3.out_b.n8 dvss 0.163419f
C842 avdd.n0 dvss 0.492818f
C843 avdd.n1 dvss 1.6981f
C844 avdd.n4 dvss 0.266474f
C845 avdd.n5 dvss 0.585389f
C846 avdd.n6 dvss 1.03476f
C847 avdd.n7 dvss 1.03476f
C848 avdd.t13 dvss 0.894926f
C849 avdd.t2 dvss 0.702496f
C850 avdd.t11 dvss 0.894926f
C851 avdd.t8 dvss 0.702496f
C852 avdd.n8 dvss 0.46232f
C853 avdd.t17 dvss 7.53658f
C854 avdd.n9 dvss 7.5153f
C855 avdd.t16 dvss 9.12027f
C856 avdd.t19 dvss 7.25381f
C857 avdd.n10 dvss 7.71793f
C858 avdd.t18 dvss 9.163919f
C859 avdd.n11 dvss 3.68652f
C860 avdd.n12 dvss 0.768588f
C861 avdd.n13 dvss 0.579746f
C862 avdd.n14 dvss 0.560241f
C863 avdd.n15 dvss 0.353066f
C864 avdd.n16 dvss 0.487874f
C865 avdd.n17 dvss 3.7478f
C866 avdd.n18 dvss 0.731215f
C867 avdd.n21 dvss 1.93441f
C868 avdd.n22 dvss 0.967373f
C869 avdd.t14 dvss 0.135207f
C870 avdd.n23 dvss 0.34342f
C871 avdd.n24 dvss 5.68989f
C872 avdd.n25 dvss 1.05169f
C873 avdd.n26 dvss 1.1887f
C874 avdd.n27 dvss 1.1887f
C875 avdd.n28 dvss 4.46094f
C876 avdd.n29 dvss 1.35368f
C877 avdd.n32 dvss 0.548551f
C878 avdd.n33 dvss 1.56238f
C879 avdd.n34 dvss 1.46595f
C880 avdd.n35 dvss 0.107384f
C881 avdd.n36 dvss 0.107943f
C882 avdd.n37 dvss 0.158157f
C883 avdd.t4 dvss 2.51038f
C884 avdd.n39 dvss 0.10415f
C885 avdd.n40 dvss 0.107943f
C886 avdd.n41 dvss 0.559667f
C887 avdd.n43 dvss 0.687088f
C888 avdd.n44 dvss 1.48367f
C889 avdd.n45 dvss 1.13727f
C890 avdd.n46 dvss 0.744579f
C891 avdd.n47 dvss 2.46523f
C892 avdd.n48 dvss 3.43088f
C893 avdd.n49 dvss 1.15288f
C894 avdd.n50 dvss 0.362301f
C895 avdd.n51 dvss 0.321745f
C896 avdd.n52 dvss 0.106191f
C897 avdd.n53 dvss 1.67879f
C898 avdd.n54 dvss 0.106191f
C899 avdd.n55 dvss 0.158157f
C900 avdd.n58 dvss 0.106191f
C901 avdd.n59 dvss 1.67879f
C902 avdd.n60 dvss 0.106191f
C903 avdd.n62 dvss 0.116928f
C904 avdd.n63 dvss 0.719248f
C905 avdd.n64 dvss 1.37927f
C906 avdd.n65 dvss 1.47231f
C907 avdd.n66 dvss 1.45902f
C908 avdd.n67 dvss 0.366507f
C909 avdd.n68 dvss 0.107943f
C910 avdd.n69 dvss 0.158157f
C911 avdd.t6 dvss 2.51038f
C912 avdd.n70 dvss 0.10415f
C913 avdd.n71 dvss 0.107943f
C914 avdd.n72 dvss 0.107384f
C915 avdd.n74 dvss 0.106191f
C916 avdd.n75 dvss 1.67879f
C917 avdd.n76 dvss 0.106191f
C918 avdd.n77 dvss 0.158157f
C919 avdd.n78 dvss 0.106191f
C920 avdd.n79 dvss 1.67879f
C921 avdd.n80 dvss 0.106191f
C922 avdd.n81 dvss 0.319178f
C923 avdd.n82 dvss 0.73302f
C924 avdd.n83 dvss 1.95073f
C925 avdd.n84 dvss 4.13419f
C926 avdd.n85 dvss 0.707422f
C927 avdd.n86 dvss 0.479606f
C928 avdd.n87 dvss 1.32047f
C929 avdd.n88 dvss 1.35617f
C930 avdd.n89 dvss 0.536684f
C931 avdd.n90 dvss 1.19042f
C932 avdd.n91 dvss 4.48227f
C933 avdd.n92 dvss 4.46094f
C934 avdd.n93 dvss 4.48227f
C935 avdd.n94 dvss 1.19042f
C936 avdd.n95 dvss 0.66577f
C937 avdd.n96 dvss 3.27742f
C938 avdd.n97 dvss 0.20944f
C939 avdd.t0 dvss 0.702496f
C940 avdd.n98 dvss 0.20944f
C941 avdd.n99 dvss 0.731637f
C942 avdd.n100 dvss 0.757787f
C943 avdd.n101 dvss 0.146948f
C944 avdd.n103 dvss 0.303016f
C945 avss.n0 dvss 0.274689f
C946 avss.n1 dvss 0.256432f
C947 avss.n2 dvss 0.199691f
C948 avss.n4 dvss 0.10291f
C949 avss.t6 dvss 0.441575f
C950 avss.t4 dvss 0.441575f
C951 avss.n9 dvss 0.832446f
C952 avss.n10 dvss 0.117588f
C953 avss.n11 dvss 0.501337f
C954 avss.n15 dvss 0.506602f
C955 avss.n17 dvss 0.506602f
C956 avss.t22 dvss 0.441575f
C957 avss.n18 dvss 0.238935f
C958 avss.t24 dvss 0.441575f
C959 avss.n19 dvss 3.28532f
C960 avss.n20 dvss 7.3481f
C961 avss.t8 dvss 0.441575f
C962 avss.n24 dvss 0.152326f
C963 avss.n27 dvss 0.238935f
C964 avss.t10 dvss 0.441575f
C965 avss.n29 dvss 0.506602f
C966 avss.n30 dvss 0.506602f
C967 avss.t0 dvss 0.441575f
C968 avss.t2 dvss 0.441575f
C969 avss.n32 dvss 0.370586f
C970 avss.n33 dvss 0.325025f
C971 avss.n34 dvss 0.132878f
C972 avss.n35 dvss 0.404741f
C973 avss.n36 dvss 2.98049f
C974 avss.t20 dvss 0.860518f
C975 avss.t12 dvss 0.732948f
C976 avss.n37 dvss 2.16357f
C977 avss.n38 dvss 1.84584f
C978 avss.t18 dvss 0.841962f
C979 avss.t16 dvss 0.732948f
C980 avss.n39 dvss 0.3741f
C981 avss.n40 dvss 0.133098f
C982 avss.t14 dvss 0.732948f
C983 avss.n41 dvss 0.133098f
C984 avss.n42 dvss 1.68799f
C985 avss.n43 dvss 0.462717f
C986 avss.n46 dvss 1.36147f
C987 avss.n47 dvss 1.03577f
C988 avss.t26 dvss 8.17429f
C989 avss.n48 dvss 7.701231f
C990 avss.t29 dvss 8.17429f
C991 avss.n49 dvss 8.01034f
C992 avss.t28 dvss 8.17429f
C993 avss.n50 dvss 7.90618f
C994 avss.n51 dvss 4.01706f
C995 avss.t27 dvss 8.17429f
C996 avss.n52 dvss 2.18128f
C997 avss.n53 dvss 4.97729f
C998 avss.n54 dvss 1.85282f
C999 avss.n55 dvss 1.94389f
C1000 avss.n56 dvss 1.85115f
C1001 avss.n58 dvss 0.227287f
C1002 avss.n59 dvss 0.265186f
C1003 avss.n60 dvss 0.643717f
C1004 avss.n61 dvss 0.274689f
C1005 avss.n62 dvss 0.354568f
C1006 avss.n64 dvss 0.102951f
C1007 avss.n68 dvss 0.238935f
C1008 avss.n71 dvss 0.10291f
C1009 avss.n73 dvss 0.117505f
C1010 avss.n75 dvss 0.79544f
C1011 avss.n76 dvss 1.9882f
C1012 avss.n77 dvss 0.79544f
C1013 avss.n79 dvss 0.117505f
C1014 avss.n80 dvss 0.117588f
C1015 avss.n81 dvss 0.455799f
C1016 avss.n82 dvss 1.20688f
C1017 avss.n83 dvss 0.606761f
C1018 avss.n84 dvss 0.354568f
C1019 avss.n86 dvss 0.102951f
C1020 avss.n89 dvss 0.238935f
C1021 avss.n92 dvss 0.152326f
C1022 avss.n94 dvss 0.162188f
C1023 avss.n95 dvss 0.241706f
C1024 inv_in.t3 dvss 0.657711f
C1025 inv_in.t11 dvss 5.68012f
C1026 inv_in.n0 dvss 5.17707f
C1027 inv_in.t5 dvss 5.52894f
C1028 inv_in.n1 dvss 2.62426f
C1029 inv_in.t6 dvss 5.52894f
C1030 inv_in.n2 dvss 2.66147f
C1031 inv_in.n3 dvss 2.79669f
C1032 inv_in.t14 dvss 5.52894f
C1033 inv_in.n4 dvss 5.29306f
C1034 inv_in.t12 dvss 5.55261f
C1035 inv_in.n5 dvss 5.28615f
C1036 inv_in.t13 dvss 5.52894f
C1037 inv_in.n6 dvss 2.66147f
C1038 inv_in.t9 dvss 5.5836f
C1039 inv_in.n7 dvss 5.39875f
C1040 inv_in.t10 dvss 5.5836f
C1041 inv_in.t2 dvss 5.5836f
C1042 inv_in.n8 dvss 5.26653f
C1043 inv_in.n9 dvss 5.40864f
C1044 inv_in.t4 dvss 5.52894f
C1045 inv_in.n10 dvss 2.66147f
C1046 inv_in.n11 dvss 2.90209f
C1047 inv_in.n12 dvss 2.75998f
C1048 inv_in.t8 dvss 5.52894f
C1049 inv_in.n13 dvss 2.62426f
C1050 inv_in.n14 dvss 2.76492f
C1051 inv_in.n15 dvss 2.76492f
C1052 inv_in.n16 dvss 2.76201f
C1053 inv_in.t7 dvss 5.52894f
C1054 inv_in.n17 dvss 5.4592f
C1055 inv_in.n18 dvss 0.82306f
C1056 inv_in.t0 dvss 0.104143f
C1057 inv_in.t1 dvss 0.647866f
C1058 inv_in.n19 dvss 2.16816f
C1059 xout.t19 dvss 0.243993f
C1060 xout.t17 dvss 0.243993f
C1061 xout.n0 dvss 2.4243f
C1062 xout.t18 dvss 0.243993f
C1063 xout.t16 dvss 0.243993f
C1064 xout.n1 dvss 1.60432f
C1065 xout.n2 dvss 6.32987f
C1066 xout.t15 dvss 0.256529f
C1067 xout.t20 dvss 0.243993f
C1068 xout.n3 dvss 1.22843f
C1069 xout.t13 dvss 0.256529f
C1070 xout.t21 dvss 0.243993f
C1071 xout.n4 dvss 1.23308f
C1072 xout.n5 dvss 2.18555f
C1073 xout.n6 dvss 8.527769f
C1074 xout.n7 dvss 3.77761f
C1075 xout.t10 dvss 0.243993f
C1076 xout.t11 dvss 0.243993f
C1077 xout.n8 dvss 1.27442f
C1078 xout.n9 dvss 1.83376f
C1079 xout.t12 dvss 0.243993f
C1080 xout.t14 dvss 0.243993f
C1081 xout.n10 dvss 1.43377f
C1082 xout.n11 dvss 1.68066f
C1083 xout.n12 dvss 1.24537f
C1084 xout.n13 dvss 0.227228f
C1085 xout.n14 dvss 0.217681f
C1086 xout.n15 dvss 0.229174f
C1087 xout.n16 dvss 4.49086f
C1088 xout.n17 dvss 0.217681f
C1089 xout.n18 dvss 0.149204f
C1090 xout.n19 dvss 2.97025f
C1091 xout.n20 dvss 3.47714f
C1092 xout.n21 dvss 4.15788f
C1093 xout.n22 dvss 4.02374f
C1094 xout.n23 dvss 0.626416f
C1095 xout.n24 dvss 0.760656f
C1096 xout.t25 dvss 1.61622f
C1097 xout.t23 dvss 1.68073f
C1098 xout.n25 dvss 1.04327f
C1099 xout.n26 dvss 0.785936f
C1100 xout.n27 dvss 8.087669f
C1101 xout.n28 dvss 9.65943f
C1102 xout.n29 dvss 1.9924f
C1103 avdd_ip.n0 dvss 0.183001f
C1104 avdd_ip.n1 dvss 0.193101f
C1105 avdd_ip.t4 dvss 0.312571f
C1106 avdd_ip.n2 dvss 25.687199f
C1107 avdd_ip.t33 dvss 0.201546p
C1108 avdd_ip.n3 dvss 42.3367f
C1109 avdd_ip.n4 dvss 31.209301f
C1110 avdd_ip.t30 dvss 12.6155f
C1111 avdd_ip.n5 dvss 8.054391f
C1112 avdd_ip.t31 dvss 12.6155f
C1113 avdd_ip.n6 dvss 7.765079f
C1114 avdd_ip.n7 dvss 10.2323f
C1115 avdd_ip.t29 dvss 12.6155f
C1116 avdd_ip.n8 dvss 11.3223f
C1117 avdd_ip.t32 dvss 12.6155f
C1118 avdd_ip.n9 dvss 11.2988f
C1119 avdd_ip.n10 dvss 11.0453f
C1120 avdd_ip.n11 dvss 25.8585f
C1121 avdd_ip.n12 dvss 11.8125f
C1122 avdd_ip.n13 dvss 15.647901f
C1123 avdd_ip.t25 dvss 0.272851f
C1124 avdd_ip.n14 dvss 0.353227f
C1125 avdd_ip.t21 dvss 0.272851f
C1126 avdd_ip.n15 dvss 1.24555f
C1127 avdd_ip.t22 dvss 0.272851f
C1128 avdd_ip.n16 dvss 1.36471f
C1129 avdd_ip.t20 dvss 0.284354f
C1130 avdd_ip.n17 dvss 1.00481f
C1131 avdd_ip.n18 dvss 1.60279f
C1132 avdd_ip.n19 dvss 0.908877f
C1133 avdd_ip.n20 dvss 0.312041f
C1134 avdd_ip.t19 dvss 0.272851f
C1135 avdd_ip.n21 dvss 0.511759f
C1136 avdd_ip.n22 dvss 1.0293f
C1137 avdd_ip.n23 dvss 1.19091f
C1138 avdd_ip.t24 dvss 0.272851f
C1139 avdd_ip.n24 dvss 1.06873f
C1140 avdd_ip.n25 dvss 4.33929f
C1141 avdd_ip.n26 dvss 15.187299f
C1142 avdd_ip.n27 dvss 15.187299f
C1143 avdd_ip.t5 dvss 19.331099f
C1144 avdd_ip.n28 dvss 1.61496f
C1145 avdd_ip.t10 dvss 0.272851f
C1146 avdd_ip.n29 dvss 5.41016f
C1147 avdd_ip.t15 dvss 0.272851f
C1148 avdd_ip.t16 dvss 0.272851f
C1149 avdd_ip.n30 dvss 2.76186f
C1150 avdd_ip.t12 dvss 0.272851f
C1151 avdd_ip.t14 dvss 0.272851f
C1152 avdd_ip.n31 dvss 1.60468f
C1153 avdd_ip.n32 dvss 2.4602f
C1154 avdd_ip.n33 dvss 6.7614f
C1155 avdd_ip.n40 dvss 0.275331f
C1156 avdd_ip.t3 dvss 0.366056f
C1157 avdd_ip.n42 dvss -24.5529f
C1158 avdd_ip.n43 dvss 24.8309f
C1159 avdd_ip.n47 dvss 2.63147f
C1160 avdd_ip.t28 dvss 0.425863f
C1161 avdd_ip.n54 dvss 0.275331f
C1162 avdd_ip.n57 dvss 0.275331f
C1163 avdd_ip.n60 dvss 2.34174f
C1164 avdd_ip.n61 dvss 3.08369f
C1165 avdd_ip.n62 dvss 7.458549f
C1166 avdd_ip.t6 dvss 0.272851f
C1167 avdd_ip.t7 dvss 0.272851f
C1168 avdd_ip.t8 dvss 0.272851f
C1169 avdd_ip.n63 dvss 2.28083f
C1170 avdd_ip.t18 dvss 0.272851f
C1171 avdd_ip.t26 dvss 0.272851f
C1172 avdd_ip.n64 dvss 2.68748f
C1173 avdd_ip.t17 dvss 0.272851f
C1174 avdd_ip.t23 dvss 0.272851f
C1175 avdd_ip.n65 dvss 1.60335f
C1176 avdd_ip.n66 dvss 2.5326f
C1177 avdd_ip.n67 dvss 6.54556f
C1178 avdd_ip.n68 dvss 5.37955f
C1179 avdd_ip.n69 dvss 12.5401f
C1180 avdd_ip.n70 dvss 7.683919f
C1181 avdd_ip.n71 dvss 8.52327f
C1182 avdd_ip.n72 dvss 8.52327f
C1183 avdd_ip.n73 dvss 32.6198f
C1184 avdd_ip.n74 dvss 7.0648f
C1185 avdd_ip.n75 dvss 2.67542f
C1186 avdd_ip.n76 dvss 5.79729f
C1187 avdd_ip.n77 dvss 37.3139f
C1188 avdd_ip.n78 dvss 13.6449f
C1189 avdd_ip.n79 dvss 32.799896f
C1190 avdd_ip.n80 dvss 32.6198f
C1191 avdd_ip.n81 dvss 32.799896f
C1192 avdd_ip.n82 dvss 8.53496f
C1193 avdd_ip.n83 dvss 8.47481f
C1194 avdd_ip.n84 dvss 3.99638f
C1195 avdd_ip.n85 dvss 32.939102f
C1196 avdd_ip.n86 dvss 7.89575f
C1197 avdd_ip.n87 dvss 2.20458f
C1198 avdd_ip.n88 dvss 5.76955f
C1199 avdd_ip.t11 dvss 0.272851f
C1200 avdd_ip.t13 dvss 0.272851f
C1201 avdd_ip.n89 dvss 2.2737f
C1202 avdd_ip.n90 dvss 0.777352f
C1203 avdd_ip.n91 dvss 1.40119f
C1204 avdd_ip.t9 dvss 19.331099f
C1205 avdd_ip.n92 dvss 16.5454f
C1206 avdd_ip.n93 dvss 1.40119f
C1207 avdd_ip.n94 dvss 2.89538f
C1208 avdd_ip.n95 dvss 1.66736f
C1209 avdd_ip.n96 dvss 7.11433f
C1210 avdd_ip.n97 dvss 23.7224f
C1211 a_9120_n9346.t3 dvss 1.47746f
C1212 a_9120_n9346.n0 dvss 3.32132f
C1213 a_9120_n9346.t1 dvss 1.67898f
C1214 a_9120_n9346.n1 dvss 2.97825f
C1215 a_9120_n9346.n2 dvss 1.80939f
C1216 avss_ip.n0 dvss 8.051339f
C1217 avss_ip.n1 dvss 2.70068f
C1218 avss_ip.n2 dvss 4.27842f
C1219 avss_ip.n4 dvss 1.42729f
C1220 avss_ip.n7 dvss 0.51324f
C1221 avss_ip.n8 dvss 1.42254f
C1222 avss_ip.n9 dvss 4.70963f
C1223 avss_ip.n10 dvss 0.982776f
C1224 avss_ip.n11 dvss 1.16687f
C1225 avss_ip.n12 dvss 0.219239f
C1226 avss_ip.n13 dvss 0.219239f
C1227 avss_ip.n14 dvss 1.65343f
C1228 avss_ip.n15 dvss 9.4519f
C1229 avss_ip.n16 dvss 0.335032f
C1230 avss_ip.n17 dvss 0.335032f
C1231 avss_ip.n18 dvss 0.312783f
C1232 avss_ip.n19 dvss 0.548526f
C1233 avss_ip.t43 dvss 0.492215f
C1234 avss_ip.n20 dvss 0.892363f
C1235 avss_ip.n21 dvss 0.664842f
C1236 avss_ip.n22 dvss 0.139099f
C1237 avss_ip.n23 dvss 2.25351f
C1238 avss_ip.n24 dvss 4.08801f
C1239 avss_ip.n26 dvss 2.98138f
C1240 avss_ip.n27 dvss 77.2165f
C1241 avss_ip.n28 dvss 0.335895f
C1242 avss_ip.t19 dvss 14.2424f
C1243 avss_ip.n29 dvss 0.408404f
C1244 avss_ip.n30 dvss 1.0842f
C1245 avss_ip.n31 dvss 15.1282f
C1246 avss_ip.n33 dvss 1.04464f
C1247 avss_ip.n34 dvss 1.24706f
C1248 avss_ip.n38 dvss 0.729328f
C1249 avss_ip.n41 dvss 0.96204f
C1250 avss_ip.n42 dvss 1.07243f
C1251 avss_ip.n43 dvss 1.991f
C1252 avss_ip.n44 dvss 0.953578f
C1253 avss_ip.n45 dvss 0.557448f
C1254 avss_ip.n46 dvss 0.874622f
C1255 avss_ip.n47 dvss 0.3217f
C1256 avss_ip.n48 dvss 0.312892f
C1257 avss_ip.n49 dvss 3.03843f
C1258 avss_ip.n50 dvss 4.61337f
C1259 avss_ip.n51 dvss 0.837054f
C1260 avss_ip.n52 dvss 0.837054f
C1261 avss_ip.t56 dvss 29.904999f
C1262 avss_ip.t0 dvss 21.299301f
C1263 avss_ip.t55 dvss 21.8722f
C1264 avss_ip.n53 dvss 4.4065f
C1265 avss_ip.n54 dvss 4.41943f
C1266 avss_ip.n55 dvss 2.63974f
C1267 avss_ip.n56 dvss 1.8376f
C1268 avss_ip.n57 dvss 1.71471f
C1269 avss_ip.n58 dvss 3.34021f
C1270 avss_ip.n59 dvss 0.19619f
C1271 avss_ip.n60 dvss 0.204413f
C1272 avss_ip.n61 dvss 0.923648f
C1273 avss_ip.n62 dvss 0.589225f
C1274 avss_ip.n63 dvss 1.73308f
C1275 avss_ip.n64 dvss 3.17891f
C1276 avss_ip.n65 dvss 0.884422f
C1277 avss_ip.n66 dvss 2.74924f
C1278 avss_ip.t32 dvss 0.127343f
C1279 avss_ip.n69 dvss 7.05607f
C1280 avss_ip.n70 dvss 6.00621f
C1281 avss_ip.n71 dvss 1.64683f
C1282 avss_ip.n72 dvss 12.9003f
C1283 avss_ip.n73 dvss 0.255846f
C1284 avss_ip.t17 dvss 6.84807f
C1285 avss_ip.n76 dvss 15.6289f
C1286 avss_ip.n77 dvss 0.642217f
C1287 avss_ip.n78 dvss 0.826164f
C1288 avss_ip.n83 dvss 1.7246f
C1289 avss_ip.n84 dvss 0.915892f
C1290 avss_ip.n85 dvss 1.61521f
C1291 avss_ip.n88 dvss 0.494835f
C1292 avss_ip.n89 dvss 1.49255f
C1293 avss_ip.t40 dvss 0.492215f
C1294 avss_ip.n90 dvss 0.732672f
C1295 avss_ip.t57 dvss 0.152854f
C1296 avss_ip.n91 dvss 0.553655f
C1297 avss_ip.n92 dvss 0.832337f
C1298 avss_ip.n93 dvss 1.46917f
C1299 avss_ip.n94 dvss 3.48304f
C1300 avss_ip.n95 dvss 1.33455f
C1301 avss_ip.n96 dvss 1.39288f
C1302 avss_ip.n97 dvss 0.408743f
C1303 avss_ip.t46 dvss 0.492215f
C1304 avss_ip.n98 dvss 1.64809f
C1305 avss_ip.n99 dvss 0.820747f
C1306 avss_ip.n100 dvss 0.85541f
C1307 avss_ip.n101 dvss 0.653769f
C1308 avss_ip.n102 dvss 0.698156f
C1309 avss_ip.n105 dvss 1.02575f
C1310 avss_ip.n107 dvss 1.26399f
C1311 avss_ip.n108 dvss 2.38643f
C1312 avss_ip.n109 dvss 2.19901f
C1313 avss_ip.n110 dvss 0.368792f
C1314 avss_ip.n111 dvss 0.375246f
C1315 avss_ip.n112 dvss 1.22227f
C1316 avss_ip.n113 dvss 0.19555f
C1317 avss_ip.n114 dvss 2.16392f
C1318 avss_ip.n115 dvss 1.61897f
C1319 avss_ip.t53 dvss 34.1232f
C1320 avss_ip.n116 dvss 17.9534f
C1321 avss_ip.n117 dvss 8.84f
C1322 avss_ip.n119 dvss 0.255936f
C1323 avss_ip.n120 dvss 0.267718f
C1324 avss_ip.n121 dvss 0.223658f
C1325 avss_ip.n122 dvss 1.77834f
C1326 avss_ip.n123 dvss 1.32272f
C1327 avss_ip.n124 dvss 0.368792f
C1328 avss_ip.n125 dvss 0.375246f
C1329 avss_ip.n126 dvss 0.640532f
C1330 avss_ip.n127 dvss 0.853581f
C1331 avss_ip.n128 dvss 13.1621f
C1332 avss_ip.n129 dvss 3.04576f
C1333 avss_ip.n130 dvss 16.1082f
C1334 avss_ip.n131 dvss 0.112631f
C1335 avss_ip.n134 dvss 0.278947f
C1336 avss_ip.n135 dvss 0.180603f
C1337 avss_ip.n139 dvss 0.217376f
C1338 avss_ip.n140 dvss 0.137585f
C1339 avss_ip.t25 dvss 0.182183f
C1340 avss_ip.n143 dvss 1.41468f
C1341 avss_ip.n144 dvss 0.161163f
C1342 avss_ip.n145 dvss 0.36541f
C1343 avss_ip.n146 dvss 0.264843f
C1344 avss_ip.n147 dvss 0.125919f
C1345 avss_ip.n148 dvss 0.280491f
C1346 avss_ip.n152 dvss 0.557772f
C1347 avss_ip.n153 dvss 0.558375f
C1348 avss_ip.n154 dvss 0.121228f
C1349 avss_ip.n155 dvss 0.317656f
C1350 avss_ip.n157 dvss 0.453901f
C1351 avss_ip.n158 dvss 0.390992f
C1352 avss_ip.n164 dvss 0.360786f
C1353 avss_ip.n165 dvss 1.96336f
C1354 avss_ip.n166 dvss 0.765038f
C1355 avss_ip.n167 dvss 0.581965f
C1356 avss_ip.n168 dvss 0.361997f
C1357 avss_ip.n169 dvss 3.05232f
C1358 avss_ip.n170 dvss 0.12516f
C1359 avss_ip.n174 dvss 0.31412f
C1360 avss_ip.n175 dvss 0.344519f
C1361 avss_ip.n176 dvss 0.387608f
C1362 avss_ip.n177 dvss 4.53066f
C1363 avss_ip.t8 dvss 1.69249f
C1364 avss_ip.t7 dvss 3.08554f
C1365 avss_ip.n180 dvss 7.44152f
C1366 avss_ip.n181 dvss 1.04285f
C1367 avss_ip.n182 dvss 10.1046f
C1368 avss_ip.n183 dvss 11.0615f
C1369 avss_ip.n184 dvss 12.1732f
C1370 avss_ip.n185 dvss 3.69637f
C1371 avss_ip.n186 dvss 7.45136f
C1372 avss_ip.n187 dvss 0.996633f
C1373 avss_ip.n188 dvss 3.38819f
C1374 avss_ip.n189 dvss 3.85472f
C1375 avss_ip.n190 dvss 6.64403f
C1376 avss_ip.n191 dvss 2.85911f
C1377 avss_ip.n192 dvss 1.79009f
C1378 avss_ip.n193 dvss 1.70665f
C1379 avss_ip.n194 dvss 1.42818f
C1380 avss_ip.n195 dvss 0.758444f
C1381 avss_ip.n196 dvss 0.223686f
C1382 avss_ip.n197 dvss 1.45123f
C1383 avss_ip.t35 dvss 3.10202f
C1384 avss_ip.t52 dvss 3.49835f
C1385 avss_ip.n199 dvss 3.34419f
C1386 avss_ip.n200 dvss 0.106377f
C1387 avss_ip.t34 dvss 3.16236f
C1388 avss_ip.t33 dvss 3.46677f
C1389 avss_ip.n201 dvss 3.37971f
C1390 avss_ip.n202 dvss 0.41933f
C1391 avss_ip.n204 dvss 0.744701f
C1392 avss_ip.n205 dvss 0.627105f
C1393 avss_ip.n206 dvss 2.9482f
C1394 avss_ip.n207 dvss 8.53732f
C1395 avss_ip.n208 dvss 3.91375f
C1396 avss_ip.n209 dvss 3.88885f
C1397 avss_ip.n210 dvss 1.06139f
C1398 avss_ip.n211 dvss 1.39201f
C1399 avss_ip.n212 dvss 1.4208f
C1400 avss_ip.n213 dvss 0.850313f
C1401 avss_ip.n215 dvss 4.42835f
C1402 avss_ip.n217 dvss 0.135164f
C1403 avss_ip.n219 dvss 0.623135f
C1404 avss_ip.n220 dvss 0.411227f
C1405 avss_ip.n221 dvss 0.644578f
C1406 avss_ip.n222 dvss 0.642217f
C1407 avss_ip.n223 dvss 0.371146f
C1408 avss_ip.n224 dvss 0.645934f
C1409 avss_ip.n225 dvss 66.9705f
C1410 avss_ip.n226 dvss 57.3493f
C1411 avss_ip.n228 dvss 3.66196f
C1412 avss_ip.n229 dvss 4.97623f
C1413 avss_ip.n230 dvss 3.73035f
C1414 avss_ip.n231 dvss 2.43323f
C1415 avss_ip.n232 dvss 0.365839f
C1416 avss_ip.n233 dvss 2.89199f
C1417 avss_ip.n234 dvss 1.29084f
C1418 avss_ip.n235 dvss 0.450859f
C1419 avss_ip.n236 dvss 2.37447f
C1420 avss_ip.t64 dvss 56.3999f
C1421 avss_ip.t63 dvss 29.106098f
C1422 avss_ip.n237 dvss 29.2517f
C1423 avss_ip.t66 dvss 29.106098f
C1424 avss_ip.n238 dvss 28.4234f
C1425 avss_ip.t65 dvss 29.106098f
C1426 avss_ip.n239 dvss 36.5448f
C1427 avss_ip.n240 dvss 6.83647f
C1428 avss_ip.n242 dvss 0.964795f
C1429 avss_ip.n243 dvss 0.352507f
C1430 avss_ip.n244 dvss 2.74861f
C1431 avss_ip.n245 dvss 1.61511f
C1432 avss_ip.n246 dvss 0.975642f
C1433 avss_ip.n247 dvss 0.608665f
C1434 avss_ip.n248 dvss 0.556808f
C1435 avss_ip.n249 dvss 0.260543f
C1436 avss_ip.n250 dvss 4.31013f
C1437 avss_ip.n253 dvss 2.3962f
C1438 avss_ip.n254 dvss 5.26518f
C1439 avss_ip.n255 dvss 4.09586f
C1440 avss_ip.n256 dvss 3.74409f
C1441 avss_ip.n257 dvss 1.063f
C1442 avss_ip.n258 dvss 4.18646f
C1443 avss_ip.n259 dvss 0.219589f
C1444 avss_ip.n260 dvss 0.835505f
C1445 avss_ip.t3 dvss 4.2182f
C1446 avss_ip.n261 dvss 0.835505f
C1447 avss_ip.n262 dvss 1.90251f
C1448 avss_ip.n263 dvss 4.73371f
C1449 avss_ip.n264 dvss 1.04285f
C1450 avss_ip.t2 dvss 0.122789p
C1451 avss_ip.t4 dvss 9.02524f
C1452 avss_ip.n266 dvss 0.394497f
C1453 avss_ip.n267 dvss 1.03579f
C1454 avss_ip.n268 dvss 1.05611f
C1455 avss_ip.n269 dvss 1.32562f
C1456 avss_ip.n270 dvss 0.787189f
C1457 avss_ip.t49 dvss 0.492215f
C1458 avss_ip.n271 dvss 0.408743f
C1459 avss_ip.n272 dvss 0.435136f
C1460 avss_ip.n273 dvss 0.591404f
C1461 avss_ip.n274 dvss 0.603247f
C1462 avss_ip.n276 dvss 0.813399f
C1463 avss_ip.n277 dvss 0.982797f
C1464 avss_ip.n278 dvss 1.41848f
C1465 avss_ip.n279 dvss 0.730783f
C1466 avss_ip.n280 dvss 0.333717f
C1467 avss_ip.n281 dvss 10.3372f
C1468 avss_ip.n282 dvss 7.42091f
C1469 avss_ip.n283 dvss 0.217128f
C1470 avss_ip.n284 dvss 0.979986f
C1471 avss_ip.n285 dvss 0.96604f
C1472 avss_ip.n286 dvss 1.75061f
C1473 avss_ip.n287 dvss 0.103199f
C1474 avss_ip.n288 dvss 0.960797f
C1475 avss_ip.n289 dvss 1.07633f
C1476 avss_ip.n290 dvss 1.55677f
C1477 avss_ip.n291 dvss 5.11571f
C1478 avss_ip.n292 dvss 4.01697f
C1479 dvdd.n0 dvss 0.231928f
C1480 dvdd.n4 dvss 0.114981f
C1481 dvdd.n5 dvss 0.114981f
C1482 dvdd.n27 dvss 0.114981f
C1483 dvdd.n29 dvss 0.114981f
C1484 dvdd.t145 dvss 0.165457f
C1485 dvdd.n38 dvss 0.47343f
C1486 dvdd.n39 dvss 0.249961f
C1487 dvdd.t73 dvss 0.165457f
C1488 dvdd.n49 dvss 1.8472f
C1489 dvdd.t175 dvss 3.83628f
C1490 dvdd.n50 dvss 3.2293f
C1491 dvdd.n51 dvss 1.13209f
C1492 dvdd.t12 dvss 0.103953f
C1493 dvdd.t27 dvss 0.103953f
C1494 dvdd.t95 dvss 0.103953f
C1495 dvdd.n275 dvss 6.53977f
C1496 dvdd.n276 dvss 9.40408f
C1497 dvdd.t178 dvss 3.83628f
C1498 dvdd.n277 dvss 6.79779f
C1499 dvdd.t177 dvss 3.83628f
C1500 dvdd.n278 dvss 3.72992f
C1501 dvdd.t176 dvss 3.83628f
C1502 dvdd.n279 dvss 3.60793f
C1503 dvdd.n280 dvss 2.57602f
C1504 dvdd.n281 dvss 0.390563f
C1505 dvdd.n290 dvss 0.466107f
C1506 dvdd.n291 dvss 0.869136f
C1507 dvdd.n292 dvss 0.243102f
C1508 dvdd.n293 dvss 0.211035f
C1509 dvdd.t147 dvss 0.222917f
C1510 dvdd.t153 dvss 0.187598f
C1511 dvdd.t155 dvss 0.187598f
C1512 dvdd.t149 dvss 0.187598f
C1513 dvdd.t151 dvss 0.140698f
C1514 dvdd.t159 dvss 0.140698f
C1515 dvdd.t141 dvss 0.187598f
C1516 dvdd.t143 dvss 0.187598f
C1517 dvdd.t157 dvss 0.187598f
C1518 dvdd.t161 dvss 0.222917f
C1519 dvdd.n295 dvss 0.211035f
C1520 dvdd.n296 dvss 0.255981f
C1521 dvdd.n297 dvss 0.773905f
C1522 dvdd.n298 dvss 0.37474f
.ends

