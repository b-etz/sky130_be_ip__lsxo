magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< pwell >>
rect -201 -100582 201 100582
<< psubdiff >>
rect -165 100512 -69 100546
rect 69 100512 165 100546
rect -165 100450 -131 100512
rect 131 100450 165 100512
rect -165 -100512 -131 -100450
rect 131 -100512 165 -100450
rect -165 -100546 -69 -100512
rect 69 -100546 165 -100512
<< psubdiffcont >>
rect -69 100512 69 100546
rect -165 -100450 -131 100450
rect 131 -100450 165 100450
rect -69 -100546 69 -100512
<< xpolycontact >>
rect -35 99984 35 100416
rect -35 -100416 35 -99984
<< xpolyres >>
rect -35 -99984 35 99984
<< locali >>
rect -165 100512 -69 100546
rect 69 100512 165 100546
rect -165 100450 -131 100512
rect 131 100450 165 100512
rect -165 -100512 -131 -100450
rect 131 -100512 165 -100450
rect -165 -100546 -69 -100512
rect 69 -100546 165 -100512
<< viali >>
rect -19 100001 19 100398
rect -19 -100398 19 -100001
<< metal1 >>
rect -25 100398 25 100410
rect -25 100001 -19 100398
rect 19 100001 25 100398
rect -25 99989 25 100001
rect -25 -100001 25 -99989
rect -25 -100398 -19 -100001
rect 19 -100398 25 -100001
rect -25 -100410 25 -100398
<< properties >>
string FIXED_BBOX -148 -100529 148 100529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1000.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 5.715meg dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
