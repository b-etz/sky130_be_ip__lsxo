* NGSPICE file created from sky130_be_ip__lsxo_rcx.ext - technology: sky130A

.subckt sky130_be_ip__lsxo_rcx ibias dout xout xin ena avss avdd standby dvss dvdd
X0 a_16620_n1869# a_15705_n2241# a_16273_n2273# dvss.t1 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1 a_20376_n2791# x7.stby_done_b dvdd.t98 dvdd.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_21036_n1869# a_19955_n2241# a_20689_n2273# dvdd.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3 a_10620_n8338# a_24220_n8172# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X4 a_16795_n2817# a_16620_n2791# a_16974_n2791# dvss.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5 dvdd.t49 ena_ip x3.in_b dvdd.t48 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X6 dvdd.t149 a_21036_n1869# a_21211_n1943# dvdd.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_18828_n2791# a_17913_n2791# a_18481_n2549# dvss.t38 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X8 a_2130_n19848# a_24530_n20014# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X9 vbreg.t0 icnode.t1 a_11526_n12394# avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X10 x7.x2.x2.CLK a_15000_n2791# dvss.t161 dvss.t160 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X11 a_18168_n1881# x7.x1.Qb2 dvss.t189 dvss.t188 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X12 tail.t9 vbp.t3 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X13 a_16317_n2791# a_16273_n2549# a_16151_n2791# dvss.t34 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X14 dvss.t109 standby_b.t0 dvss_ip dvss.t108 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X15 a_9120_n9346.t4 a_24220_n9832# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X16 a_16795_n1943# a_16620_n1869# a_16974_n1881# dvss.t87 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X17 x7.ena_done_b.t1 a_21775_n2247# dvdd.t156 dvdd.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X18 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X19 a_20121_n2241# a_19955_n2241# dvdd.t99 dvdd.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_2130_n21176# a_24530_n21342# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X21 ibias_ip.t10 standby_33.t3 ibias.t1 ibias.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X22 xout.t18 vbreg.t9 avdd_ip.t27 avdd_ip.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X23 inv_m1 inv_in.t1 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X24 a_2132_n15590# a_18932_n15756# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X25 dout_ip.t3 inv_m2 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X26 a_20733_n2791# a_20689_n2549# a_20567_n2791# dvss.t206 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X27 inv_in.t2 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X28 x7.x1.x2.CLK a_15000_n1881# dvss.t165 dvss.t164 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X29 avdd_ip.t29 avss_ip sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X30 a_16317_n1881# a_16273_n2273# a_16151_n1869# dvss.t166 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X31 x7.stby_done_b a_21775_n2791# dvss.t18 dvss.t17 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X32 a_14009_n2701# x7.clk_disable dvss.t136 dvss.t14 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.07665 ps=0.785 w=0.42 l=0.15
X33 dvss.t12 standby_ip x4.in_b dvss.t11 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X34 dvss.t212 a_2971_n1521# ena_ip dvss.t211 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X35 dvss.t111 standby_b.t1 a_16317_n2791# dvss.t110 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X36 avdd_ip.t30 avss_ip sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X37 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X38 dvss.t19 x7.ena_done_b.t2 a_14035_n1997# dvss.t7 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X39 x7.stby_done_b a_21775_n2791# dvdd.t34 dvdd.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X40 a_2132_n17582# a_18932_n17416# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X41 inv_m1 inv_in.t3 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X42 avss.t26 avdd.t16 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X43 a_10620_n9666# a_24220_n9832# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X44 a_20733_n1881# a_20689_n2273# a_20567_n1869# dvss.t75 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X45 dvdd.t89 x7.x2.x2.CLK a_15539_n2791# dvdd.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X46 a_16782_n2425# a_15705_n2791# a_16620_n2791# dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X47 dvdd_ip inv_m1 inv_m2 dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X48 a_4857_n1521# standby.t0 dvdd.t116 dvdd.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X49 avdd_ip.t0 x3.out_b.t3 avdd.t1 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X50 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X51 a_20121_n2791# a_19955_n2791# dvss.t49 dvss.t48 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X52 dvss.t33 ena_ip a_16317_n1881# dvss.t32 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X53 x7.x1.Qb2 a_19567_n2247# dvss.t77 dvss.t76 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X54 dvss.t178 ena.t0 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X55 dvdd.t110 a_19003_n2817# a_19567_n2791# dvdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X56 avss_ip vg1.t0 vg1.t1 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X57 a_21145_n1869# a_19955_n2241# a_21036_n1869# dvss.t105 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X58 avdd_ip.t20 vbreg.t10 avdd_ip.t19 avdd_ip.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X59 a_21211_n2817# standby_b.t2 dvdd.t102 dvdd.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X60 avss_ip xin.t6 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=23.6118 ps=175.6 w=4 l=0.5
X61 a_19003_n2817# a_18828_n2791# a_19182_n2791# dvss.t78 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X62 a_15000_n1881# dout_ip.t4 dvdd.t32 dvdd.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
X63 a_2132_n17250# a_18932_n17416# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X64 a_20121_n2241# a_19955_n2241# dvss.t104 dvss.t103 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X65 dvss_ip ibias_ip.t11 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=5.8 ps=45.8 w=2 l=2
X66 a_10620_n9666# a_24220_n9500# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X67 a_18359_n1869# a_17913_n2241# a_18263_n1869# dvss.t197 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X68 xout.t17 vbreg.t11 avdd_ip.t26 avdd_ip.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X69 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=75
X70 vbreg.t2 vg2.t5 vrb.t4 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X71 a_18525_n2791# a_18481_n2549# a_18359_n2791# dvss.t137 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X72 a_2130_n20844# a_24530_n21010# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X73 a_15083_n2791# dout_ip.t5 a_15000_n2791# dvss.t16 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X74 a_21036_n1869# a_20121_n2241# a_20689_n2273# dvss.t95 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X75 dvss_ip standby_b.t3 dvss.t151 dvss.t150 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X76 a_2132_n15590# a_18932_n15424# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X77 a_14285_n2079# x7.ena_done_b.t3 a_14285_n2281# dvdd.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X78 a_19003_n1943# a_18828_n1869# a_19182_n1881# dvss.t45 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X79 vn.t2 xin.t7 vn.t1 dvdd_ip sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X80 avss.t17 standby_b.t4 standby_33.t1 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X81 a_10620_n7674# a_24220_n7840# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X82 ibias_ip.t9 ibias_ip.t8 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X83 avdd.t18 x3.out_b.t4 avdd_ip.t28 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X84 a_15960_n2791# x7.x2.Qb1 dvdd.t128 dvdd.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X85 a_2130_n19516# a_24530_n19682# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X86 xin.t8 avdd_ip.t5 sky130_fd_pr__diode_pd2nw_05v5 perim=1.8e+06 area=2.025e+11
X87 a_20579_n2247# ena_ip dvdd.t47 dvdd.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X88 dvdd.t173 a_2971_n1521# ena_ip dvdd.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X89 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X90 a_15083_n1881# dout_ip.t6 a_15000_n1881# dvss.t174 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X91 a_18525_n1881# a_18481_n2273# a_18359_n1869# dvss.t50 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X92 a_18168_n2791# x7.x2.Qb2 dvdd.t107 dvdd.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X93 dvss.t153 standby_b.t5 a_18525_n2791# dvss.t152 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X94 xin_buf xout.t23 tail.t10 dvdd_ip sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X95 a_16273_n2549# a_16055_n2791# dvdd.t101 dvdd.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X96 dvss.t101 x7.stby_done_b a_15083_n2791# dvss.t100 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X97 xout.t8 xin.t9 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X98 x7.x1.x4.Q a_21211_n1943# dvss.t184 dvss.t183 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X99 dvdd.t97 x7.stby_done_b a_15000_n2791# dvdd.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X100 a_14009_n2404# standby_ip a_14285_n2079# dvdd.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X101 dvss_ip standby_b.t6 dvss.t113 dvss.t112 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X102 avdd_ip.t21 vbreg.t12 xout.t16 avdd_ip.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X103 tail.t8 vbp.t4 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X104 a_2130_n20844# a_24530_n20678# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X105 a_16729_n1869# a_15539_n2241# a_16620_n1869# dvss.t74 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X106 avss_ip vg2.t4 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X107 dvdd_ip vbp.t5 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=19.865 ps=155.56 w=2 l=2
X108 a_16273_n2273# a_16055_n1869# dvdd.t169 dvdd.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X109 a_2132_n15258# a_18932_n15424# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X110 a_18990_n2425# a_17913_n2791# a_18828_n2791# dvdd.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X111 a_14285_n2281# x7.stby_done_b dvdd.t96 dvdd.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X112 avdd_ip.t25 vbreg.t13 avdd_ip.t24 avdd_ip.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X113 dvss.t31 ena_ip a_18525_n1881# dvss.t30 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X114 dvdd.t162 a_21211_n1943# a_21775_n2247# dvdd.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X115 dvss.t91 x7.ena_done_b.t4 a_15083_n1881# dvss.t90 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X116 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X117 a_16795_n1943# ena_ip dvdd.t45 dvdd.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X118 dvss.t13 standby.t1 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X119 dvss.t115 standby_b.t7 dvss_ip dvss.t114 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X120 a_2130_n19516# a_24530_n19350# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X121 dvdd.t94 a_14009_n2404# x7.clk_disable dvdd.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X122 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X123 dvdd_ip standby_ip dvdd.t29 dvdd.t28 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X124 a_16163_n2247# ena_ip dvdd.t43 dvdd.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X125 a_2132_n16918# a_18932_n17084# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X126 dvdd.t105 x7.x2.Qb2 a_19955_n2791# dvdd.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X127 a_19003_n1943# ena_ip dvdd.t41 dvdd.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X128 inv_in.t4 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X129 a_10620_n9334# a_24220_n9500# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X130 dvss.t195 a_21211_n2817# a_21775_n2791# dvss.t194 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X131 a_3134_n13324# vrb.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=75
X132 dvdd_ip standby_ip dvdd.t27 dvdd.t26 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X133 a_16974_n2791# standby_b.t8 dvss.t117 dvss.t116 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X134 x7.x1.x2.Q a_16795_n1943# dvss.t173 dvss.t172 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X135 a_2132_n17582# a_18932_n17748# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X136 dvdd.t174 x7.x1.x2.CLK a_15539_n2241# dvdd.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X137 dvdd_ip vbp.t6 tail.t7 dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X138 a_19182_n2791# standby_b.t9 dvss.t119 dvss.t118 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X139 dvss.t129 a_19003_n2817# a_18937_n2791# dvss.t128 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X140 avss_ip avss_ip avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X141 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X142 dout_ip.t1 inv_m2 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X143 a_15705_n2791# a_15539_n2791# dvdd.t71 dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X144 avdd.t19 x3.out_b.t5 x3.out.t0 avdd.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X145 dvdd.t137 a_16795_n2817# a_16782_n2425# dvdd.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X146 dvss.t182 a_21211_n1943# a_21775_n2247# dvss.t181 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X147 xout.t5 xin.t10 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X148 avss_ip avss_ip avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X149 a_16974_n1881# ena_ip dvss.t29 dvss.t28 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X150 dvdd.t152 a_16795_n1943# a_17359_n2247# dvdd.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X151 xin.t5 a_24530_n22338# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X152 avss_ip x3.out.t3 avss.t25 avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X153 dvss.t135 x7.clk_disable dout_filt dvss.t134 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X154 a_16055_n2791# a_15539_n2791# a_15960_n2791# dvss.t54 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X155 dvdd.t25 standby_ip dvdd_ip dvdd.t24 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X156 standby_33.t0 x4.out_b.t3 avdd.t3 avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X157 a_16055_n1869# a_15705_n2241# a_15960_n1881# dvdd.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X158 dvdd_ip vbp.t7 tail.t6 dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X159 a_20471_n2791# a_20121_n2791# a_20376_n2791# dvdd.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X160 avss_ip xout.t24 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
**devattr s=257843176,88584 d=257843176,88584
X161 tail.t5 vbp.t8 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X162 dvdd.t109 a_19003_n2817# a_18990_n2425# dvdd.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X163 a_10620_n9334# a_24220_n9168# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X164 a_19182_n1881# ena_ip dvss.t27 dvss.t26 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X165 avdd_ip.t23 vbreg.t14 xout.t15 avdd_ip.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X166 avss_ip xin.t11 xout.t6 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X167 xin_buf xout.t25 xin_buf dvdd_ip sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=2.32 ps=17.16 w=4 l=2
X168 a_3134_n13324# avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=75
X169 a_21036_n2791# a_19955_n2791# a_20689_n2549# dvdd.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X170 dvss.t44 a_19003_n1943# a_18937_n1869# dvss.t43 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X171 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X172 a_18937_n2791# a_17747_n2791# a_18828_n2791# dvss.t133 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X173 dvss.t159 a_16795_n2817# a_17359_n2791# dvss.t158 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X174 a_16273_n2273# a_16055_n1869# dvss.t199 dvss.t198 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X175 dvdd.t87 a_16620_n1869# a_16795_n1943# dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X176 x7.x1.x2.Q a_16795_n1943# dvdd.t151 dvdd.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X177 a_2130_n20512# a_24530_n20678# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X178 avss_ip xin.t12 xout.t21 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X179 dvdd.t163 a_21036_n2791# a_21211_n2817# dvdd.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X180 x4.out_b.t1 standby_ip avss.t3 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X181 a_18481_n2549# a_18263_n2791# dvdd.t142 dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X182 dvss_ip inv_m1 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=7.9025 ps=61.46 w=0.5 l=1
X183 ibias_ip.t7 ibias_ip.t6 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X184 dvss.t89 x7.x2.x2.CLK a_15539_n2791# dvss.t88 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X185 xout.t22 xin.t13 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X186 a_2132_n14926# a_18932_n15092# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X187 dvdd.t120 x7.clk_disable a_14357_n2743# dvdd.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.005 as=0.0672 ps=0.85 w=0.64 l=0.15
X188 vn.t7 vn.t5 vn.t6 dvss_ip sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X189 a_20567_n2791# a_20121_n2791# a_20471_n2791# dvss.t201 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X190 dvdd.t23 standby_ip dvdd_ip dvdd.t22 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X191 dvss_ip dout_filt dout.t0 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=1
X192 a_20471_n1869# a_19955_n2241# a_20376_n1881# dvss.t102 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X193 a_18481_n2273# a_18263_n1869# dvdd.t7 dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X194 avss.t9 x3.out.t4 avss_ip avss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X195 dvss.t171 a_16795_n1943# a_17359_n2247# dvss.t170 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X196 x7.x1.Qb1 a_17359_n2247# dvdd.t129 dvdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X197 dvdd_ip vbp.t9 tail.t4 dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X198 avss.t27 avdd.t15 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X199 x7.x2.x2.Q a_16795_n2817# dvdd.t135 dvdd.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X200 a_14035_n2743# dout_ip.t7 dout_filt dvss.t14 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X201 dvss.t214 x7.x1.x2.CLK a_15539_n2241# dvss.t213 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X202 dout_ip.t0 inv_m2 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X203 xin_buf vn.t8 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X204 avdd_ip.t22 vbreg.t15 vg1.t3 avdd_ip.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X205 a_2130_n19848# a_24530_n19682# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X206 vrb.t3 vg2.t6 vbreg.t5 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X207 a_18828_n1869# a_17913_n2241# a_18481_n2273# dvss.t196 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X208 x7.x2.Qb1 a_17359_n2791# dvss.t4 dvss.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X209 a_2130_n20512# a_24530_n20346# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X210 dvdd.t82 a_20689_n2273# a_20579_n2247# dvdd.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X211 x7.x1.x2.CLK a_15000_n1881# dvdd.t143 dvdd.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X212 dvdd_ip standby_ip dvdd.t21 dvdd.t20 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X213 a_2132_n14926# a_18932_n14760# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X214 x7.x2.Qb1 a_17359_n2791# dvdd.t5 dvdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X215 x7.x1.x3.Q a_19003_n1943# dvss.t42 dvss.t41 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X216 xout.t0 xin.t14 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X217 avdd.t10 x3.out_b.t6 avdd_ip.t3 avdd.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X218 a_16273_n2549# a_16055_n2791# dvss.t107 dvss.t106 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X219 a_16151_n2791# a_15705_n2791# a_16055_n2791# dvss.t56 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X220 vg1.t4 xin.t4 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X221 avss_ip xin.t15 xout.t1 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X222 dvss_ip inv_m1 inv_m2 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X223 a_2130_n19184# a_24530_n19018# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X224 dvdd_ip vbp.t10 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X225 inv_in.t5 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X226 dvdd.t155 a_4857_n1521# standby_ip dvdd.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X227 a_14035_n1997# ena_ip a_14009_n2404# dvss.t7 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X228 a_17913_n2791# a_17747_n2791# dvdd.t114 dvdd.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X229 a_4857_n1521# standby.t2 dvss.t36 dvss.t35 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X230 a_10620_n9002# a_24220_n9168# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X231 a_18263_n2791# a_17747_n2791# a_18168_n2791# dvss.t132 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X232 a_14009_n2404# standby_b.t10 a_14035_n2281# dvss.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X233 a_16620_n1869# a_15539_n2241# a_16273_n2273# dvdd.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X234 a_18263_n1869# a_17913_n2241# a_18168_n1881# dvdd.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X235 a_10620_n9002# a_24220_n8836# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X236 dvdd.t165 x7.x1.Qb2 a_19955_n2241# dvdd.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X237 a_2130_n20180# a_24530_n20346# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X238 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X239 x3.out_b.t2 x3.out.t5 avdd.t7 avdd.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X240 xout.t2 xin.t16 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X241 avdd.t8 standby_33.t4 x4.out_b.t2 avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X242 a_20579_n2247# a_19955_n2241# a_20471_n1869# dvdd.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X243 dvdd.t144 a_16273_n2273# a_16163_n2247# dvdd.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X244 a_15000_n2791# dout_ip.t8 dvdd.t153 dvdd.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
X245 dvdd.t61 a_18828_n1869# a_19003_n1943# dvdd.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X246 a_2130_n22172# a_24530_n22006# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X247 avss_ip xin.t17 xout.t3 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X248 avdd_ip.t31 avss_ip sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X249 a_15705_n2241# a_15539_n2241# dvdd.t79 dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X250 a_2130_n21840# a_24530_n22006# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X251 avdd_ip.t18 vbreg.t16 xout.t14 avdd_ip.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X252 dvdd.t127 x7.x2.Qb1 a_17747_n2791# dvdd.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X253 a_2132_n16586# a_18932_n16420# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X254 avss_ip xin.t18 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X255 a_10620_n8670# a_24220_n8836# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X256 xin_buf vn.t9 xin_buf dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=2.32 ps=17.16 w=4 l=2
X257 x7.x1.Qb2 a_19567_n2247# dvdd.t84 dvdd.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X258 a_2132_n17250# a_18932_n17084# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X259 a_14009_n2701# x7.clk_disable dvdd.t118 dvdd.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.10855 ps=1.005 w=0.42 l=0.15
X260 dvss.t123 x7.x2.Qb2 a_19955_n2791# dvss.t122 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X261 dvss.t10 standby_ip x7.clkin dvss.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X262 dvss_ip ibias_ip.t12 vbp.t2 dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X263 inv_in.t6 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X264 a_22601_n15524.t1 vbreg.t17 a_22601_n15524.t0 avdd_ip.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X265 a_20579_n2425# standby_b.t11 dvdd.t103 dvdd.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X266 a_16163_n2247# a_15539_n2241# a_16055_n1869# dvdd.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X267 avss_ip xin.t19 xout.t4 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X268 x7.x2.Qb2 a_19567_n2791# dvss.t86 dvss.t85 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X269 vbreg.t4 vg1.t5 vbreg.t3 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X270 vg1.t6 xin.t3 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X271 avss_ip x3.out.t6 avss.t11 avss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X272 x3.in_b ena_ip dvss.t25 dvss.t24 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X273 x7.x2.Qb2 a_19567_n2791# dvdd.t86 dvdd.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X274 dvss.t187 x7.x1.Qb2 a_19955_n2241# dvss.t186 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X275 a_15705_n2791# a_15539_n2791# dvss.t53 dvss.t52 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X276 standby_33.t2 standby_b.t12 avss.t15 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X277 vbreg.t6 vg2.t7 vrb.t2 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X278 tail.t11 xin.t20 vn.t0 dvdd_ip sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X279 dout_ip.t2 inv_m2 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X280 dvdd.t175 dvss.t202 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X281 dvdd.t160 a_21211_n1943# a_21198_n2247# dvdd.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X282 a_2130_n20180# a_24530_n20014# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X283 dvdd_ip vbp.t11 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X284 a_20376_n2791# x7.stby_done_b dvss.t99 dvss.t98 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X285 a_18828_n1869# a_17747_n2241# a_18481_n2273# dvdd.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X286 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X287 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X288 a_16795_n2817# standby_b.t13 dvdd.t130 dvdd.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X289 a_2132_n14594# a_18932_n14428# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X290 a_15705_n2241# a_15539_n2241# dvss.t73 dvss.t72 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X291 x3.out.t2 x3.in_b avss.t23 avss.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X292 a_16163_n2425# standby_b.t14 dvdd.t131 dvdd.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X293 inv_in.t7 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X294 a_2132_n15258# a_18932_n15092# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X295 a_19003_n2817# standby_b.t15 dvdd.t72 dvdd.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X296 dvdd.t67 a_18481_n2273# a_18371_n2247# dvdd.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X297 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X298 a_20376_n1881# x7.ena_done_b.t5 dvss.t93 dvss.t92 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X299 dvdd_ip inv_m1 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=1
X300 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X301 dvss.t60 standby_b.t16 dvss_ip dvss.t59 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X302 vg1.t7 xin.t2 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X303 a_2130_n19184# a_24530_n19350# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X304 a_10620_n8670# a_24220_n8504# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X305 a_17913_n2241# a_17747_n2241# dvdd.t171 dvdd.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X306 x7.x2.x4.Q a_21211_n2817# dvss.t193 dvss.t192 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X307 dvss_ip ibias_ip.t4 ibias_ip.t5 dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X308 a_21198_n2247# a_20121_n2241# a_21036_n1869# dvdd.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X309 a_20689_n2273# a_20471_n1869# dvss.t139 dvss.t138 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X310 x7.x1.x4.Q a_21211_n1943# dvdd.t158 dvdd.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X311 xout.t20 vbreg.t18 xout.t19 avdd_ip.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X312 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X313 a_2132_n16918# a_18932_n16752# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X314 avss_ip vg2.t3 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X315 a_16055_n2791# a_15705_n2791# a_15960_n2791# dvdd.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X316 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=75
X317 avss.t21 x3.in_b x3.out.t1 avss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X318 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X319 dvss_ip standby_b.t17 dvss.t62 dvss.t61 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X320 a_18371_n2247# ena_ip dvdd.t39 dvdd.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X321 a_2130_n21508# a_24530_n21674# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X322 a_18371_n2247# a_17747_n2241# a_18263_n1869# dvdd.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X323 vbreg.t8 vbreg.t7 avdd_ip.t17 avdd_ip.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X324 a_16620_n2791# a_15705_n2791# a_16273_n2549# dvss.t55 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X325 x7.x2.x4.Q a_21211_n2817# dvdd.t168 dvdd.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X326 dvdd.t3 a_16620_n2791# a_16795_n2817# dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X327 dvss_ip standby_b.t18 dvss.t80 dvss.t79 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X328 a_2130_n22172# a_24530_n22338# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X329 a_10620_n8338# a_24220_n8504# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X330 dvdd.t126 x7.x1.Qb1 a_17747_n2241# dvdd.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X331 dvdd.t19 standby_ip dvdd_ip dvdd.t18 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X332 inv_in.t8 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X333 a_2132_n16586# a_18932_n16752# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X334 a_17913_n2791# a_17747_n2791# dvss.t131 dvss.t130 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X335 a_16055_n1869# a_15539_n2241# a_15960_n1881# dvss.t71 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X336 x7.x2.x2.Q a_16795_n2817# dvss.t157 dvss.t156 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X337 avdd_ip.t32 avss_ip sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X338 x7.ena_done_b.t0 a_21775_n2247# dvss.t177 dvss.t176 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X339 avss_ip vg2.t2 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X340 avss_ip avss_ip avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X341 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X342 a_20689_n2549# a_20471_n2791# dvss.t70 dvss.t69 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X343 dvss.t82 standby_b.t19 dvss_ip dvss.t81 sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X344 dvdd.t59 a_19003_n1943# a_19567_n2247# dvdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X345 dvdd_ip a_9120_n9346.t2 a_9120_n9346.t3 dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X346 dvdd.t167 a_21211_n2817# a_21775_n2791# dvdd.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X347 a_20376_n1881# x7.ena_done_b.t6 dvdd.t76 dvdd.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X348 a_18937_n1869# a_17747_n2241# a_18828_n1869# dvss.t210 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X349 avss_ip xin.t21 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
**devattr s=257843176,88584 d=257843176,88584
X350 dvdd_ip vbp.t12 tail.t3 dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X351 a_21211_n2817# a_21036_n2791# a_21390_n2791# dvss.t185 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X352 tail.t2 vbp.t13 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X353 a_17913_n2241# a_17747_n2241# dvss.t209 dvss.t208 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X354 dvdd.t170 a_20689_n2549# a_20579_n2425# dvdd.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X355 dvdd_ip standby_ip dvdd.t17 dvdd.t16 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X356 a_20567_n1869# a_20121_n2241# a_20471_n1869# dvss.t94 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X357 dvdd.t176 dvss.t203 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X358 dvss.t127 a_19003_n2817# a_19567_n2791# dvss.t126 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X359 a_18481_n2273# a_18263_n1869# dvss.t6 dvss.t5 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X360 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X361 dvss_ip vn.t3 vn.t4 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X362 a_2130_n18852# a_24530_n19018# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X363 dvss.t147 x7.x2.Qb1 a_17747_n2791# dvss.t146 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X364 dvdd.t177 dvss.t204 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X365 avss.t28 avdd.t14 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X366 avss.t1 standby_ip x4.out_b.t0 avss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X367 icnode.t0 vg2.t8 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X368 avdd_ip.t16 vbreg.t19 xout.t13 avdd_ip.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X369 a_21211_n1943# a_21036_n1869# a_21390_n1881# dvss.t167 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X370 a_15960_n2791# x7.x2.Qb1 dvss.t145 dvss.t144 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X371 a_11526_n12394# icnode.t1 a_8268_n12482.t0 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X372 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X373 dvss.t40 a_19003_n1943# a_19567_n2247# dvss.t39 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X374 xout.t12 vbreg.t20 avdd_ip.t15 avdd_ip.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X375 dvss.t175 a_4857_n1521# standby_ip dvss.t35 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X376 a_14009_n2404# standby_ip dvss.t8 dvss.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X377 inv_in.t9 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X378 dvdd_ip vbp.t0 vbp.t1 dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X379 a_2132_n14594# a_18932_n14760# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X380 a_16620_n2791# a_15539_n2791# a_16273_n2549# dvdd.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X381 dvss.t143 x7.x1.Qb1 a_17747_n2241# dvss.t142 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X382 a_18263_n2791# a_17913_n2791# a_18168_n2791# dvdd.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X383 dvdd.t133 a_16795_n2817# a_17359_n2791# dvdd.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X384 a_2971_n1521# ena.t1 dvss.t58 dvss.t57 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X385 dvss.t84 standby_b.t20 a_20733_n2791# dvss.t83 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X386 a_15960_n1881# x7.x1.Qb1 dvss.t141 dvss.t140 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X387 a_14035_n2281# x7.stby_done_b dvss.t97 dvss.t7 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X388 a_20579_n2425# a_19955_n2791# a_20471_n2791# dvdd.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X389 a_21145_n2791# a_19955_n2791# a_21036_n2791# dvss.t47 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X390 dvdd.t51 a_16273_n2549# a_16163_n2425# dvdd.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X391 a_16151_n1869# a_15705_n2241# a_16055_n1869# dvss.t0 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X392 a_2130_n18852# xout.t7 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X393 dvdd.t85 a_18828_n2791# a_19003_n2817# dvdd.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X394 a_16782_n2247# a_15705_n2241# a_16620_n1869# dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X395 x3.out_b.t1 ena_ip avss.t7 avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X396 dvss.t96 a_14009_n2404# x7.clk_disable dvss.t7 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X397 avss.t29 avdd.t13 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X398 dvdd.t15 standby_ip dvdd_ip dvdd.t14 sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X399 a_18481_n2549# a_18263_n2791# dvss.t163 dvss.t162 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X400 a_18359_n2791# a_17913_n2791# a_18263_n2791# dvss.t37 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X401 avdd_ip.t4 x3.out_b.t7 avdd.t12 avdd.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X402 a_18263_n1869# a_17747_n2241# a_18168_n1881# dvss.t207 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X403 dvss.t23 ena_ip a_20733_n1881# dvss.t22 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X404 x7.x2.x3.Q a_19003_n2817# dvss.t125 dvss.t124 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X405 xout.t11 vbreg.t21 avdd_ip.t14 avdd_ip.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X406 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X407 x7.x1.x3.Q a_19003_n1943# dvdd.t57 dvdd.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X408 a_21036_n2791# a_20121_n2791# a_20689_n2549# dvss.t200 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X409 dvss.t64 standby_b.t21 dvss_ip dvss.t63 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X410 avdd_ip.t33 icnode.t1 sky130_fd_pr__cap_mim_m3_1 l=20 w=20
X411 a_21211_n1943# ena_ip dvdd.t37 dvdd.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X412 inv_in.t10 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X413 inv_in.t11 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X414 a_10620_n8006# a_24220_n8172# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X415 avdd_ip.t13 vbreg.t22 xout.t10 avdd_ip.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X416 a_2130_n21840# a_24530_n21674# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X417 inv_in.t12 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X418 a_10620_n8006# a_24220_n7840# dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X419 avdd.t5 x3.out_b.t8 avdd_ip.t1 avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X420 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X421 avss.t5 ena_ip x3.out_b.t0 avss.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X422 a_2132_n16254# a_18932_n16420# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X423 a_16163_n2425# a_15539_n2791# a_16055_n2791# dvdd.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X424 tail.t1 vbp.t14 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X425 a_8268_n12482.t0 a_8268_n12482.t1 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X426 x7.x2.x3.Q a_19003_n2817# dvdd.t108 dvdd.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X427 dvss.t15 a_14009_n2701# a_14035_n2743# dvss.t14 sky130_fd_pr__nfet_01v8 ad=0.07665 pd=0.785 as=0.0441 ps=0.63 w=0.42 l=0.15
X428 x7.x2.x2.CLK a_15000_n2791# dvdd.t139 dvdd.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X429 dvdd_ip vbp.t15 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X430 a_21390_n2791# standby_b.t22 dvss.t66 dvss.t65 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X431 dvss.t191 a_21211_n2817# a_21145_n2791# dvss.t190 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X432 vg1.t8 xin.t1 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X433 dvss_ip standby_b.t23 dvss.t68 dvss.t67 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X434 inv_in.t13 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X435 a_16729_n2791# a_15539_n2791# a_16620_n2791# dvss.t51 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X436 a_9120_n9346.t1 a_9120_n9346.t0 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X437 a_2130_n21176# a_24530_n21010# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X438 a_2132_n17914# vg1.t2 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X439 a_15960_n1881# x7.x1.Qb1 dvdd.t124 dvdd.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X440 a_20121_n2791# a_19955_n2791# dvdd.t63 dvdd.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X441 dvdd.t166 a_21211_n2817# a_21198_n2425# dvdd.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X442 a_14357_n2743# dout_ip.t9 dout_filt dvdd.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X443 a_2971_n1521# ena.t2 dvdd.t141 dvdd.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X444 a_21390_n1881# ena_ip dvss.t21 dvss.t20 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X445 x4.in_b standby_ip dvdd.t13 dvdd.t12 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X446 dvss_ip ibias_ip.t2 ibias_ip.t3 dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X447 avss_ip x3.out.t7 avss.t13 avss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X448 a_18828_n2791# a_17747_n2791# a_18481_n2549# dvdd.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X449 a_18168_n1881# x7.x1.Qb2 dvdd.t164 dvdd.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X450 dvdd.t178 dvss.t205 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X451 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X452 dvss.t180 a_21211_n1943# a_21145_n1869# dvss.t179 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X453 a_14285_n2281# ena_ip a_14285_n2079# dvdd.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X454 avdd_ip.t12 vbreg.t23 avdd_ip.t11 avdd_ip.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X455 a_2132_n16254# a_18932_n16088# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X456 a_20689_n2549# a_20471_n2791# dvdd.t74 dvdd.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X457 dvdd.t78 x7.ena_done_b.t7 a_15000_n1881# dvdd.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X458 dvdd.t146 standby_b.t24 a_14285_n2281# dvdd.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X459 dvdd.t121 a_18481_n2549# a_18371_n2425# dvdd.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X460 dvdd_ip vbp.t16 tail.t0 dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X461 xout.t9 vbreg.t24 avdd_ip.t9 avdd_ip.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X462 a_18990_n2247# a_17913_n2241# a_18828_n1869# dvdd.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X463 a_20689_n2273# a_20471_n1869# dvdd.t122 dvdd.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X464 dvss_ip ibias_ip.t13 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X465 vg1.t9 xin.t0 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X466 avss.t19 x3.out.t8 avss_ip avss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X467 avss_ip avss_ip avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X468 a_2132_n17914# a_18932_n17748# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X469 a_2132_n14262# a_18932_n14428# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X470 a_21198_n2425# a_20121_n2791# a_21036_n2791# dvdd.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X471 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X472 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X473 dvss.t155 a_16795_n2817# a_16729_n2791# dvss.t154 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X474 inv_in.t14 xin_buf sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X475 dvdd_ip vbp.t17 dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X476 dvdd_ip standby_ip dvdd.t11 dvdd.t10 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X477 avss_ip vg2.t1 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X478 a_2132_n15922# a_18932_n16088# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X479 a_18371_n2425# standby_b.t25 dvdd.t147 dvdd.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X480 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X481 a_18371_n2425# a_17747_n2791# a_18263_n2791# dvdd.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X482 ibias_ip.t1 ibias_ip.t0 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X483 dvss.t169 a_16795_n1943# a_16729_n1869# dvss.t168 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X484 dout.t1 dout_filt dvdd_ip dvdd_ip sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X485 a_2132_n14262# vg2.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X486 dvdd.t150 a_16795_n1943# a_16782_n2247# dvdd.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X487 avdd_ip.t8 vbreg.t25 avdd_ip.t7 avdd_ip.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X488 xout.t26 avdd_ip.t2 sky130_fd_pr__diode_pd2nw_05v5 perim=1.8e+06 area=2.025e+11
X489 a_20471_n2791# a_19955_n2791# a_20376_n2791# dvss.t46 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X490 x7.x1.Qb1 a_17359_n2247# dvss.t149 dvss.t148 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X491 a_20471_n1869# a_20121_n2241# a_20376_n1881# dvdd.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X492 dvdd.t9 standby_ip dvdd_ip dvdd.t8 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X493 a_2130_n21508# a_24530_n21342# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X494 a_10620_n7674# inv_in.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X495 dvdd.t55 a_19003_n1943# a_18990_n2247# dvdd.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X496 dvdd_ip dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X497 a_18168_n2791# x7.x2.Qb2 dvss.t121 dvss.t120 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X498 vrb.t1 vg2.t9 vbreg.t1 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X499 a_2132_n15922# a_18932_n15756# avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
R0 dvss.n623 dvss.n622 844724
R1 dvss.n146 dvss.n145 148018
R2 dvss.n650 dvss.n17 121073
R3 dvss.n144 dvss.n44 20785.4
R4 dvss.n145 dvss.n144 13161.6
R5 dvss.n43 dvss.n42 10590.5
R6 dvss.n142 dvss.n40 8607.23
R7 dvss.n562 dvss.n546 8366.71
R8 dvss.n546 dvss.n92 8366.71
R9 dvss.n544 dvss.n92 8366.71
R10 dvss.n562 dvss.n544 8366.71
R11 dvss.n613 dvss.n612 5881.35
R12 dvss.n88 dvss.n40 5784.65
R13 dvss.n624 dvss.n31 5227.07
R14 dvss.n32 dvss.n31 5083.5
R15 dvss.n612 dvss.n44 4954.5
R16 dvss.n229 dvss.n227 4604.94
R17 dvss.n603 dvss.n44 4392.82
R18 dvss.n101 dvss.n93 4247.09
R19 dvss.n541 dvss.n93 4247.09
R20 dvss.n101 dvss.n94 4247.09
R21 dvss.n541 dvss.n94 4247.09
R22 dvss.n213 dvss.n206 4247.09
R23 dvss.n218 dvss.n206 4247.09
R24 dvss.n213 dvss.n207 4247.09
R25 dvss.n218 dvss.n207 4247.09
R26 dvss.n623 dvss.n32 3898.89
R27 dvss.n622 dvss.n621 3764.56
R28 dvss.n625 dvss.n624 3697.38
R29 dvss.n227 dvss.n90 3234.36
R30 dvss.n29 dvss.n15 2798.56
R31 dvss.n653 dvss.n15 2798.56
R32 dvss.n29 dvss.n16 2798.56
R33 dvss.n653 dvss.n16 2798.56
R34 dvss.n589 dvss.n55 2798.56
R35 dvss.n56 dvss.n55 2798.56
R36 dvss.n589 dvss.n60 2798.56
R37 dvss.n60 dvss.n56 2798.56
R38 dvss.n543 dvss.n542 2575.49
R39 dvss.n624 dvss.n623 2562.64
R40 dvss.n613 dvss.n43 2543.9
R41 dvss.n233 dvss.n83 2397.52
R42 dvss.n303 dvss.n302 2387.64
R43 dvss.n436 dvss.n146 2316.35
R44 dvss.n143 dvss.n142 2162.81
R45 dvss.n566 dvss.n90 2000.34
R46 dvss.n649 dvss.n18 1686.66
R47 dvss.n304 dvss.n303 1680.95
R48 dvss.n630 dvss.n626 1407.97
R49 dvss.n636 dvss.n626 1407.97
R50 dvss.n636 dvss.n627 1407.97
R51 dvss.n586 dvss.n62 1407.97
R52 dvss.n70 dvss.n62 1407.97
R53 dvss.n586 dvss.n63 1407.97
R54 dvss.n70 dvss.n63 1407.97
R55 dvss.n34 dvss.n32 1313.59
R56 dvss.n681 dvss.n0 1212.38
R57 dvss.n588 dvss.n61 1202.51
R58 dvss.n220 dvss.n7 1198.25
R59 dvss.n302 dvss.n301 1198.25
R60 dvss.n289 dvss.n235 1198.25
R61 dvss.n518 dvss.n109 1198.25
R62 dvss.n478 dvss.n126 1198.25
R63 dvss.n438 dvss.n437 1198.25
R64 dvss.n435 dvss.n434 1198.25
R65 dvss.n209 dvss.n164 1198.25
R66 dvss.n210 dvss.n181 1198.25
R67 dvss.n315 dvss.n200 1198.25
R68 dvss.n305 dvss.n304 1198.25
R69 dvss.n639 dvss.n638 1198.25
R70 dvss.n73 dvss.n72 1198.25
R71 dvss.n651 dvss.n650 1184.03
R72 dvss.n681 dvss.n680 1175.19
R73 dvss.n615 dvss.n35 1127.15
R74 dvss.n42 dvss.n41 1064.88
R75 dvss.t92 dvss.t103 935.78
R76 dvss.t188 dvss.t208 935.78
R77 dvss.t140 dvss.t72 935.78
R78 dvss.n574 dvss.n85 927.908
R79 dvss.n145 dvss.n49 900.194
R80 dvss.n620 dvss.n35 884.347
R81 dvss.n554 dvss.n553 784.03
R82 dvss.n561 dvss.n560 783.962
R83 dvss.n553 dvss.n552 783.75
R84 dvss.n561 dvss.n551 783.683
R85 dvss.n235 dvss.t164 748.625
R86 dvss.n614 dvss.n613 720.655
R87 dvss.t48 dvss.t98 717.851
R88 dvss.t130 dvss.t120 717.851
R89 dvss.t181 dvss.t183 689.909
R90 dvss.t183 dvss.t167 689.909
R91 dvss.t39 dvss.t41 689.909
R92 dvss.t41 dvss.t45 689.909
R93 dvss.t172 dvss.t170 689.909
R94 dvss.t87 dvss.t172 689.909
R95 dvss.n211 dvss.t52 655.918
R96 dvss.n652 dvss.n651 639.12
R97 dvss.n598 dvss.n597 626.816
R98 dvss.n30 dvss.t24 618.75
R99 dvss.n652 dvss.t24 618.75
R100 dvss.t75 dvss.t94 609.174
R101 dvss.t50 dvss.t197 609.174
R102 dvss.t0 dvss.t166 609.174
R103 dvss.n84 dvss.n81 585
R104 dvss.n84 dvss.n61 585
R105 dvss.n605 dvss.n604 585
R106 dvss.n604 dvss.n603 585
R107 dvss.n229 dvss.n107 585
R108 dvss.n229 dvss.n228 585
R109 dvss.n230 dvss.n83 585
R110 dvss.n91 dvss.n83 585
R111 dvss.n571 dvss.n570 585
R112 dvss.n572 dvss.n571 585
R113 dvss.n569 dvss.n88 585
R114 dvss.n88 dvss.n86 585
R115 dvss.t160 dvss.n200 574.28
R116 dvss.n437 dvss.t176 554.129
R117 dvss.n126 dvss.t76 554.129
R118 dvss.t148 dvss.n109 554.129
R119 dvss.t20 dvss.t179 546.789
R120 dvss.t26 dvss.t43 546.789
R121 dvss.t168 dvss.t28 546.789
R122 dvss.t192 dvss.t194 529.24
R123 dvss.t185 dvss.t192 529.24
R124 dvss.t124 dvss.t126 529.24
R125 dvss.t78 dvss.t124 529.24
R126 dvss.t156 dvss.t158 529.24
R127 dvss.t2 dvss.t156 529.24
R128 dvss.t138 dvss.t22 484.404
R129 dvss.t5 dvss.t30 484.404
R130 dvss.t32 dvss.t198 484.404
R131 dvss.t201 dvss.t206 467.307
R132 dvss.t37 dvss.t137 467.307
R133 dvss.t56 dvss.t34 467.307
R134 dvss.n615 dvss.n39 467.033
R135 dvss.t164 dvss.t90 447.707
R136 dvss.n303 dvss.n220 426.382
R137 dvss.n435 dvss.t17 425.08
R138 dvss.t85 dvss.n209 425.08
R139 dvss.t3 dvss.n210 425.08
R140 dvss.t190 dvss.t65 419.45
R141 dvss.t128 dvss.t118 419.45
R142 dvss.t154 dvss.t116 419.45
R143 dvss.n638 dvss.n637 419.18
R144 dvss.n597 dvss.n50 404.022
R145 dvss.t105 dvss.t95 400
R146 dvss.t210 dvss.t196 400
R147 dvss.t1 dvss.t74 400
R148 dvss.n630 dvss.n629 390.825
R149 dvss.t83 dvss.t69 371.594
R150 dvss.t152 dvss.t162 371.594
R151 dvss.t110 dvss.t106 371.594
R152 dvss.n651 dvss.t211 366.435
R153 dvss.t95 dvss.t138 363.303
R154 dvss.t196 dvss.t5 363.303
R155 dvss.t198 dvss.t1 363.303
R156 dvss.t176 dvss.t181 355.964
R157 dvss.t76 dvss.t39 355.964
R158 dvss.t170 dvss.t148 355.964
R159 dvss.t179 dvss.t105 352.295
R160 dvss.t94 dvss.t102 352.295
R161 dvss.t43 dvss.t210 352.295
R162 dvss.t197 dvss.t207 352.295
R163 dvss.t74 dvss.t168 352.295
R164 dvss.t102 dvss.t92 348.625
R165 dvss.t207 dvss.t188 348.625
R166 dvss.t71 dvss.t140 348.625
R167 dvss.n637 dvss.n625 344.228
R168 dvss.t100 dvss.t160 343.442
R169 dvss.n233 dvss.n229 335.039
R170 dvss.t167 dvss.t20 333.945
R171 dvss.t45 dvss.t26 333.945
R172 dvss.t28 dvss.t87 333.945
R173 dvss.n85 dvss.n84 331.606
R174 dvss.n228 dvss.t71 326.606
R175 dvss.n615 dvss.n40 310.599
R176 dvss.n41 dvss.n35 308.933
R177 dvss.n437 dvss.n436 308.257
R178 dvss.t103 dvss.t186 308.257
R179 dvss.t208 dvss.t142 308.257
R180 dvss.n638 dvss 308.139
R181 dvss.n283 dvss.t141 307.536
R182 dvss.n512 dvss.t189 307.536
R183 dvss.n472 dvss.t93 307.536
R184 dvss.n161 dvss.t99 307.536
R185 dvss.n178 dvss.t121 307.536
R186 dvss.n321 dvss.t145 307.536
R187 dvss.t200 dvss.t47 306.846
R188 dvss.t38 dvss.t133 306.846
R189 dvss.t55 dvss.t51 306.846
R190 dvss.n70 dvss.n69 292.5
R191 dvss.n71 dvss.n70 292.5
R192 dvss.n68 dvss.n63 292.5
R193 dvss.t13 dvss.n63 292.5
R194 dvss.n586 dvss.n585 292.5
R195 dvss.n587 dvss.n586 292.5
R196 dvss.n64 dvss.n62 292.5
R197 dvss.t13 dvss.n62 292.5
R198 dvss.n633 dvss.n627 292.5
R199 dvss.n636 dvss.n635 292.5
R200 dvss.n637 dvss.n636 292.5
R201 dvss.n628 dvss.n626 292.5
R202 dvss.t178 dvss.n626 292.5
R203 dvss.n631 dvss.n630 292.5
R204 dvss.t174 dvss 289.909
R205 dvss.t69 dvss.t200 278.695
R206 dvss.t162 dvss.t38 278.695
R207 dvss.t106 dvss.t55 278.695
R208 dvss.n217 dvss.n215 276.286
R209 dvss dvss.n126 275.229
R210 dvss dvss.n109 275.229
R211 dvss.n235 dvss 275.229
R212 dvss.n302 dvss 275.229
R213 dvss.t9 dvss.n0 273.678
R214 dvss.n542 dvss.t9 273.678
R215 dvss.t194 dvss.t17 273.065
R216 dvss.t126 dvss.t85 273.065
R217 dvss.t158 dvss.t3 273.065
R218 dvss.t47 dvss.t190 270.25
R219 dvss.t46 dvss.t201 270.25
R220 dvss.t133 dvss.t128 270.25
R221 dvss.t132 dvss.t37 270.25
R222 dvss.t51 dvss.t154 270.25
R223 dvss.t98 dvss.t46 267.435
R224 dvss.t120 dvss.t132 267.435
R225 dvss.t54 dvss.t144 267.435
R226 dvss.t22 dvss.t75 264.221
R227 dvss.t30 dvss.t50 264.221
R228 dvss.t166 dvss.t32 264.221
R229 dvss.t90 dvss.t174 264.221
R230 dvss.n611 dvss.n45 258.5
R231 dvss.t65 dvss.t185 256.175
R232 dvss.t118 dvss.t78 256.175
R233 dvss.t116 dvss.t2 256.175
R234 dvss.n543 dvss.t81 255.168
R235 dvss.n256 dvss.t173 246.817
R236 dvss.n485 dvss.t42 246.817
R237 dvss.n445 dvss.t184 246.817
R238 dvss.n151 dvss.t193 246.817
R239 dvss.n386 dvss.t125 246.817
R240 dvss.n347 dvss.t157 246.817
R241 dvss.t57 dvss.t211 244.291
R242 dvss.t186 dvss 238.532
R243 dvss.t142 dvss 238.532
R244 dvss dvss.t213 238.532
R245 dvss.n436 dvss.n435 236.469
R246 dvss.t122 dvss.t48 236.469
R247 dvss.t146 dvss.t130 236.469
R248 dvss.t52 dvss.t88 236.469
R249 dvss.n61 dvss.n42 236.023
R250 dvss.n588 dvss.n587 230.855
R251 dvss.n325 dvss.t135 229.185
R252 dvss.n522 dvss.n521 227.357
R253 dvss.n97 dvss.t10 219.8
R254 dvss.n540 dvss.n95 217.329
R255 dvss.n215 dvss.n214 217.225
R256 dvss.n249 dvss.n248 214.742
R257 dvss.n123 dvss.n122 214.742
R258 dvss.n140 dvss.n139 214.742
R259 dvss.n150 dvss.n149 214.742
R260 dvss.n392 dvss.n166 214.742
R261 dvss.n353 dvss.n183 214.742
R262 dvss.n571 dvss.n87 213.325
R263 dvss.n209 dvss 211.132
R264 dvss.n210 dvss 211.132
R265 dvss dvss.n200 211.132
R266 dvss.n304 dvss 211.132
R267 dvss.n263 dvss.n245 209.254
R268 dvss.n492 dvss.n119 209.254
R269 dvss.n452 dvss.n136 209.254
R270 dvss.n154 dvss.n153 209.254
R271 dvss.n172 dvss.n171 209.254
R272 dvss.n189 dvss.n188 209.254
R273 dvss.t81 dvss.t61 208.894
R274 dvss.t61 dvss.t114 208.894
R275 dvss.t114 dvss.t67 208.894
R276 dvss.t67 dvss.t63 208.894
R277 dvss.t150 dvss.t108 208.894
R278 dvss.t108 dvss.t79 208.894
R279 dvss.t59 dvss.t112 208.894
R280 dvss.n526 dvss.n525 203.619
R281 dvss.t206 dvss.t83 202.688
R282 dvss.t137 dvss.t152 202.688
R283 dvss.t34 dvss.t110 202.688
R284 dvss.t16 dvss.t100 202.688
R285 dvss.n666 dvss.n6 202.067
R286 dvss.n604 dvss.n45 202.048
R287 dvss.n3 dvss.n2 200.516
R288 dvss.n237 dvss.n236 199.739
R289 dvss.n271 dvss.n270 199.739
R290 dvss.n111 dvss.n110 199.739
R291 dvss.n500 dvss.n499 199.739
R292 dvss.n128 dvss.n127 199.739
R293 dvss.n460 dvss.n459 199.739
R294 dvss.n412 dvss.n158 199.739
R295 dvss.n399 dvss.n163 199.739
R296 dvss.n373 dvss.n175 199.739
R297 dvss.n360 dvss.n180 199.739
R298 dvss.n334 dvss.n192 199.739
R299 dvss.n199 dvss.n198 199.739
R300 dvss.n24 dvss.n23 199.739
R301 dvss.n75 dvss.n74 199.739
R302 dvss.n540 dvss.n539 198.024
R303 dvss.n587 dvss.t11 187.785
R304 dvss.n295 dvss.n294 185
R305 dvss.n205 dvss.n204 185
R306 dvss.n679 dvss.n678 185
R307 dvss dvss.t122 182.982
R308 dvss dvss.t146 182.982
R309 dvss.n28 dvss.n12 181.835
R310 dvss.n28 dvss.n27 181.835
R311 dvss.n58 dvss.n57 181.835
R312 dvss.n59 dvss.n58 181.835
R313 dvss.n629 dvss.n627 174.962
R314 dvss.n212 dvss.t54 166.091
R315 dvss.n234 dvss.t72 161.469
R316 dvss.n31 dvss.n30 155.325
R317 dvss.n219 dvss.t16 154.831
R318 dvss.n95 dvss.n93 148.029
R319 dvss.t213 dvss.n234 146.79
R320 dvss.n218 dvss.n217 146.25
R321 dvss.n219 dvss.n218 146.25
R322 dvss.n214 dvss.n213 146.25
R323 dvss.n213 dvss.n212 146.25
R324 dvss.n96 dvss.n94 146.25
R325 dvss.n94 dvss.t9 146.25
R326 dvss.n93 dvss.t9 146.25
R327 dvss.n102 dvss.n95 143.809
R328 dvss.n577 dvss.n81 143.196
R329 dvss.t35 dvss 141.269
R330 dvss.t88 dvss.t134 140.756
R331 dvss dvss.t14 140.144
R332 dvss.n545 dvss.n86 129.567
R333 dvss.n574 dvss.n83 128.583
R334 dvss.n217 dvss.n216 127.487
R335 dvss.n72 dvss.n33 122.319
R336 dvss.t112 dvss.n572 120.312
R337 dvss.n58 dvss.n56 117.001
R338 dvss.n56 dvss.n33 117.001
R339 dvss.n60 dvss.n59 117.001
R340 dvss.t11 dvss.n60 117.001
R341 dvss.n590 dvss.n589 117.001
R342 dvss.n589 dvss.n588 117.001
R343 dvss.n57 dvss.n55 117.001
R344 dvss.t11 dvss.n55 117.001
R345 dvss.n654 dvss.n653 117.001
R346 dvss.n653 dvss.n652 117.001
R347 dvss.n16 dvss.n12 117.001
R348 dvss.t24 dvss.n16 117.001
R349 dvss.n29 dvss.n28 117.001
R350 dvss.n30 dvss.n29 117.001
R351 dvss.n27 dvss.n15 117.001
R352 dvss.t24 dvss.n15 117.001
R353 dvss.n573 dvss.t79 113.703
R354 dvss.n232 dvss.n231 108.201
R355 dvss.n622 dvss.n33 105.091
R356 dvss.n212 dvss.t56 104.159
R357 dvss.n654 dvss.n13 102.025
R358 dvss.n655 dvss.n654 102.025
R359 dvss.n590 dvss.n52 102.025
R360 dvss.n590 dvss.n54 102.025
R361 dvss.n648 dvss.n19 101.874
R362 dvss.t63 dvss.n91 101.803
R363 dvss.n245 dvss.t29 100.001
R364 dvss.n119 dvss.t27 100.001
R365 dvss.n136 dvss.t21 100.001
R366 dvss.n153 dvss.t66 100.001
R367 dvss.n171 dvss.t119 100.001
R368 dvss.n188 dvss.t117 100.001
R369 dvss.n599 dvss.n598 98.4337
R370 dvss.n573 dvss.t59 95.1928
R371 dvss.n631 dvss.n628 91.4829
R372 dvss.n69 dvss.n64 91.4829
R373 dvss.n545 dvss.n43 85.938
R374 dvss.n53 dvss.t12 83.7183
R375 dvss.n646 dvss.t25 83.7183
R376 dvss.n142 dvss.n45 81.509
R377 dvss.n629 dvss.t178 81.1932
R378 dvss dvss.t57 80.5052
R379 dvss.n655 dvss.n12 79.8123
R380 dvss.n27 dvss.n13 79.8123
R381 dvss.n59 dvss.n52 79.8123
R382 dvss.n57 dvss.n54 79.8123
R383 dvss.n617 dvss.n616 73.2369
R384 dvss.n616 dvss.n615 73.1255
R385 dvss.n615 dvss.n614 73.1255
R386 dvss.n294 dvss.t165 72.8576
R387 dvss.n270 dvss.t33 72.8576
R388 dvss.n499 dvss.t31 72.8576
R389 dvss.n459 dvss.t23 72.8576
R390 dvss.n204 dvss.t161 72.8576
R391 dvss.n158 dvss.t84 72.8576
R392 dvss.n175 dvss.t153 72.8576
R393 dvss.n192 dvss.t111 72.8576
R394 dvss.n41 dvss.n39 72.01
R395 dvss.n521 dvss.n107 71.4371
R396 dvss.n245 dvss.t169 70.0005
R397 dvss.n119 dvss.t44 70.0005
R398 dvss.n136 dvss.t180 70.0005
R399 dvss.n153 dvss.t191 70.0005
R400 dvss.n171 dvss.t129 70.0005
R401 dvss.n188 dvss.t155 70.0005
R402 dvss.n69 dvss.n68 69.6045
R403 dvss.n635 dvss.n628 69.0306
R404 dvss dvss.t13 68.912
R405 dvss.n208 dvss.n196 68.8106
R406 dvss dvss.n219 67.5629
R407 dvss.n585 dvss.n64 66.3131
R408 dvss.n632 dvss.n631 65.475
R409 dvss.n527 dvss.n526 64.5768
R410 dvss.n564 dvss.t150 63.462
R411 dvss.t144 dvss.n211 61.9327
R412 dvss.n270 dvss.t199 60.5809
R413 dvss.n499 dvss.t6 60.5809
R414 dvss.n459 dvss.t139 60.5809
R415 dvss.n158 dvss.t70 60.5809
R416 dvss.n175 dvss.t163 60.5809
R417 dvss.n192 dvss.t107 60.5809
R418 dvss.n294 dvss.t91 58.5719
R419 dvss.n204 dvss.t101 58.5719
R420 dvss.n619 dvss.n617 57.4606
R421 dvss.n599 dvss.n49 57.2559
R422 dvss.n248 dvss.t171 57.1434
R423 dvss.n122 dvss.t40 57.1434
R424 dvss.n139 dvss.t182 57.1434
R425 dvss.n149 dvss.t195 57.1434
R426 dvss.n166 dvss.t127 57.1434
R427 dvss.n183 dvss.t159 57.1434
R428 dvss.n614 dvss.n42 54.0496
R429 dvss.n678 dvss.t15 52.8576
R430 dvss.n678 dvss.t136 51.4291
R431 dvss.n576 dvss.n575 45.2502
R432 dvss.n85 dvss.n39 44.978
R433 dvss.t134 dvss 42.227
R434 dvss.n216 dvss.n207 41.7862
R435 dvss.t134 dvss.n207 41.7862
R436 dvss.n215 dvss.n206 41.7862
R437 dvss.t134 dvss.n206 41.7862
R438 dvss.n541 dvss.n540 41.7862
R439 dvss.n542 dvss.n541 41.7862
R440 dvss.n102 dvss.n101 41.7862
R441 dvss.n101 dvss.n0 41.7862
R442 dvss.n554 dvss.n546 41.7862
R443 dvss.n546 dvss.n545 41.7862
R444 dvss.n552 dvss.n544 41.7862
R445 dvss.n544 dvss.n543 41.7862
R446 dvss.n231 dvss.n230 40.2432
R447 dvss.n677 dvss.n676 40.0735
R448 dvss.n236 dvss.t73 38.5719
R449 dvss.n236 dvss.t214 38.5719
R450 dvss.n110 dvss.t209 38.5719
R451 dvss.n110 dvss.t143 38.5719
R452 dvss.n127 dvss.t104 38.5719
R453 dvss.n127 dvss.t187 38.5719
R454 dvss.n163 dvss.t49 38.5719
R455 dvss.n163 dvss.t123 38.5719
R456 dvss.n180 dvss.t131 38.5719
R457 dvss.n180 dvss.t147 38.5719
R458 dvss.n198 dvss.t53 38.5719
R459 dvss.n198 dvss.t89 38.5719
R460 dvss.n634 dvss.n633 37.6894
R461 dvss.n584 dvss.n65 37.4862
R462 dvss.n611 dvss.n40 36.1883
R463 dvss.t13 dvss.t11 36.179
R464 dvss.n72 dvss.n71 36.179
R465 dvss.n6 dvss.t19 36.0005
R466 dvss.n565 dvss.n563 35.6976
R467 dvss.n537 dvss.n536 35.5421
R468 dvss.n670 dvss.n5 34.6358
R469 dvss.n671 dvss.n670 34.6358
R470 dvss.n672 dvss.n671 34.6358
R471 dvss.n300 dvss.n225 34.6358
R472 dvss.n293 dvss.n226 34.6358
R473 dvss.n276 dvss.n241 34.6358
R474 dvss.n277 dvss.n276 34.6358
R475 dvss.n278 dvss.n277 34.6358
R476 dvss.n278 dvss.n239 34.6358
R477 dvss.n282 dvss.n239 34.6358
R478 dvss.n264 dvss.n243 34.6358
R479 dvss.n268 dvss.n243 34.6358
R480 dvss.n269 dvss.n268 34.6358
R481 dvss.n272 dvss.n269 34.6358
R482 dvss.n251 dvss.n108 34.6358
R483 dvss.n255 dvss.n254 34.6358
R484 dvss.n257 dvss.n255 34.6358
R485 dvss.n261 dvss.n246 34.6358
R486 dvss.n262 dvss.n261 34.6358
R487 dvss.n505 dvss.n115 34.6358
R488 dvss.n506 dvss.n505 34.6358
R489 dvss.n507 dvss.n506 34.6358
R490 dvss.n507 dvss.n113 34.6358
R491 dvss.n511 dvss.n113 34.6358
R492 dvss.n493 dvss.n117 34.6358
R493 dvss.n497 dvss.n117 34.6358
R494 dvss.n498 dvss.n497 34.6358
R495 dvss.n501 dvss.n498 34.6358
R496 dvss.n480 dvss.n479 34.6358
R497 dvss.n484 dvss.n483 34.6358
R498 dvss.n486 dvss.n484 34.6358
R499 dvss.n490 dvss.n120 34.6358
R500 dvss.n491 dvss.n490 34.6358
R501 dvss.n465 dvss.n132 34.6358
R502 dvss.n466 dvss.n465 34.6358
R503 dvss.n467 dvss.n466 34.6358
R504 dvss.n467 dvss.n130 34.6358
R505 dvss.n471 dvss.n130 34.6358
R506 dvss.n453 dvss.n134 34.6358
R507 dvss.n457 dvss.n134 34.6358
R508 dvss.n458 dvss.n457 34.6358
R509 dvss.n461 dvss.n458 34.6358
R510 dvss.n440 dvss.n439 34.6358
R511 dvss.n444 dvss.n443 34.6358
R512 dvss.n446 dvss.n444 34.6358
R513 dvss.n450 dvss.n137 34.6358
R514 dvss.n451 dvss.n450 34.6358
R515 dvss.n433 dvss.n147 34.6358
R516 dvss.n429 dvss.n428 34.6358
R517 dvss.n428 dvss.n427 34.6358
R518 dvss.n424 dvss.n423 34.6358
R519 dvss.n423 dvss.n422 34.6358
R520 dvss.n419 dvss.n418 34.6358
R521 dvss.n418 dvss.n417 34.6358
R522 dvss.n417 dvss.n156 34.6358
R523 dvss.n413 dvss.n156 34.6358
R524 dvss.n411 dvss.n410 34.6358
R525 dvss.n410 dvss.n159 34.6358
R526 dvss.n406 dvss.n159 34.6358
R527 dvss.n406 dvss.n405 34.6358
R528 dvss.n405 dvss.n404 34.6358
R529 dvss.n394 dvss.n393 34.6358
R530 dvss.n391 dvss.n167 34.6358
R531 dvss.n387 dvss.n167 34.6358
R532 dvss.n385 dvss.n384 34.6358
R533 dvss.n384 dvss.n169 34.6358
R534 dvss.n380 dvss.n379 34.6358
R535 dvss.n379 dvss.n378 34.6358
R536 dvss.n378 dvss.n173 34.6358
R537 dvss.n374 dvss.n173 34.6358
R538 dvss.n372 dvss.n371 34.6358
R539 dvss.n371 dvss.n176 34.6358
R540 dvss.n367 dvss.n176 34.6358
R541 dvss.n367 dvss.n366 34.6358
R542 dvss.n366 dvss.n365 34.6358
R543 dvss.n355 dvss.n354 34.6358
R544 dvss.n352 dvss.n184 34.6358
R545 dvss.n348 dvss.n184 34.6358
R546 dvss.n346 dvss.n345 34.6358
R547 dvss.n345 dvss.n186 34.6358
R548 dvss.n341 dvss.n340 34.6358
R549 dvss.n340 dvss.n190 34.6358
R550 dvss.n336 dvss.n190 34.6358
R551 dvss.n336 dvss.n335 34.6358
R552 dvss.n333 dvss.n193 34.6358
R553 dvss.n329 dvss.n193 34.6358
R554 dvss.n329 dvss.n328 34.6358
R555 dvss.n328 dvss.n195 34.6358
R556 dvss.n322 dvss.n195 34.6358
R557 dvss.n314 dvss.n202 34.6358
R558 dvss.n309 dvss.n308 34.6358
R559 dvss.n23 dvss.t58 33.462
R560 dvss.n23 dvss.t212 33.462
R561 dvss.n74 dvss.t36 33.462
R562 dvss.n74 dvss.t175 33.462
R563 dvss.n2 dvss.t96 33.2313
R564 dvss.n24 dvss.n21 31.5123
R565 dvss.n254 dvss.n249 31.2476
R566 dvss.n483 dvss.n123 31.2476
R567 dvss.n443 dvss.n140 31.2476
R568 dvss.n429 dvss.n150 31.2476
R569 dvss.n392 dvss.n391 31.2476
R570 dvss.n353 dvss.n352 31.2476
R571 dvss.t7 dvss.t14 30.4092
R572 dvss dvss.n681 30.4092
R573 dvss.n616 dvss.n37 30.2484
R574 dvss.n284 dvss.n283 29.7417
R575 dvss.n513 dvss.n512 29.7417
R576 dvss.n473 dvss.n472 29.7417
R577 dvss.n400 dvss.n161 29.7417
R578 dvss.n361 dvss.n178 29.7417
R579 dvss.n321 dvss.n320 29.7417
R580 dvss.n80 dvss.n37 28.5338
R581 dvss.n538 dvss.n99 28.3255
R582 dvss.n527 dvss.n100 27.9866
R583 dvss.n256 dvss.n246 27.8593
R584 dvss.n485 dvss.n120 27.8593
R585 dvss.n445 dvss.n137 27.8593
R586 dvss.n424 dvss.n151 27.8593
R587 dvss.n386 dvss.n385 27.8593
R588 dvss.n347 dvss.n346 27.8593
R589 dvss.n676 dvss.n3 25.977
R590 dvss.n228 dvss.t0 25.6886
R591 dvss.n248 dvss.t149 25.4291
R592 dvss.n122 dvss.t77 25.4291
R593 dvss.n139 dvss.t177 25.4291
R594 dvss.n149 dvss.t18 25.4291
R595 dvss.n166 dvss.t86 25.4291
R596 dvss.n183 dvss.t4 25.4291
R597 dvss.n2 dvss.t97 24.9236
R598 dvss.n6 dvss.t8 24.9236
R599 dvss.n562 dvss.n561 24.3755
R600 dvss.n563 dvss.n562 24.3755
R601 dvss.n553 dvss.n92 24.3755
R602 dvss.n563 dvss.n92 24.3755
R603 dvss.n296 dvss.n225 23.7737
R604 dvss.n310 dvss.n309 23.7737
R605 dvss.n665 dvss.n7 23.7181
R606 dvss.n301 dvss.n300 23.7181
R607 dvss.n289 dvss.n226 23.7181
R608 dvss.n289 dvss.n288 23.7181
R609 dvss.n518 dvss.n108 23.7181
R610 dvss.n518 dvss.n517 23.7181
R611 dvss.n479 dvss.n478 23.7181
R612 dvss.n478 dvss.n477 23.7181
R613 dvss.n439 dvss.n438 23.7181
R614 dvss.n434 dvss.n433 23.7181
R615 dvss.n398 dvss.n164 23.7181
R616 dvss.n394 dvss.n164 23.7181
R617 dvss.n359 dvss.n181 23.7181
R618 dvss.n355 dvss.n181 23.7181
R619 dvss.n316 dvss.n315 23.7181
R620 dvss.n315 dvss.n314 23.7181
R621 dvss.n308 dvss.n305 23.7181
R622 dvss.n639 dvss.n26 23.7181
R623 dvss.n76 dvss.n73 23.7181
R624 dvss.n666 dvss.n5 22.9652
R625 dvss.n284 dvss.n237 22.9652
R626 dvss.n513 dvss.n111 22.9652
R627 dvss.n473 dvss.n128 22.9652
R628 dvss.n400 dvss.n399 22.9652
R629 dvss.n361 dvss.n360 22.9652
R630 dvss.n320 dvss.n199 22.9652
R631 dvss.n537 dvss.n533 22.1054
R632 dvss.n232 dvss.n107 21.7695
R633 dvss.n98 dvss.n97 21.753
R634 dvss.n666 dvss.n665 21.4593
R635 dvss.n288 dvss.n237 21.4593
R636 dvss.n517 dvss.n111 21.4593
R637 dvss.n477 dvss.n128 21.4593
R638 dvss.n399 dvss.n398 21.4593
R639 dvss.n360 dvss.n359 21.4593
R640 dvss.n316 dvss.n199 21.4593
R641 dvss.n680 dvss.n679 21.4265
R642 dvss.n552 dvss.t82 21.1687
R643 dvss.n554 dvss.t113 21.1687
R644 dvss.n220 dvss.t7 21.1543
R645 dvss.n295 dvss.n293 20.9718
R646 dvss.n205 dvss.n202 20.9718
R647 dvss.n576 dvss.n37 20.1009
R648 dvss.n617 dvss.n36 20.0732
R649 dvss.n528 dvss.n527 18.7867
R650 dvss.n559 dvss.n555 18.4515
R651 dvss.n558 dvss.n556 18.4515
R652 dvss.n549 dvss.n548 18.4515
R653 dvss.n550 dvss.n547 18.4515
R654 dvss.n672 dvss.n3 18.4476
R655 dvss.n263 dvss.n262 17.6946
R656 dvss.n492 dvss.n491 17.6946
R657 dvss.n452 dvss.n451 17.6946
R658 dvss.n422 dvss.n154 17.6946
R659 dvss.n172 dvss.n169 17.6946
R660 dvss.n189 dvss.n186 17.6946
R661 dvss.t178 dvss.n625 16.6567
R662 dvss dvss.n24 15.0593
R663 dvss dvss.n75 15.0593
R664 dvss.n283 dvss.n282 14.6829
R665 dvss.n512 dvss.n511 14.6829
R666 dvss.n472 dvss.n471 14.6829
R667 dvss.n404 dvss.n161 14.6829
R668 dvss.n365 dvss.n178 14.6829
R669 dvss.n322 dvss.n321 14.6829
R670 dvss.n594 dvss.n593 14.3573
R671 dvss.n570 dvss.n568 13.8612
R672 dvss.n71 dvss.t35 13.7828
R673 dvss.n99 dvss.n98 13.2836
R674 dvss.n606 dvss.n47 13.0628
R675 dvss.n610 dvss.n609 12.2414
R676 dvss.n97 dvss.n95 11.7338
R677 dvss.n581 dvss.n54 10.5081
R678 dvss.n597 dvss.n596 10.2484
R679 dvss.n592 dvss.n52 10.2179
R680 dvss.n656 dvss.n655 10.1264
R681 dvss.n649 dvss.n648 9.79535
R682 dvss.n582 dvss.n79 9.76662
R683 dvss.n596 dvss.n38 9.49353
R684 dvss.n80 dvss.n79 9.30109
R685 dvss.n306 dvss.n305 9.3005
R686 dvss.n324 dvss.n195 9.3005
R687 dvss.n323 dvss.n322 9.3005
R688 dvss.n321 dvss.n197 9.3005
R689 dvss.n320 dvss.n319 9.3005
R690 dvss.n318 dvss.n199 9.3005
R691 dvss.n317 dvss.n316 9.3005
R692 dvss.n315 dvss.n201 9.3005
R693 dvss.n314 dvss.n313 9.3005
R694 dvss.n312 dvss.n202 9.3005
R695 dvss.n311 dvss.n310 9.3005
R696 dvss.n309 dvss.n203 9.3005
R697 dvss.n308 dvss.n307 9.3005
R698 dvss.n434 dvss.n105 9.3005
R699 dvss.n433 dvss.n432 9.3005
R700 dvss.n431 dvss.n147 9.3005
R701 dvss.n430 dvss.n429 9.3005
R702 dvss.n428 dvss.n148 9.3005
R703 dvss.n427 dvss.n426 9.3005
R704 dvss.n425 dvss.n424 9.3005
R705 dvss.n423 dvss.n152 9.3005
R706 dvss.n422 dvss.n421 9.3005
R707 dvss.n420 dvss.n419 9.3005
R708 dvss.n418 dvss.n155 9.3005
R709 dvss.n417 dvss.n416 9.3005
R710 dvss.n415 dvss.n156 9.3005
R711 dvss.n414 dvss.n413 9.3005
R712 dvss.n411 dvss.n157 9.3005
R713 dvss.n410 dvss.n409 9.3005
R714 dvss.n408 dvss.n159 9.3005
R715 dvss.n407 dvss.n406 9.3005
R716 dvss.n405 dvss.n160 9.3005
R717 dvss.n404 dvss.n403 9.3005
R718 dvss.n402 dvss.n161 9.3005
R719 dvss.n401 dvss.n400 9.3005
R720 dvss.n399 dvss.n162 9.3005
R721 dvss.n398 dvss.n397 9.3005
R722 dvss.n396 dvss.n164 9.3005
R723 dvss.n395 dvss.n394 9.3005
R724 dvss.n393 dvss.n165 9.3005
R725 dvss.n391 dvss.n390 9.3005
R726 dvss.n389 dvss.n167 9.3005
R727 dvss.n388 dvss.n387 9.3005
R728 dvss.n385 dvss.n168 9.3005
R729 dvss.n384 dvss.n383 9.3005
R730 dvss.n382 dvss.n169 9.3005
R731 dvss.n381 dvss.n380 9.3005
R732 dvss.n379 dvss.n170 9.3005
R733 dvss.n378 dvss.n377 9.3005
R734 dvss.n376 dvss.n173 9.3005
R735 dvss.n375 dvss.n374 9.3005
R736 dvss.n372 dvss.n174 9.3005
R737 dvss.n371 dvss.n370 9.3005
R738 dvss.n369 dvss.n176 9.3005
R739 dvss.n368 dvss.n367 9.3005
R740 dvss.n366 dvss.n177 9.3005
R741 dvss.n365 dvss.n364 9.3005
R742 dvss.n363 dvss.n178 9.3005
R743 dvss.n362 dvss.n361 9.3005
R744 dvss.n360 dvss.n179 9.3005
R745 dvss.n359 dvss.n358 9.3005
R746 dvss.n357 dvss.n181 9.3005
R747 dvss.n356 dvss.n355 9.3005
R748 dvss.n354 dvss.n182 9.3005
R749 dvss.n352 dvss.n351 9.3005
R750 dvss.n350 dvss.n184 9.3005
R751 dvss.n349 dvss.n348 9.3005
R752 dvss.n346 dvss.n185 9.3005
R753 dvss.n345 dvss.n344 9.3005
R754 dvss.n343 dvss.n186 9.3005
R755 dvss.n342 dvss.n341 9.3005
R756 dvss.n340 dvss.n339 9.3005
R757 dvss.n338 dvss.n190 9.3005
R758 dvss.n337 dvss.n336 9.3005
R759 dvss.n335 dvss.n191 9.3005
R760 dvss.n333 dvss.n332 9.3005
R761 dvss.n331 dvss.n193 9.3005
R762 dvss.n330 dvss.n329 9.3005
R763 dvss.n328 dvss.n327 9.3005
R764 dvss.n438 dvss.n106 9.3005
R765 dvss.n439 dvss.n141 9.3005
R766 dvss.n441 dvss.n440 9.3005
R767 dvss.n443 dvss.n442 9.3005
R768 dvss.n444 dvss.n138 9.3005
R769 dvss.n447 dvss.n446 9.3005
R770 dvss.n448 dvss.n137 9.3005
R771 dvss.n450 dvss.n449 9.3005
R772 dvss.n451 dvss.n135 9.3005
R773 dvss.n454 dvss.n453 9.3005
R774 dvss.n455 dvss.n134 9.3005
R775 dvss.n457 dvss.n456 9.3005
R776 dvss.n458 dvss.n133 9.3005
R777 dvss.n462 dvss.n461 9.3005
R778 dvss.n463 dvss.n132 9.3005
R779 dvss.n465 dvss.n464 9.3005
R780 dvss.n466 dvss.n131 9.3005
R781 dvss.n468 dvss.n467 9.3005
R782 dvss.n469 dvss.n130 9.3005
R783 dvss.n471 dvss.n470 9.3005
R784 dvss.n472 dvss.n129 9.3005
R785 dvss.n474 dvss.n473 9.3005
R786 dvss.n475 dvss.n128 9.3005
R787 dvss.n477 dvss.n476 9.3005
R788 dvss.n478 dvss.n125 9.3005
R789 dvss.n479 dvss.n124 9.3005
R790 dvss.n481 dvss.n480 9.3005
R791 dvss.n483 dvss.n482 9.3005
R792 dvss.n484 dvss.n121 9.3005
R793 dvss.n487 dvss.n486 9.3005
R794 dvss.n488 dvss.n120 9.3005
R795 dvss.n490 dvss.n489 9.3005
R796 dvss.n491 dvss.n118 9.3005
R797 dvss.n494 dvss.n493 9.3005
R798 dvss.n495 dvss.n117 9.3005
R799 dvss.n497 dvss.n496 9.3005
R800 dvss.n498 dvss.n116 9.3005
R801 dvss.n502 dvss.n501 9.3005
R802 dvss.n503 dvss.n115 9.3005
R803 dvss.n505 dvss.n504 9.3005
R804 dvss.n506 dvss.n114 9.3005
R805 dvss.n508 dvss.n507 9.3005
R806 dvss.n509 dvss.n113 9.3005
R807 dvss.n511 dvss.n510 9.3005
R808 dvss.n512 dvss.n112 9.3005
R809 dvss.n514 dvss.n513 9.3005
R810 dvss.n515 dvss.n111 9.3005
R811 dvss.n517 dvss.n516 9.3005
R812 dvss.n519 dvss.n518 9.3005
R813 dvss.n250 dvss.n108 9.3005
R814 dvss.n252 dvss.n251 9.3005
R815 dvss.n254 dvss.n253 9.3005
R816 dvss.n255 dvss.n247 9.3005
R817 dvss.n258 dvss.n257 9.3005
R818 dvss.n259 dvss.n246 9.3005
R819 dvss.n261 dvss.n260 9.3005
R820 dvss.n262 dvss.n244 9.3005
R821 dvss.n265 dvss.n264 9.3005
R822 dvss.n266 dvss.n243 9.3005
R823 dvss.n268 dvss.n267 9.3005
R824 dvss.n269 dvss.n242 9.3005
R825 dvss.n273 dvss.n272 9.3005
R826 dvss.n274 dvss.n241 9.3005
R827 dvss.n276 dvss.n275 9.3005
R828 dvss.n277 dvss.n240 9.3005
R829 dvss.n279 dvss.n278 9.3005
R830 dvss.n280 dvss.n239 9.3005
R831 dvss.n282 dvss.n281 9.3005
R832 dvss.n283 dvss.n238 9.3005
R833 dvss.n285 dvss.n284 9.3005
R834 dvss.n286 dvss.n237 9.3005
R835 dvss.n288 dvss.n287 9.3005
R836 dvss.n290 dvss.n289 9.3005
R837 dvss.n291 dvss.n226 9.3005
R838 dvss.n293 dvss.n292 9.3005
R839 dvss.n297 dvss.n296 9.3005
R840 dvss.n298 dvss.n225 9.3005
R841 dvss.n300 dvss.n299 9.3005
R842 dvss.n301 dvss.n224 9.3005
R843 dvss.n662 dvss.n7 9.3005
R844 dvss.n667 dvss.n666 9.3005
R845 dvss.n673 dvss.n672 9.3005
R846 dvss.n671 dvss.n4 9.3005
R847 dvss.n670 dvss.n669 9.3005
R848 dvss.n668 dvss.n5 9.3005
R849 dvss.n665 dvss.n664 9.3005
R850 dvss.n674 dvss.n3 9.3005
R851 dvss.n676 dvss.n675 9.3005
R852 dvss.n640 dvss.n639 9.3005
R853 dvss.n24 dvss.n20 9.3005
R854 dvss.n26 dvss.n25 9.3005
R855 dvss.n644 dvss.n13 9.3005
R856 dvss.n77 dvss.n76 9.3005
R857 dvss.n73 dvss.n67 9.3005
R858 dvss.n635 dvss.n634 8.88939
R859 dvss.n68 dvss.n65 8.77764
R860 dvss.n528 dvss.n103 8.43597
R861 dvss.n271 dvss.n241 7.90638
R862 dvss.n500 dvss.n115 7.90638
R863 dvss.n460 dvss.n132 7.90638
R864 dvss.n412 dvss.n411 7.90638
R865 dvss.n373 dvss.n372 7.90638
R866 dvss.n334 dvss.n333 7.90638
R867 dvss.n620 dvss.n619 7.40556
R868 dvss.n621 dvss.n620 7.40556
R869 dvss.n603 dvss.n602 7.17831
R870 dvss.n75 dvss.n66 7.17078
R871 dvss.n26 dvss 7.15344
R872 dvss.n76 dvss 7.15344
R873 dvss.n569 dvss.n50 7.1196
R874 dvss.n257 dvss.n256 6.77697
R875 dvss.n486 dvss.n485 6.77697
R876 dvss.n446 dvss.n445 6.77697
R877 dvss.n427 dvss.n151 6.77697
R878 dvss.n387 dvss.n386 6.77697
R879 dvss.n348 dvss.n347 6.77697
R880 dvss.n538 dvss.n537 6.7205
R881 dvss.n216 dvss.n196 6.7005
R882 dvss.n679 dvss.n677 6.56103
R883 dvss.n525 dvss.n104 6.53261
R884 dvss.n230 dvss.n82 6.36591
R885 dvss.n602 dvss.n601 5.73579
R886 dvss.n621 dvss.n34 5.34031
R887 dvss.n598 dvss.n47 5.31835
R888 dvss.n565 dvss.n564 5.28896
R889 dvss.n572 dvss.n86 5.28896
R890 dvss.n609 dvss.n47 4.48642
R891 dvss.n555 dvss.t80 4.3505
R892 dvss.n555 dvss.t60 4.3505
R893 dvss.n556 dvss.t151 4.3505
R894 dvss.n556 dvss.t109 4.3505
R895 dvss.n548 dvss.t68 4.3505
R896 dvss.n548 dvss.t64 4.3505
R897 dvss.n547 dvss.t62 4.3505
R898 dvss.n547 dvss.t115 4.3505
R899 dvss.n529 dvss.n528 4.00961
R900 dvss.n577 dvss.n576 3.89404
R901 dvss.n583 dvss.n582 3.84425
R902 dvss.n602 dvss.n17 3.58941
R903 dvss.n579 dvss.n36 3.56414
R904 dvss.n584 dvss.n583 3.54405
R905 dvss.n251 dvss.n249 3.38874
R906 dvss.n480 dvss.n123 3.38874
R907 dvss.n440 dvss.n140 3.38874
R908 dvss.n150 dvss.n147 3.38874
R909 dvss.n393 dvss.n392 3.38874
R910 dvss.n354 dvss.n353 3.38874
R911 dvss.n666 dvss 3.29747
R912 dvss.n680 dvss.n1 3.21038
R913 dvss.n539 dvss.n96 3.01827
R914 dvss.n650 dvss.n649 2.88227
R915 dvss.n567 dvss.n566 2.75993
R916 dvss.n566 dvss.n565 2.75993
R917 dvss.n568 dvss.n87 2.75993
R918 dvss.n564 dvss.n87 2.75993
R919 dvss.n563 dvss.n91 2.64473
R920 dvss.n264 dvss.n263 2.63579
R921 dvss.n493 dvss.n492 2.63579
R922 dvss.n453 dvss.n452 2.63579
R923 dvss.n419 dvss.n154 2.63579
R924 dvss.n380 dvss.n172 2.63579
R925 dvss.n341 dvss.n189 2.63579
R926 dvss.n632 dvss.n22 2.47305
R927 dvss.n67 dvss.n65 2.41042
R928 dvss.n634 dvss.n22 2.33976
R929 dvss.n530 dvss.n96 2.3185
R930 dvss.n575 dvss.n82 1.98969
R931 dvss.n677 dvss.n1 1.93239
R932 dvss.n41 dvss.n36 1.92484
R933 dvss.n272 dvss.n271 1.88285
R934 dvss.n501 dvss.n500 1.88285
R935 dvss.n461 dvss.n460 1.88285
R936 dvss.n413 dvss.n412 1.88285
R937 dvss.n374 dvss.n373 1.88285
R938 dvss.n335 dvss.n334 1.88285
R939 dvss.n103 dvss.n102 1.85983
R940 dvss.n597 dvss.n46 1.80934
R941 dvss.n560 dvss.n559 1.57196
R942 dvss.n551 dvss.n550 1.57139
R943 dvss.n208 dvss.n194 1.5505
R944 dvss.n618 dvss.n18 1.48151
R945 dvss.n34 dvss.n18 1.48151
R946 dvss.n585 dvss.n584 1.46336
R947 dvss.n654 dvss.n14 1.32907
R948 dvss.n591 dvss.n590 1.32907
R949 dvss.n530 dvss.n529 1.21052
R950 dvss.n326 dvss.n196 1.11858
R951 dvss.n566 dvss.n87 1.10724
R952 dvss.n571 dvss.n88 1.10724
R953 dvss.n579 dvss.n37 1.01868
R954 dvss.n567 dvss.n89 0.899376
R955 dvss.n618 dvss.n19 0.804872
R956 dvss.n593 dvss.n38 0.778315
R957 dvss.n575 dvss.n574 0.774309
R958 dvss.n574 dvss.n573 0.774309
R959 dvss.n214 dvss.n208 0.649775
R960 dvss.n296 dvss.n295 0.630008
R961 dvss.n310 dvss.n205 0.630008
R962 dvss.n536 dvss.n89 0.629714
R963 dvss.n620 dvss.n18 0.538751
R964 dvss.n610 dvss.n46 0.533285
R965 dvss.n233 dvss.n232 0.519117
R966 dvss.n234 dvss.n233 0.519117
R967 dvss.n535 dvss.n533 0.482579
R968 dvss.t202 dvss.n657 0.474702
R969 dvss.n657 dvss.n656 0.447064
R970 dvss.n529 dvss.n100 0.443357
R971 dvss.n531 dvss.n530 0.443357
R972 dvss.n227 dvss.n104 0.428132
R973 dvss.n227 dvss.n146 0.428132
R974 dvss.n522 dvss.n104 0.411509
R975 dvss.n616 dvss.n38 0.362946
R976 dvss.n526 dvss.n90 0.355045
R977 dvss.n211 dvss.n90 0.355045
R978 dvss.n604 dvss.n601 0.336965
R979 dvss.n600 dvss.n17 0.328522
R980 dvss.n103 dvss 0.326572
R981 dvss.n605 dvss.n600 0.326101
R982 dvss.n592 dvss.n11 0.313726
R983 dvss.n557 dvss.n82 0.277008
R984 dvss.n662 dvss.n661 0.274194
R985 dvss.n534 dvss.n51 0.271039
R986 dvss.n583 dvss.n78 0.262597
R987 dvss.n611 dvss.n610 0.2605
R988 dvss.n612 dvss.n611 0.2605
R989 dvss.n539 dvss.n538 0.248336
R990 dvss.n81 dvss.n80 0.218682
R991 dvss.n608 dvss.n48 0.210906
R992 dvss.n642 dvss.n641 0.206439
R993 dvss.n595 dvss.n48 0.202526
R994 dvss.n187 dvss.t205 0.189075
R995 dvss.n525 dvss.n524 0.181217
R996 dvss.n633 dvss.n632 0.178278
R997 dvss.n582 dvss.n581 0.170143
R998 dvss.n607 dvss.n606 0.166164
R999 dvss.n601 dvss.n600 0.155797
R1000 dvss dvss.n660 0.150986
R1001 dvss.n51 dvss.n50 0.145813
R1002 dvss.n325 dvss 0.142307
R1003 dvss.n222 dvss 0.140841
R1004 dvss.n660 dvss.n659 0.13579
R1005 dvss.n607 dvss.n599 0.130165
R1006 dvss.n223 dvss 0.127978
R1007 dvss.n223 dvss.n222 0.123227
R1008 dvss.n532 dvss.n531 0.122311
R1009 dvss.n523 dvss.n106 0.121873
R1010 dvss.n324 dvss.n323 0.120292
R1011 dvss.n323 dvss.n197 0.120292
R1012 dvss.n319 dvss.n197 0.120292
R1013 dvss.n319 dvss.n318 0.120292
R1014 dvss.n318 dvss.n317 0.120292
R1015 dvss.n313 dvss.n312 0.120292
R1016 dvss.n311 dvss.n203 0.120292
R1017 dvss.n307 dvss.n203 0.120292
R1018 dvss.n668 dvss.n667 0.120292
R1019 dvss.n669 dvss.n668 0.120292
R1020 dvss.n669 dvss.n4 0.120292
R1021 dvss.n673 dvss.n4 0.120292
R1022 dvss.n674 dvss.n673 0.120292
R1023 dvss.n675 dvss.n674 0.120292
R1024 dvss.n144 dvss.n143 0.104964
R1025 dvss.n312 dvss 0.104667
R1026 dvss.n594 dvss.n51 0.103194
R1027 dvss.n326 dvss 0.0999624
R1028 dvss.n667 dvss 0.0968542
R1029 dvss.n643 dvss 0.0941255
R1030 dvss.n606 dvss.n605 0.0879466
R1031 dvss.n648 dvss.n647 0.0850455
R1032 dvss.n66 dvss 0.080434
R1033 dvss.n221 dvss 0.0781256
R1034 dvss.n77 dvss.n66 0.0777204
R1035 dvss.n645 dvss 0.0770968
R1036 dvss.n578 dvss.n577 0.0749
R1037 dvss.n524 dvss.n523 0.0737044
R1038 dvss.n568 dvss.n567 0.0724101
R1039 dvss.n570 dvss.n569 0.0724101
R1040 dvss.t204 dvss.t203 0.070611
R1041 dvss.n560 dvss.n554 0.0678684
R1042 dvss.n658 dvss.t202 0.0675999
R1043 dvss.n552 dvss.n551 0.0671667
R1044 dvss.n595 dvss.n594 0.06684
R1045 dvss.n222 dvss.n221 0.0638562
R1046 dvss.n557 dvss 0.0633141
R1047 dvss.n581 dvss.n580 0.0614929
R1048 dvss.n659 dvss.t205 0.060491
R1049 dvss.n201 dvss 0.0603958
R1050 dvss.n313 dvss 0.0603958
R1051 dvss dvss.n306 0.0603958
R1052 dvss.n664 dvss 0.0603958
R1053 dvss.n657 dvss.n11 0.0595861
R1054 dvss.n221 dvss.n8 0.0586797
R1055 dvss.n98 dvss.n9 0.0559625
R1056 dvss.n143 dvss.n49 0.0535781
R1057 dvss.n608 dvss.n607 0.0533794
R1058 dvss.n1 dvss 0.0525833
R1059 dvss.n14 dvss 0.0515042
R1060 dvss.n25 dvss.n20 0.0480207
R1061 dvss.n643 dvss.n642 0.0476863
R1062 dvss.n524 dvss.n105 0.0461989
R1063 dvss.n550 dvss.n549 0.0457733
R1064 dvss.n325 dvss.n324 0.0447708
R1065 dvss.n658 dvss.n10 0.0405094
R1066 dvss.n642 dvss.n21 0.0402727
R1067 dvss.n593 dvss.n592 0.0393298
R1068 dvss.n531 dvss.n100 0.0374705
R1069 dvss.n619 dvss.n618 0.0354727
R1070 dvss dvss.n591 0.0347199
R1071 dvss.n559 dvss 0.0346686
R1072 dvss.n580 dvss.n579 0.0341957
R1073 dvss dvss.n201 0.0330521
R1074 dvss.n306 dvss 0.0330521
R1075 dvss.n19 dvss.n11 0.0323493
R1076 dvss.n656 dvss 0.0323446
R1077 dvss.n534 dvss.n89 0.0321327
R1078 dvss.n48 dvss.n46 0.0315
R1079 dvss.n581 dvss.n578 0.0306418
R1080 dvss.n532 dvss.n99 0.0284126
R1081 dvss dvss.n662 0.0271393
R1082 dvss.n592 dvss 0.0255
R1083 dvss.n641 dvss.n22 0.0247851
R1084 dvss.n641 dvss.n640 0.0242603
R1085 dvss.n25 dvss 0.0242603
R1086 dvss.n21 dvss 0.0242603
R1087 dvss.n536 dvss.n535 0.0239848
R1088 dvss.n664 dvss 0.0239375
R1089 dvss.n647 dvss.n645 0.0230951
R1090 dvss.n549 dvss.n10 0.0228519
R1091 dvss.n317 dvss 0.0226354
R1092 dvss.n307 dvss 0.0226354
R1093 dvss.n78 dvss 0.0215598
R1094 dvss.n8 dvss 0.0206613
R1095 dvss.n231 dvss.n9 0.0206307
R1096 dvss.n663 dvss 0.0199672
R1097 dvss.n523 dvss.n522 0.0192879
R1098 dvss.n521 dvss.n520 0.0189524
R1099 dvss.n596 dvss.n595 0.0189524
R1100 dvss.n558 dvss.n557 0.0184385
R1101 dvss.n67 dvss 0.0174837
R1102 dvss.n578 dvss.n79 0.0174213
R1103 dvss.n609 dvss.n608 0.0166458
R1104 dvss dvss.n311 0.016125
R1105 dvss.n432 dvss.n431 0.015957
R1106 dvss.n431 dvss.n430 0.015957
R1107 dvss.n430 dvss.n148 0.015957
R1108 dvss.n426 dvss.n148 0.015957
R1109 dvss.n426 dvss.n425 0.015957
R1110 dvss.n425 dvss.n152 0.015957
R1111 dvss.n421 dvss.n152 0.015957
R1112 dvss.n421 dvss.n420 0.015957
R1113 dvss.n420 dvss.n155 0.015957
R1114 dvss.n416 dvss.n155 0.015957
R1115 dvss.n416 dvss.n415 0.015957
R1116 dvss.n415 dvss.n414 0.015957
R1117 dvss.n414 dvss.n157 0.015957
R1118 dvss.n409 dvss.n157 0.015957
R1119 dvss.n409 dvss.n408 0.015957
R1120 dvss.n408 dvss.n407 0.015957
R1121 dvss.n407 dvss.n160 0.015957
R1122 dvss.n403 dvss.n160 0.015957
R1123 dvss.n403 dvss.n402 0.015957
R1124 dvss.n402 dvss.n401 0.015957
R1125 dvss.n401 dvss.n162 0.015957
R1126 dvss.n397 dvss.n162 0.015957
R1127 dvss.n395 dvss.n165 0.015957
R1128 dvss.n390 dvss.n165 0.015957
R1129 dvss.n390 dvss.n389 0.015957
R1130 dvss.n389 dvss.n388 0.015957
R1131 dvss.n388 dvss.n168 0.015957
R1132 dvss.n383 dvss.n168 0.015957
R1133 dvss.n383 dvss.n382 0.015957
R1134 dvss.n382 dvss.n381 0.015957
R1135 dvss.n381 dvss.n170 0.015957
R1136 dvss.n377 dvss.n170 0.015957
R1137 dvss.n377 dvss.n376 0.015957
R1138 dvss.n376 dvss.n375 0.015957
R1139 dvss.n375 dvss.n174 0.015957
R1140 dvss.n370 dvss.n174 0.015957
R1141 dvss.n370 dvss.n369 0.015957
R1142 dvss.n369 dvss.n368 0.015957
R1143 dvss.n368 dvss.n177 0.015957
R1144 dvss.n364 dvss.n177 0.015957
R1145 dvss.n364 dvss.n363 0.015957
R1146 dvss.n363 dvss.n362 0.015957
R1147 dvss.n362 dvss.n179 0.015957
R1148 dvss.n358 dvss.n179 0.015957
R1149 dvss.n356 dvss.n182 0.015957
R1150 dvss.n351 dvss.n182 0.015957
R1151 dvss.n351 dvss.n350 0.015957
R1152 dvss.n350 dvss.n349 0.015957
R1153 dvss.n349 dvss.n185 0.015957
R1154 dvss.n344 dvss.n185 0.015957
R1155 dvss.n344 dvss.n343 0.015957
R1156 dvss.n343 dvss.n342 0.015957
R1157 dvss.n339 dvss.n338 0.015957
R1158 dvss.n338 dvss.n337 0.015957
R1159 dvss.n337 dvss.n191 0.015957
R1160 dvss.n332 dvss.n191 0.015957
R1161 dvss.n332 dvss.n331 0.015957
R1162 dvss.n331 dvss.n330 0.015957
R1163 dvss.n326 dvss.n325 0.0141555
R1164 dvss.n644 dvss.n643 0.0140978
R1165 dvss.n640 dvss 0.0139298
R1166 dvss.n441 dvss.n141 0.0125293
R1167 dvss.n442 dvss.n441 0.0125293
R1168 dvss.n442 dvss.n138 0.0125293
R1169 dvss.n447 dvss.n138 0.0125293
R1170 dvss.n448 dvss.n447 0.0125293
R1171 dvss.n449 dvss.n448 0.0125293
R1172 dvss.n449 dvss.n135 0.0125293
R1173 dvss.n454 dvss.n135 0.0125293
R1174 dvss.n455 dvss.n454 0.0125293
R1175 dvss.n456 dvss.n455 0.0125293
R1176 dvss.n456 dvss.n133 0.0125293
R1177 dvss.n462 dvss.n133 0.0125293
R1178 dvss.n463 dvss.n462 0.0125293
R1179 dvss.n464 dvss.n463 0.0125293
R1180 dvss.n464 dvss.n131 0.0125293
R1181 dvss.n468 dvss.n131 0.0125293
R1182 dvss.n469 dvss.n468 0.0125293
R1183 dvss.n470 dvss.n469 0.0125293
R1184 dvss.n470 dvss.n129 0.0125293
R1185 dvss.n474 dvss.n129 0.0125293
R1186 dvss.n475 dvss.n474 0.0125293
R1187 dvss.n476 dvss.n475 0.0125293
R1188 dvss.n481 dvss.n124 0.0125293
R1189 dvss.n482 dvss.n481 0.0125293
R1190 dvss.n482 dvss.n121 0.0125293
R1191 dvss.n487 dvss.n121 0.0125293
R1192 dvss.n488 dvss.n487 0.0125293
R1193 dvss.n489 dvss.n488 0.0125293
R1194 dvss.n489 dvss.n118 0.0125293
R1195 dvss.n494 dvss.n118 0.0125293
R1196 dvss.n495 dvss.n494 0.0125293
R1197 dvss.n496 dvss.n495 0.0125293
R1198 dvss.n496 dvss.n116 0.0125293
R1199 dvss.n502 dvss.n116 0.0125293
R1200 dvss.n503 dvss.n502 0.0125293
R1201 dvss.n504 dvss.n503 0.0125293
R1202 dvss.n504 dvss.n114 0.0125293
R1203 dvss.n508 dvss.n114 0.0125293
R1204 dvss.n509 dvss.n508 0.0125293
R1205 dvss.n510 dvss.n509 0.0125293
R1206 dvss.n510 dvss.n112 0.0125293
R1207 dvss.n514 dvss.n112 0.0125293
R1208 dvss.n515 dvss.n514 0.0125293
R1209 dvss.n516 dvss.n515 0.0125293
R1210 dvss.n252 dvss.n250 0.0125293
R1211 dvss.n253 dvss.n252 0.0125293
R1212 dvss.n253 dvss.n247 0.0125293
R1213 dvss.n258 dvss.n247 0.0125293
R1214 dvss.n259 dvss.n258 0.0125293
R1215 dvss.n260 dvss.n259 0.0125293
R1216 dvss.n260 dvss.n244 0.0125293
R1217 dvss.n265 dvss.n244 0.0125293
R1218 dvss.n266 dvss.n265 0.0125293
R1219 dvss.n267 dvss.n266 0.0125293
R1220 dvss.n267 dvss.n242 0.0125293
R1221 dvss.n273 dvss.n242 0.0125293
R1222 dvss.n274 dvss.n273 0.0125293
R1223 dvss.n275 dvss.n274 0.0125293
R1224 dvss.n275 dvss.n240 0.0125293
R1225 dvss.n279 dvss.n240 0.0125293
R1226 dvss.n280 dvss.n279 0.0125293
R1227 dvss.n281 dvss.n280 0.0125293
R1228 dvss.n281 dvss.n238 0.0125293
R1229 dvss.n285 dvss.n238 0.0125293
R1230 dvss.n286 dvss.n285 0.0125293
R1231 dvss.n287 dvss.n286 0.0125293
R1232 dvss.n292 dvss.n291 0.0125293
R1233 dvss.n298 dvss.n297 0.0125293
R1234 dvss.n299 dvss.n298 0.0125293
R1235 dvss.n339 dvss.n187 0.0122608
R1236 dvss dvss.n558 0.0110353
R1237 dvss.n292 dvss 0.0109603
R1238 dvss.n78 dvss.n77 0.0106902
R1239 dvss.n659 dvss.t204 0.0106199
R1240 dvss.n580 dvss.n53 0.0101631
R1241 dvss.n327 dvss.n194 0.0099086
R1242 dvss.n661 dvss.n8 0.00990439
R1243 dvss.n660 dvss.n9 0.00933152
R1244 dvss.n675 dvss.n1 0.0083125
R1245 dvss.n642 dvss.n20 0.00824793
R1246 dvss.n535 dvss.n534 0.00822968
R1247 dvss.n432 dvss 0.00822849
R1248 dvss dvss.n396 0.00822849
R1249 dvss dvss.n395 0.00822849
R1250 dvss dvss.n357 0.00822849
R1251 dvss dvss.n356 0.00822849
R1252 dvss.n647 dvss.n646 0.00789958
R1253 dvss.n330 dvss.n194 0.00654839
R1254 dvss.n141 dvss 0.00651464
R1255 dvss dvss.n125 0.00651464
R1256 dvss dvss.n124 0.00651464
R1257 dvss.n250 dvss 0.00651464
R1258 dvss.n290 dvss 0.00651464
R1259 dvss.n291 dvss 0.00651464
R1260 dvss dvss.n224 0.00651464
R1261 dvss.n520 dvss.n519 0.00573013
R1262 dvss dvss.n1 0.00570833
R1263 dvss.n557 dvss.n10 0.00519818
R1264 dvss.n661 dvss 0.00481034
R1265 dvss dvss.n105 0.00470027
R1266 dvss.n396 dvss 0.00470027
R1267 dvss.n357 dvss 0.00470027
R1268 dvss.n342 dvss.n187 0.00419624
R1269 dvss.n645 dvss.n644 0.00411776
R1270 dvss dvss.n106 0.00376883
R1271 dvss.n125 dvss 0.00376883
R1272 dvss.n519 dvss 0.00376883
R1273 dvss dvss.n290 0.00376883
R1274 dvss.n224 dvss 0.00376883
R1275 dvss.t203 dvss.n658 0.00351108
R1276 dvss.n397 dvss 0.00335618
R1277 dvss.n358 dvss 0.00335618
R1278 dvss.n476 dvss 0.0027228
R1279 dvss.n516 dvss 0.0027228
R1280 dvss.n287 dvss 0.0027228
R1281 dvss.n299 dvss 0.0027228
R1282 dvss.n297 dvss 0.00206904
R1283 dvss dvss.n663 0.00180208
R1284 dvss.n533 dvss.n532 0.00156293
R1285 dvss.n663 dvss 0.00152459
R1286 dvss.n327 dvss.n326 0.00150806
R1287 dvss.n520 dvss 0.00128452
R1288 dvss dvss.n223 0.00077533
R1289 dvss.n646 dvss.n14 0.000632135
R1290 dvss.n591 dvss.n53 0.000588652
R1291 dvdd.n295 dvdd.n286 5128.23
R1292 dvdd.n295 dvdd.n287 5128.23
R1293 dvdd.n293 dvdd.n287 5128.23
R1294 dvdd.n293 dvdd.n286 5128.23
R1295 dvdd.n42 dvdd.n5 1736.47
R1296 dvdd.n45 dvdd.n4 1736.47
R1297 dvdd.n30 dvdd.n27 1736.47
R1298 dvdd.n33 dvdd.n29 1736.47
R1299 dvdd.n255 dvdd.t146 838.817
R1300 dvdd.n69 dvdd.t169 806.511
R1301 dvdd.n69 dvdd.t101 806.511
R1302 dvdd.n90 dvdd.t7 806.511
R1303 dvdd.n90 dvdd.t142 806.511
R1304 dvdd.n111 dvdd.t122 806.511
R1305 dvdd.n111 dvdd.t74 806.511
R1306 dvdd.n292 dvdd.n284 787.447
R1307 dvdd.n292 dvdd.n285 786.827
R1308 dvdd.n56 dvdd.t32 668.683
R1309 dvdd.n56 dvdd.t153 668.683
R1310 dvdd.n227 dvdd.t124 667.778
R1311 dvdd.n227 dvdd.t128 667.778
R1312 dvdd.n189 dvdd.t164 667.778
R1313 dvdd.n189 dvdd.t107 667.778
R1314 dvdd.n151 dvdd.t76 667.778
R1315 dvdd.n151 dvdd.t98 667.778
R1316 dvdd.n296 dvdd.n284 604.574
R1317 dvdd.n73 dvdd.n71 604.457
R1318 dvdd.n73 dvdd.n72 604.457
R1319 dvdd.n94 dvdd.n92 604.457
R1320 dvdd.n94 dvdd.n93 604.457
R1321 dvdd.n115 dvdd.n113 604.457
R1322 dvdd.n115 dvdd.n114 604.457
R1323 dvdd.n232 dvdd.n61 604.394
R1324 dvdd.n232 dvdd.n62 604.394
R1325 dvdd.n194 dvdd.n82 604.394
R1326 dvdd.n194 dvdd.n83 604.394
R1327 dvdd.n156 dvdd.n103 604.394
R1328 dvdd.n156 dvdd.n104 604.394
R1329 dvdd.n220 dvdd.n67 601.679
R1330 dvdd.n220 dvdd.n68 601.679
R1331 dvdd.n182 dvdd.n88 601.679
R1332 dvdd.n182 dvdd.n89 601.679
R1333 dvdd.n144 dvdd.n109 601.679
R1334 dvdd.n144 dvdd.n110 601.679
R1335 dvdd.n260 dvdd.n259 585
R1336 dvdd.t35 dvdd.t145 556.386
R1337 dvdd.n246 dvdd 538.664
R1338 dvdd.n18 dvdd 535.705
R1339 dvdd.n11 dvdd 535.705
R1340 dvdd.t93 dvdd 473.521
R1341 dvdd.t75 dvdd.t62 448.146
R1342 dvdd.t106 dvdd.t113 448.146
R1343 dvdd.t123 dvdd.t70 448.146
R1344 dvdd.n296 dvdd.n285 423.062
R1345 dvdd.t161 dvdd.t157 367.579
R1346 dvdd.t58 dvdd.t56 367.579
R1347 dvdd.t132 dvdd.t134 367.579
R1348 dvdd.n274 dvdd.t33 360.005
R1349 dvdd.t73 dvdd.t46 330.654
R1350 dvdd.t6 dvdd.t38 330.654
R1351 dvdd.t100 dvdd.t42 330.654
R1352 dvdd.n43 dvdd.n4 314.781
R1353 dvdd.n44 dvdd.n5 314.781
R1354 dvdd.n31 dvdd.n29 314.781
R1355 dvdd.n32 dvdd.n27 314.781
R1356 dvdd.n23 dvdd.n17 312.053
R1357 dvdd.n9 dvdd.n8 312.051
R1358 dvdd.n266 dvdd.n256 312.051
R1359 dvdd.t117 dvdd.t119 304.829
R1360 dvdd.t145 dvdd.t95 284.113
R1361 dvdd.t157 dvdd.t148 275.265
R1362 dvdd.t56 dvdd.t60 275.265
R1363 dvdd.t134 dvdd.t2 275.265
R1364 dvdd.t95 dvdd.t93 275.235
R1365 dvdd.n271 dvdd.t138 261.837
R1366 dvdd.t115 dvdd.t154 260.437
R1367 dvdd.t140 dvdd.t172 260.437
R1368 dvdd.n207 dvdd.n76 259.707
R1369 dvdd.n207 dvdd.n75 259.707
R1370 dvdd.n169 dvdd.n97 259.707
R1371 dvdd.n169 dvdd.n96 259.707
R1372 dvdd.n131 dvdd.n118 259.707
R1373 dvdd.n131 dvdd.n117 259.707
R1374 dvdd.t138 dvdd.t77 258.481
R1375 dvdd.n273 dvdd.t83 253.446
R1376 dvdd.n272 dvdd.t4 253.446
R1377 dvdd.t30 dvdd.t90 248.599
R1378 dvdd.t90 dvdd.t35 248.599
R1379 dvdd.n201 dvdd.n80 242.607
R1380 dvdd.n163 dvdd.n101 242.607
R1381 dvdd.n125 dvdd.n123 242.607
R1382 dvdd.n201 dvdd.n79 242.607
R1383 dvdd.n163 dvdd.n100 242.607
R1384 dvdd.n125 dvdd.n122 242.607
R1385 dvdd.t81 dvdd.t64 234.982
R1386 dvdd.t66 dvdd.t111 234.982
R1387 dvdd.t50 dvdd.t68 234.982
R1388 dvdd dvdd.n270 232.445
R1389 dvdd.n0 dvdd.t13 228.215
R1390 dvdd.n0 dvdd.t49 228.215
R1391 dvdd.n239 dvdd.n59 215.123
R1392 dvdd.n239 dvdd.n238 215.123
R1393 dvdd.t119 dvdd.t80 213.084
R1394 dvdd.n41 dvdd.n3 185.225
R1395 dvdd.n46 dvdd.n3 185.225
R1396 dvdd.n34 dvdd.n28 185.225
R1397 dvdd.n28 dvdd.n26 185.225
R1398 dvdd.t36 dvdd.t159 181.273
R1399 dvdd.t40 dvdd.t54 181.273
R1400 dvdd.t44 dvdd.t136 181.273
R1401 dvdd.t65 dvdd.t73 166.167
R1402 dvdd.t64 dvdd.t91 166.167
R1403 dvdd.t112 dvdd.t6 166.167
R1404 dvdd.t111 dvdd.t52 166.167
R1405 dvdd.t69 dvdd.t100 166.167
R1406 dvdd.t68 dvdd.t1 166.167
R1407 dvdd.t33 dvdd.t161 162.81
R1408 dvdd.t46 dvdd.t81 162.81
R1409 dvdd.t83 dvdd.t58 162.81
R1410 dvdd.t38 dvdd.t66 162.81
R1411 dvdd.t4 dvdd.t132 162.81
R1412 dvdd.t42 dvdd.t50 162.81
R1413 dvdd.t14 dvdd.n293 161.316
R1414 dvdd.n295 dvdd.t28 161.316
R1415 dvdd.t91 dvdd.t75 154.417
R1416 dvdd.t52 dvdd.t106 154.417
R1417 dvdd.t1 dvdd.t123 154.417
R1418 dvdd.t77 dvdd.t31 147.703
R1419 dvdd.n75 dvdd.t87 147.111
R1420 dvdd.n76 dvdd.t3 147.111
R1421 dvdd.n96 dvdd.t61 147.111
R1422 dvdd.n97 dvdd.t85 147.111
R1423 dvdd.n117 dvdd.t149 147.111
R1424 dvdd.n118 dvdd.t163 147.111
R1425 dvdd.t92 dvdd.t65 144.346
R1426 dvdd.t53 dvdd.t112 144.346
R1427 dvdd.t0 dvdd.t69 144.346
R1428 dvdd.t148 dvdd.t36 140.989
R1429 dvdd.t159 dvdd.t92 140.989
R1430 dvdd.t62 dvdd.t104 140.989
R1431 dvdd.t60 dvdd.t40 140.989
R1432 dvdd.t54 dvdd.t53 140.989
R1433 dvdd.t113 dvdd.t125 140.989
R1434 dvdd.t2 dvdd.t44 140.989
R1435 dvdd.t136 dvdd.t0 140.989
R1436 dvdd.t70 dvdd.t88 140.989
R1437 dvdd.t31 dvdd 132.597
R1438 dvdd dvdd.n273 125.883
R1439 dvdd dvdd.n272 125.883
R1440 dvdd dvdd.n271 125.883
R1441 dvdd.t20 dvdd.t14 121.245
R1442 dvdd.t22 dvdd.t20 121.245
R1443 dvdd.t16 dvdd.t22 121.245
R1444 dvdd.t18 dvdd.t16 121.245
R1445 dvdd.t8 dvdd.t26 121.245
R1446 dvdd.t10 dvdd.t8 121.245
R1447 dvdd.t24 dvdd.t10 121.245
R1448 dvdd.t28 dvdd.t24 121.245
R1449 dvdd.n71 dvdd.t150 119.608
R1450 dvdd.n72 dvdd.t137 119.608
R1451 dvdd.n92 dvdd.t55 119.608
R1452 dvdd.n93 dvdd.t109 119.608
R1453 dvdd.n113 dvdd.t160 119.608
R1454 dvdd.n114 dvdd.t166 119.608
R1455 dvdd.t104 dvdd 109.1
R1456 dvdd.t125 dvdd 109.1
R1457 dvdd.t88 dvdd 109.1
R1458 dvdd.n75 dvdd.t151 108.413
R1459 dvdd.n76 dvdd.t135 108.413
R1460 dvdd.n96 dvdd.t57 108.413
R1461 dvdd.n97 dvdd.t108 108.413
R1462 dvdd.n117 dvdd.t158 108.413
R1463 dvdd.n118 dvdd.t168 108.413
R1464 dvdd.n271 dvdd.n55 106.559
R1465 dvdd.n272 dvdd.n54 106.559
R1466 dvdd.n273 dvdd.n53 106.559
R1467 dvdd.n47 dvdd.n2 105.412
R1468 dvdd.n40 dvdd.n2 105.412
R1469 dvdd.n37 dvdd.n36 105.412
R1470 dvdd.n36 dvdd.n35 105.412
R1471 dvdd dvdd.t117 100.624
R1472 dvdd.n67 dvdd.t144 93.81
R1473 dvdd.n68 dvdd.t51 93.81
R1474 dvdd.n88 dvdd.t67 93.81
R1475 dvdd.n89 dvdd.t121 93.81
R1476 dvdd.n109 dvdd.t82 93.81
R1477 dvdd.n110 dvdd.t170 93.81
R1478 dvdd dvdd.t115 91.745
R1479 dvdd dvdd.t140 91.745
R1480 dvdd dvdd.t30 88.7855
R1481 dvdd.n259 dvdd.t118 86.7743
R1482 dvdd.n47 dvdd.n46 79.8123
R1483 dvdd.n41 dvdd.n40 79.8123
R1484 dvdd.n35 dvdd.n34 79.8123
R1485 dvdd.n37 dvdd.n26 79.8123
R1486 dvdd.n59 dvdd.t78 74.7554
R1487 dvdd.n238 dvdd.t97 74.7554
R1488 dvdd.n67 dvdd.t43 63.3219
R1489 dvdd.n68 dvdd.t131 63.3219
R1490 dvdd.n71 dvdd.t45 63.3219
R1491 dvdd.n72 dvdd.t130 63.3219
R1492 dvdd.n88 dvdd.t39 63.3219
R1493 dvdd.n89 dvdd.t147 63.3219
R1494 dvdd.n92 dvdd.t41 63.3219
R1495 dvdd.n93 dvdd.t72 63.3219
R1496 dvdd.n109 dvdd.t47 63.3219
R1497 dvdd.n110 dvdd.t103 63.3219
R1498 dvdd.n113 dvdd.t37 63.3219
R1499 dvdd.n114 dvdd.t102 63.3219
R1500 dvdd.n79 dvdd.t152 61.9829
R1501 dvdd.n100 dvdd.t59 61.9829
R1502 dvdd.n122 dvdd.t162 61.9829
R1503 dvdd.n80 dvdd.t133 61.9826
R1504 dvdd.n101 dvdd.t110 61.9826
R1505 dvdd.n123 dvdd.t167 61.9826
R1506 dvdd.n259 dvdd.t120 61.05
R1507 dvdd.n294 dvdd.t18 60.6225
R1508 dvdd.t26 dvdd.n294 60.6225
R1509 dvdd.n292 dvdd.t15 60.3236
R1510 dvdd.n296 dvdd.t29 60.3236
R1511 dvdd.n297 dvdd.n283 54.7085
R1512 dvdd.n298 dvdd.n282 54.7085
R1513 dvdd.n290 dvdd.n289 54.7085
R1514 dvdd.n291 dvdd.n288 54.7085
R1515 dvdd.n61 dvdd.t79 41.5552
R1516 dvdd.n61 dvdd.t174 41.5552
R1517 dvdd.n62 dvdd.t71 41.5552
R1518 dvdd.n62 dvdd.t89 41.5552
R1519 dvdd.n82 dvdd.t171 41.5552
R1520 dvdd.n82 dvdd.t126 41.5552
R1521 dvdd.n83 dvdd.t114 41.5552
R1522 dvdd.n83 dvdd.t127 41.5552
R1523 dvdd.n103 dvdd.t99 41.5552
R1524 dvdd.n103 dvdd.t165 41.5552
R1525 dvdd.n104 dvdd.t63 41.5552
R1526 dvdd.n104 dvdd.t105 41.5552
R1527 dvdd.n46 dvdd.n45 37.0005
R1528 dvdd.n42 dvdd.n41 37.0005
R1529 dvdd.n34 dvdd.n33 37.0005
R1530 dvdd.n30 dvdd.n26 37.0005
R1531 dvdd.n17 dvdd.t116 36.1587
R1532 dvdd.n17 dvdd.t155 36.1587
R1533 dvdd.n8 dvdd.t141 36.1587
R1534 dvdd.n8 dvdd.t173 36.1587
R1535 dvdd.n256 dvdd.t96 35.4605
R1536 dvdd.n250 dvdd.n249 34.6358
R1537 dvdd.n254 dvdd.n245 34.6358
R1538 dvdd.n265 dvdd.n257 34.6358
R1539 dvdd.n231 dvdd.n63 34.6358
R1540 dvdd.n221 dvdd.n65 34.6358
R1541 dvdd.n225 dvdd.n65 34.6358
R1542 dvdd.n226 dvdd.n225 34.6358
R1543 dvdd.n219 dvdd.n218 34.6358
R1544 dvdd.n213 dvdd.n212 34.6358
R1545 dvdd.n214 dvdd.n213 34.6358
R1546 dvdd.n200 dvdd.n199 34.6358
R1547 dvdd.n202 dvdd.n77 34.6358
R1548 dvdd.n206 dvdd.n77 34.6358
R1549 dvdd.n193 dvdd.n84 34.6358
R1550 dvdd.n183 dvdd.n86 34.6358
R1551 dvdd.n187 dvdd.n86 34.6358
R1552 dvdd.n188 dvdd.n187 34.6358
R1553 dvdd.n181 dvdd.n180 34.6358
R1554 dvdd.n175 dvdd.n174 34.6358
R1555 dvdd.n176 dvdd.n175 34.6358
R1556 dvdd.n162 dvdd.n161 34.6358
R1557 dvdd.n164 dvdd.n98 34.6358
R1558 dvdd.n168 dvdd.n98 34.6358
R1559 dvdd.n155 dvdd.n105 34.6358
R1560 dvdd.n145 dvdd.n107 34.6358
R1561 dvdd.n149 dvdd.n107 34.6358
R1562 dvdd.n150 dvdd.n149 34.6358
R1563 dvdd.n143 dvdd.n142 34.6358
R1564 dvdd.n137 dvdd.n136 34.6358
R1565 dvdd.n138 dvdd.n137 34.6358
R1566 dvdd.n124 dvdd.n52 34.6358
R1567 dvdd.n126 dvdd.n119 34.6358
R1568 dvdd.n130 dvdd.n119 34.6358
R1569 dvdd.n239 dvdd.n58 33.8829
R1570 dvdd.n227 dvdd.n226 32.377
R1571 dvdd.n189 dvdd.n188 32.377
R1572 dvdd.n151 dvdd.n150 32.377
R1573 dvdd.n214 dvdd.n69 32.0005
R1574 dvdd.n176 dvdd.n90 32.0005
R1575 dvdd.n138 dvdd.n111 32.0005
R1576 dvdd.n240 dvdd.n239 31.624
R1577 dvdd.n202 dvdd.n201 31.2476
R1578 dvdd.n164 dvdd.n163 31.2476
R1579 dvdd.n126 dvdd.n125 31.2476
R1580 dvdd.n5 dvdd.n3 30.8338
R1581 dvdd.n4 dvdd.n2 30.8338
R1582 dvdd.n36 dvdd.n27 30.8338
R1583 dvdd.n29 dvdd.n28 30.8338
R1584 dvdd.n79 dvdd.t129 30.1745
R1585 dvdd.n100 dvdd.t84 30.1745
R1586 dvdd.n122 dvdd.t156 30.1745
R1587 dvdd.n80 dvdd.t5 30.1738
R1588 dvdd.n101 dvdd.t86 30.1738
R1589 dvdd.n123 dvdd.t34 30.1738
R1590 dvdd.n208 dvdd.n73 30.1181
R1591 dvdd.n170 dvdd.n94 30.1181
R1592 dvdd.n132 dvdd.n115 30.1181
R1593 dvdd.n43 dvdd.n42 29.6618
R1594 dvdd.n45 dvdd.n44 29.6618
R1595 dvdd.n31 dvdd.n30 29.6618
R1596 dvdd.n33 dvdd.n32 29.6618
R1597 dvdd.n59 dvdd.t143 28.5349
R1598 dvdd.n238 dvdd.t139 28.5349
R1599 dvdd.n261 dvdd.n257 28.2952
R1600 dvdd dvdd.n245 27.8593
R1601 dvdd.n256 dvdd.t94 26.5955
R1602 dvdd.n260 dvdd.n258 25.2079
R1603 dvdd.n22 dvdd.n18 23.7181
R1604 dvdd.n11 dvdd.n10 23.7181
R1605 dvdd.n249 dvdd.n246 23.7181
R1606 dvdd.n233 dvdd.n55 23.7181
R1607 dvdd.n199 dvdd.n54 23.7181
R1608 dvdd.n195 dvdd.n54 23.7181
R1609 dvdd.n161 dvdd.n53 23.7181
R1610 dvdd.n157 dvdd.n53 23.7181
R1611 dvdd.n274 dvdd.n52 23.7181
R1612 dvdd.n58 dvdd.n55 23.7181
R1613 dvdd.n232 dvdd.n231 22.9652
R1614 dvdd.n194 dvdd.n193 22.9652
R1615 dvdd.n156 dvdd.n155 22.9652
R1616 dvdd.n267 dvdd.n255 22.5887
R1617 dvdd.n266 dvdd.n265 22.5887
R1618 dvdd.n267 dvdd.n266 21.8358
R1619 dvdd.n233 dvdd.n232 21.4593
R1620 dvdd.n195 dvdd.n194 21.4593
R1621 dvdd.n157 dvdd.n156 21.4593
R1622 dvdd.n212 dvdd.n73 20.3299
R1623 dvdd.n174 dvdd.n94 20.3299
R1624 dvdd.n136 dvdd.n115 20.3299
R1625 dvdd.n255 dvdd.n254 19.9534
R1626 dvdd.n240 dvdd.n56 19.577
R1627 dvdd.n270 dvdd.n56 18.4476
R1628 dvdd.n227 dvdd.n63 18.0711
R1629 dvdd.n189 dvdd.n84 18.0711
R1630 dvdd.n151 dvdd.n105 18.0711
R1631 dvdd.n23 dvdd 15.8123
R1632 dvdd dvdd.n9 15.8123
R1633 dvdd.n296 dvdd.n295 13.2148
R1634 dvdd.n293 dvdd.n292 13.2148
R1635 dvdd.n38 dvdd.n37 10.0436
R1636 dvdd.n35 dvdd.n1 9.59217
R1637 dvdd.n218 dvdd.n69 9.41227
R1638 dvdd.n180 dvdd.n90 9.41227
R1639 dvdd.n142 dvdd.n111 9.41227
R1640 dvdd.n19 dvdd.n18 9.3005
R1641 dvdd.n22 dvdd.n21 9.3005
R1642 dvdd.n10 dvdd.n6 9.3005
R1643 dvdd.n12 dvdd.n11 9.3005
R1644 dvdd.n40 dvdd.n39 9.3005
R1645 dvdd.n48 dvdd.n47 9.3005
R1646 dvdd.n262 dvdd.n261 9.3005
R1647 dvdd.n263 dvdd.n257 9.3005
R1648 dvdd.n265 dvdd.n264 9.3005
R1649 dvdd.n266 dvdd.n243 9.3005
R1650 dvdd.n255 dvdd.n244 9.3005
R1651 dvdd.n254 dvdd.n253 9.3005
R1652 dvdd.n252 dvdd.n245 9.3005
R1653 dvdd.n251 dvdd.n250 9.3005
R1654 dvdd.n249 dvdd.n248 9.3005
R1655 dvdd.n247 dvdd.n246 9.3005
R1656 dvdd.n270 dvdd.n269 9.3005
R1657 dvdd.n275 dvdd.n274 9.3005
R1658 dvdd.n120 dvdd.n52 9.3005
R1659 dvdd.n124 dvdd.n121 9.3005
R1660 dvdd.n127 dvdd.n126 9.3005
R1661 dvdd.n128 dvdd.n119 9.3005
R1662 dvdd.n130 dvdd.n129 9.3005
R1663 dvdd.n131 dvdd.n116 9.3005
R1664 dvdd.n133 dvdd.n132 9.3005
R1665 dvdd.n134 dvdd.n115 9.3005
R1666 dvdd.n136 dvdd.n135 9.3005
R1667 dvdd.n137 dvdd.n112 9.3005
R1668 dvdd.n139 dvdd.n138 9.3005
R1669 dvdd.n140 dvdd.n111 9.3005
R1670 dvdd.n142 dvdd.n141 9.3005
R1671 dvdd.n143 dvdd.n108 9.3005
R1672 dvdd.n146 dvdd.n145 9.3005
R1673 dvdd.n147 dvdd.n107 9.3005
R1674 dvdd.n149 dvdd.n148 9.3005
R1675 dvdd.n150 dvdd.n106 9.3005
R1676 dvdd.n152 dvdd.n151 9.3005
R1677 dvdd.n153 dvdd.n105 9.3005
R1678 dvdd.n155 dvdd.n154 9.3005
R1679 dvdd.n156 dvdd.n102 9.3005
R1680 dvdd.n158 dvdd.n157 9.3005
R1681 dvdd.n159 dvdd.n53 9.3005
R1682 dvdd.n161 dvdd.n160 9.3005
R1683 dvdd.n162 dvdd.n99 9.3005
R1684 dvdd.n165 dvdd.n164 9.3005
R1685 dvdd.n166 dvdd.n98 9.3005
R1686 dvdd.n168 dvdd.n167 9.3005
R1687 dvdd.n169 dvdd.n95 9.3005
R1688 dvdd.n171 dvdd.n170 9.3005
R1689 dvdd.n172 dvdd.n94 9.3005
R1690 dvdd.n174 dvdd.n173 9.3005
R1691 dvdd.n175 dvdd.n91 9.3005
R1692 dvdd.n177 dvdd.n176 9.3005
R1693 dvdd.n178 dvdd.n90 9.3005
R1694 dvdd.n180 dvdd.n179 9.3005
R1695 dvdd.n181 dvdd.n87 9.3005
R1696 dvdd.n184 dvdd.n183 9.3005
R1697 dvdd.n185 dvdd.n86 9.3005
R1698 dvdd.n187 dvdd.n186 9.3005
R1699 dvdd.n188 dvdd.n85 9.3005
R1700 dvdd.n190 dvdd.n189 9.3005
R1701 dvdd.n191 dvdd.n84 9.3005
R1702 dvdd.n193 dvdd.n192 9.3005
R1703 dvdd.n194 dvdd.n81 9.3005
R1704 dvdd.n196 dvdd.n195 9.3005
R1705 dvdd.n197 dvdd.n54 9.3005
R1706 dvdd.n199 dvdd.n198 9.3005
R1707 dvdd.n200 dvdd.n78 9.3005
R1708 dvdd.n203 dvdd.n202 9.3005
R1709 dvdd.n204 dvdd.n77 9.3005
R1710 dvdd.n206 dvdd.n205 9.3005
R1711 dvdd.n207 dvdd.n74 9.3005
R1712 dvdd.n209 dvdd.n208 9.3005
R1713 dvdd.n210 dvdd.n73 9.3005
R1714 dvdd.n212 dvdd.n211 9.3005
R1715 dvdd.n213 dvdd.n70 9.3005
R1716 dvdd.n215 dvdd.n214 9.3005
R1717 dvdd.n216 dvdd.n69 9.3005
R1718 dvdd.n218 dvdd.n217 9.3005
R1719 dvdd.n219 dvdd.n66 9.3005
R1720 dvdd.n222 dvdd.n221 9.3005
R1721 dvdd.n223 dvdd.n65 9.3005
R1722 dvdd.n225 dvdd.n224 9.3005
R1723 dvdd.n226 dvdd.n64 9.3005
R1724 dvdd.n228 dvdd.n227 9.3005
R1725 dvdd.n229 dvdd.n63 9.3005
R1726 dvdd.n231 dvdd.n230 9.3005
R1727 dvdd.n232 dvdd.n60 9.3005
R1728 dvdd.n234 dvdd.n233 9.3005
R1729 dvdd.n235 dvdd.n55 9.3005
R1730 dvdd.n236 dvdd.n58 9.3005
R1731 dvdd.n239 dvdd.n237 9.3005
R1732 dvdd.n239 dvdd.n57 9.3005
R1733 dvdd.n241 dvdd.n240 9.3005
R1734 dvdd.n242 dvdd.n56 9.3005
R1735 dvdd.n268 dvdd.n267 9.3005
R1736 dvdd.n208 dvdd.n207 9.03579
R1737 dvdd.n170 dvdd.n169 9.03579
R1738 dvdd.n132 dvdd.n131 9.03579
R1739 dvdd.n286 dvdd.n284 7.70883
R1740 dvdd.n294 dvdd.n286 7.70883
R1741 dvdd.n287 dvdd.n285 7.70883
R1742 dvdd.n294 dvdd.n287 7.70883
R1743 dvdd.n24 dvdd.n23 7.17001
R1744 dvdd.n9 dvdd.n7 7.15376
R1745 dvdd.n283 dvdd.t11 7.14175
R1746 dvdd.n283 dvdd.t25 7.14175
R1747 dvdd.n282 dvdd.t27 7.14175
R1748 dvdd.n282 dvdd.t9 7.14175
R1749 dvdd.n289 dvdd.t17 7.14175
R1750 dvdd.n289 dvdd.t19 7.14175
R1751 dvdd.n288 dvdd.t21 7.14175
R1752 dvdd.n288 dvdd.t23 7.14175
R1753 dvdd.n250 dvdd 6.77697
R1754 dvdd.n44 dvdd.t48 6.70818
R1755 dvdd.t48 dvdd.n43 6.70818
R1756 dvdd.n32 dvdd.t12 6.70818
R1757 dvdd.t12 dvdd.n31 6.70818
R1758 dvdd dvdd.n22 6.4005
R1759 dvdd.n10 dvdd 6.4005
R1760 dvdd.n221 dvdd.n220 6.02403
R1761 dvdd.n207 dvdd.n206 6.02403
R1762 dvdd.n183 dvdd.n182 6.02403
R1763 dvdd.n169 dvdd.n168 6.02403
R1764 dvdd.n145 dvdd.n144 6.02403
R1765 dvdd.n131 dvdd.n130 6.02403
R1766 dvdd.n220 dvdd.n219 3.76521
R1767 dvdd.n182 dvdd.n181 3.76521
R1768 dvdd.n144 dvdd.n143 3.76521
R1769 dvdd.n201 dvdd.n200 3.38874
R1770 dvdd.n163 dvdd.n162 3.38874
R1771 dvdd.n125 dvdd.n124 3.38874
R1772 dvdd.n297 dvdd.n296 1.66909
R1773 dvdd.n292 dvdd.n291 1.57188
R1774 dvdd.n36 dvdd.n0 1.32907
R1775 dvdd.n2 dvdd.n0 1.32907
R1776 dvdd.n261 dvdd.n260 1.23559
R1777 dvdd.n276 dvdd.n275 0.637387
R1778 dvdd.n276 dvdd.n51 0.496845
R1779 dvdd dvdd.n268 0.438
R1780 dvdd.n50 dvdd.n49 0.432317
R1781 dvdd.n16 dvdd 0.42713
R1782 dvdd dvdd.n16 0.32387
R1783 dvdd.n268 dvdd 0.313
R1784 dvdd.n247 dvdd.n51 0.280448
R1785 dvdd.n51 dvdd 0.232271
R1786 dvdd.n7 dvdd 0.203706
R1787 dvdd.n13 dvdd 0.167167
R1788 dvdd.n19 dvdd 0.164848
R1789 dvdd.n258 dvdd 0.159538
R1790 dvdd.n38 dvdd.n15 0.141704
R1791 dvdd.n262 dvdd.n258 0.141672
R1792 dvdd.n38 dvdd.n25 0.139389
R1793 dvdd.n14 dvdd.n6 0.127236
R1794 dvdd.n264 dvdd.n243 0.120292
R1795 dvdd.n252 dvdd.n251 0.120292
R1796 dvdd.n253 dvdd.n252 0.120292
R1797 dvdd.n253 dvdd.n244 0.120292
R1798 dvdd.n121 dvdd.n120 0.120292
R1799 dvdd.n127 dvdd.n121 0.120292
R1800 dvdd.n128 dvdd.n127 0.120292
R1801 dvdd.n129 dvdd.n128 0.120292
R1802 dvdd.n129 dvdd.n116 0.120292
R1803 dvdd.n133 dvdd.n116 0.120292
R1804 dvdd.n134 dvdd.n133 0.120292
R1805 dvdd.n135 dvdd.n134 0.120292
R1806 dvdd.n135 dvdd.n112 0.120292
R1807 dvdd.n139 dvdd.n112 0.120292
R1808 dvdd.n140 dvdd.n139 0.120292
R1809 dvdd.n141 dvdd.n140 0.120292
R1810 dvdd.n141 dvdd.n108 0.120292
R1811 dvdd.n146 dvdd.n108 0.120292
R1812 dvdd.n147 dvdd.n146 0.120292
R1813 dvdd.n148 dvdd.n147 0.120292
R1814 dvdd.n148 dvdd.n106 0.120292
R1815 dvdd.n152 dvdd.n106 0.120292
R1816 dvdd.n153 dvdd.n152 0.120292
R1817 dvdd.n154 dvdd.n153 0.120292
R1818 dvdd.n154 dvdd.n102 0.120292
R1819 dvdd.n158 dvdd.n102 0.120292
R1820 dvdd.n160 dvdd.n99 0.120292
R1821 dvdd.n165 dvdd.n99 0.120292
R1822 dvdd.n166 dvdd.n165 0.120292
R1823 dvdd.n167 dvdd.n166 0.120292
R1824 dvdd.n167 dvdd.n95 0.120292
R1825 dvdd.n171 dvdd.n95 0.120292
R1826 dvdd.n172 dvdd.n171 0.120292
R1827 dvdd.n173 dvdd.n172 0.120292
R1828 dvdd.n173 dvdd.n91 0.120292
R1829 dvdd.n177 dvdd.n91 0.120292
R1830 dvdd.n178 dvdd.n177 0.120292
R1831 dvdd.n179 dvdd.n178 0.120292
R1832 dvdd.n179 dvdd.n87 0.120292
R1833 dvdd.n184 dvdd.n87 0.120292
R1834 dvdd.n185 dvdd.n184 0.120292
R1835 dvdd.n186 dvdd.n185 0.120292
R1836 dvdd.n186 dvdd.n85 0.120292
R1837 dvdd.n190 dvdd.n85 0.120292
R1838 dvdd.n191 dvdd.n190 0.120292
R1839 dvdd.n192 dvdd.n191 0.120292
R1840 dvdd.n192 dvdd.n81 0.120292
R1841 dvdd.n196 dvdd.n81 0.120292
R1842 dvdd.n198 dvdd.n78 0.120292
R1843 dvdd.n203 dvdd.n78 0.120292
R1844 dvdd.n204 dvdd.n203 0.120292
R1845 dvdd.n205 dvdd.n204 0.120292
R1846 dvdd.n205 dvdd.n74 0.120292
R1847 dvdd.n209 dvdd.n74 0.120292
R1848 dvdd.n210 dvdd.n209 0.120292
R1849 dvdd.n211 dvdd.n210 0.120292
R1850 dvdd.n211 dvdd.n70 0.120292
R1851 dvdd.n215 dvdd.n70 0.120292
R1852 dvdd.n216 dvdd.n215 0.120292
R1853 dvdd.n217 dvdd.n216 0.120292
R1854 dvdd.n217 dvdd.n66 0.120292
R1855 dvdd.n222 dvdd.n66 0.120292
R1856 dvdd.n223 dvdd.n222 0.120292
R1857 dvdd.n224 dvdd.n223 0.120292
R1858 dvdd.n224 dvdd.n64 0.120292
R1859 dvdd.n228 dvdd.n64 0.120292
R1860 dvdd.n229 dvdd.n228 0.120292
R1861 dvdd.n230 dvdd.n229 0.120292
R1862 dvdd.n230 dvdd.n60 0.120292
R1863 dvdd.n234 dvdd.n60 0.120292
R1864 dvdd.n237 dvdd.n236 0.120292
R1865 dvdd.n241 dvdd.n57 0.120292
R1866 dvdd.n242 dvdd.n241 0.120292
R1867 dvdd.n277 dvdd.n276 0.109494
R1868 dvdd.n15 dvdd.n14 0.109053
R1869 dvdd.n268 dvdd.n244 0.107271
R1870 dvdd.n14 dvdd 0.0983618
R1871 dvdd dvdd.n262 0.0981562
R1872 dvdd.n251 dvdd 0.0968542
R1873 dvdd.n281 dvdd.n280 0.0944312
R1874 dvdd.n278 dvdd.n277 0.0856755
R1875 dvdd.n279 dvdd.n278 0.0856755
R1876 dvdd.n237 dvdd 0.0812292
R1877 dvdd dvdd.n6 0.0803611
R1878 dvdd.n280 dvdd.n279 0.0777774
R1879 dvdd.n14 dvdd.n7 0.070241
R1880 dvdd.n25 dvdd.n24 0.0685285
R1881 dvdd.n268 dvdd 0.063
R1882 dvdd.n264 dvdd 0.0603958
R1883 dvdd dvdd.n263 0.0603958
R1884 dvdd.n248 dvdd 0.0603958
R1885 dvdd.n120 dvdd 0.0603958
R1886 dvdd.n159 dvdd 0.0603958
R1887 dvdd.n160 dvdd 0.0603958
R1888 dvdd.n197 dvdd 0.0603958
R1889 dvdd.n198 dvdd 0.0603958
R1890 dvdd.n235 dvdd 0.0603958
R1891 dvdd.n236 dvdd 0.0603958
R1892 dvdd.n269 dvdd 0.0603958
R1893 dvdd dvdd.n13 0.0595278
R1894 dvdd.n21 dvdd.n16 0.0535523
R1895 dvdd.n12 dvdd 0.0508472
R1896 dvdd.n291 dvdd.n290 0.0456945
R1897 dvdd.n39 dvdd.n38 0.0456858
R1898 dvdd.n20 dvdd 0.0405
R1899 dvdd dvdd.n57 0.0395625
R1900 dvdd dvdd.n297 0.0385435
R1901 dvdd dvdd.n247 0.0382604
R1902 dvdd.n39 dvdd.n0 0.0379437
R1903 dvdd.n21 dvdd 0.0339302
R1904 dvdd.n13 dvdd.n12 0.0334861
R1905 dvdd.n275 dvdd 0.03175
R1906 dvdd dvdd.n159 0.03175
R1907 dvdd dvdd.n197 0.03175
R1908 dvdd dvdd.n235 0.03175
R1909 dvdd.n269 dvdd 0.03175
R1910 dvdd.n24 dvdd.n16 0.0300191
R1911 dvdd.n248 dvdd 0.0239375
R1912 dvdd.n49 dvdd.n0 0.0233041
R1913 dvdd.n263 dvdd 0.0226354
R1914 dvdd dvdd.n158 0.0226354
R1915 dvdd dvdd.n196 0.0226354
R1916 dvdd dvdd.n234 0.0226354
R1917 dvdd dvdd.n242 0.0226354
R1918 dvdd.n299 dvdd.n298 0.0219531
R1919 dvdd.n15 dvdd 0.0210592
R1920 dvdd.n20 dvdd.n19 0.0205
R1921 dvdd.n48 dvdd.n1 0.0182365
R1922 dvdd.n25 dvdd 0.0179419
R1923 dvdd.n49 dvdd.n48 0.0151396
R1924 dvdd.n290 dvdd.n281 0.0150881
R1925 dvdd dvdd.n20 0.0121279
R1926 dvdd.n299 dvdd.n281 0.00936728
R1927 dvdd.n268 dvdd.n243 0.0083125
R1928 dvdd.n277 dvdd.t178 0.0083125
R1929 dvdd.n278 dvdd.t177 0.0083125
R1930 dvdd.n279 dvdd.t176 0.0083125
R1931 dvdd.n50 dvdd.t175 0.0083125
R1932 dvdd.n298 dvdd 0.00765103
R1933 dvdd.n280 dvdd.n50 0.00754239
R1934 dvdd.n1 dvdd 0.00176689
R1935 dvdd.n299 dvdd 0.001125
R1936 icnode.t1 icnode.t0 84.1171
R1937 vbreg.n21 vbreg.t0 244.944
R1938 vbreg.n49 vbreg.n2 202.542
R1939 vbreg.n40 vbreg.n10 201.036
R1940 vbreg.n33 vbreg.n7 200.282
R1941 vbreg.n20 vbreg.n21 0.962138
R1942 vbreg.n35 vbreg.n10 179.201
R1943 vbreg.n2 vbreg.n24 178.447
R1944 vbreg.n35 vbreg.n7 176.941
R1945 vbreg.n42 vbreg.n24 160.376
R1946 vbreg.n35 vbreg.n19 116.609
R1947 vbreg.n35 vbreg.n15 116.609
R1948 vbreg.n30 vbreg.n10 116.609
R1949 vbreg.n17 vbreg.n10 116.609
R1950 vbreg.n44 vbreg.n24 116.609
R1951 vbreg.n56 vbreg.n24 116.609
R1952 vbreg.n53 vbreg.n2 116.609
R1953 vbreg.n2 vbreg.n25 116.609
R1954 vbreg.n18 vbreg.n7 116.609
R1955 vbreg.n16 vbreg.n7 116.609
R1956 vbreg.n42 vbreg.n26 115.005
R1957 vbreg.n42 vbreg.n40 110.683
R1958 vbreg.t13 vbreg.n31 86.3125
R1959 vbreg.n14 vbreg.t10 88.4838
R1960 vbreg.n18 vbreg.t14 86.3125
R1961 vbreg.t12 vbreg.n16 86.3125
R1962 vbreg.t23 vbreg.n12 88.4979
R1963 vbreg.n51 vbreg.t25 86.3125
R1964 vbreg.t17 vbreg.n38 86.3125
R1965 vbreg.n28 vbreg.t18 86.3125
R1966 vbreg.n15 vbreg.t9 86.3125
R1967 vbreg.n19 vbreg.t11 86.3125
R1968 vbreg.n37 vbreg.t15 86.3125
R1969 vbreg.n29 vbreg.t16 86.3125
R1970 vbreg.n57 vbreg.t7 86.3125
R1971 vbreg.n43 vbreg.t20 86.3125
R1972 vbreg.n55 vbreg.t19 86.3125
R1973 vbreg.n54 vbreg.t22 86.3125
R1974 vbreg.n47 vbreg.t21 86.3125
R1975 vbreg.n52 vbreg.t24 86.3125
R1976 vbreg.n16 vbreg.n14 2.64048
R1977 vbreg.n38 vbreg.n37 72.5338
R1978 vbreg.n12 vbreg.n47 2.18593
R1979 vbreg.n18 vbreg.n31 72.5338
R1980 vbreg.n29 vbreg.n28 72.5338
R1981 vbreg.n52 vbreg.n51 72.5338
R1982 vbreg.n15 vbreg.n17 71.7809
R1983 vbreg.n57 vbreg.n56 71.7809
R1984 vbreg.n19 vbreg.n30 71.7809
R1985 vbreg.n28 vbreg.n26 71.7809
R1986 vbreg.n44 vbreg.n43 71.7809
R1987 vbreg.n16 vbreg.n15 71.5299
R1988 vbreg.n13 vbreg.n18 2.62088
R1989 vbreg.n55 vbreg.n25 71.2789
R1990 vbreg.n54 vbreg.n53 71.2789
R1991 vbreg.n38 vbreg.n23 60.7378
R1992 vbreg.n11 vbreg.t8 60.1061
R1993 vbreg.n32 vbreg.t13 55.9125
R1994 vbreg.n32 vbreg.t10 55.9125
R1995 vbreg.t14 vbreg.n34 55.9125
R1996 vbreg.n34 vbreg.t12 55.9125
R1997 vbreg.n48 vbreg.t23 55.9125
R1998 vbreg.n48 vbreg.t25 55.9125
R1999 vbreg.n39 vbreg.t17 55.9125
R2000 vbreg.n39 vbreg.t18 55.9125
R2001 vbreg.t9 vbreg.n36 55.9125
R2002 vbreg.n36 vbreg.t11 55.9125
R2003 vbreg.n27 vbreg.t15 55.9125
R2004 vbreg.t16 vbreg.n27 55.9125
R2005 vbreg.n41 vbreg.t7 55.9125
R2006 vbreg.n41 vbreg.t20 55.9125
R2007 vbreg.n45 vbreg.t19 55.9125
R2008 vbreg.t22 vbreg.n45 55.9125
R2009 vbreg.t21 vbreg.n46 55.9125
R2010 vbreg.n46 vbreg.t24 55.9125
R2011 vbreg.n33 vbreg.n32 30.4005
R2012 vbreg.n49 vbreg.n48 30.4005
R2013 vbreg.n36 vbreg.n35 30.4005
R2014 vbreg.n27 vbreg.n10 30.4005
R2015 vbreg.n40 vbreg.n39 30.4005
R2016 vbreg.n42 vbreg.n41 30.4005
R2017 vbreg.n45 vbreg.n24 30.4005
R2018 vbreg.n46 vbreg.n2 30.4005
R2019 vbreg.n34 vbreg.n7 30.4005
R2020 vbreg.n21 vbreg.t1 22.4019
R2021 vbreg.n22 vbreg.t5 21.1527
R2022 vbreg.n21 vbreg.t6 21.0621
R2023 vbreg.n42 vbreg.n11 2.00645
R2024 vbreg.n11 vbreg.n23 15.0573
R2025 vbreg.n57 vbreg.n23 11.7966
R2026 vbreg.n21 vbreg.n22 0.632464
R2027 vbreg.n40 vbreg.n3 3.01598
R2028 vbreg.n51 vbreg.n50 2.92951
R2029 vbreg.n4 vbreg.n31 2.92951
R2030 vbreg.n50 vbreg.n49 2.3255
R2031 vbreg.n0 vbreg.n2 2.3255
R2032 vbreg.n38 vbreg.n3 2.3255
R2033 vbreg.n55 vbreg.n3 2.3255
R2034 vbreg.n0 vbreg.n54 2.3255
R2035 vbreg.n52 vbreg.n0 2.3255
R2036 vbreg.n4 vbreg.n33 2.3255
R2037 vbreg.n5 vbreg.n7 2.3255
R2038 vbreg.n37 vbreg.n9 2.3255
R2039 vbreg.n9 vbreg.n10 2.3255
R2040 vbreg.n29 vbreg.n9 2.3255
R2041 vbreg.n28 vbreg.n8 2.3255
R2042 vbreg.n43 vbreg.n8 2.3255
R2043 vbreg.n3 vbreg.n57 2.3255
R2044 vbreg.n8 vbreg.n11 1.77359
R2045 vbreg.n3 vbreg.n20 1.69825
R2046 vbreg.n47 vbreg.n25 1.2554
R2047 vbreg.n53 vbreg.n52 1.2554
R2048 vbreg.n20 vbreg.t2 21.8362
R2049 vbreg.n21 vbreg.t4 21.6418
R2050 vbreg.n22 vbreg.t3 21.6076
R2051 vbreg.n19 vbreg.n13 2.62088
R2052 vbreg.n9 vbreg.n15 2.82746
R2053 vbreg.n6 vbreg.n5 0.489702
R2054 vbreg.n9 vbreg.n6 0.553315
R2055 vbreg.n1 vbreg.n0 0.420519
R2056 vbreg.n9 vbreg.n8 1.22324
R2057 vbreg.n6 vbreg.n35 2.715
R2058 vbreg.n12 vbreg.n0 1.45199
R2059 vbreg.n50 vbreg.n0 1.13148
R2060 vbreg.n5 vbreg.n4 1.12454
R2061 vbreg.n1 vbreg.n3 0.237615
R2062 vbreg.n5 vbreg.n13 0.795018
R2063 vbreg.n14 vbreg.n5 0.776083
R2064 vbreg.n3 vbreg.n11 0.753999
R2065 vbreg.n37 vbreg.n17 0.753441
R2066 vbreg.n56 vbreg.n55 0.753441
R2067 vbreg.n30 vbreg.n29 0.753441
R2068 vbreg.n43 vbreg.n26 0.753441
R2069 vbreg.n54 vbreg.n44 0.753441
R2070 vbreg.n1 vbreg.n24 2.61619
R2071 vbp.n3 vbp.n4 26.3414
R2072 vbp.n0 vbp 26.2397
R2073 vbp vbp.t1 112.21
R2074 vbp.n5 vbp.t12 21.3971
R2075 vbp.t10 vbp.n7 21.2714
R2076 vbp.n1 vbp.t13 21.3971
R2077 vbp.n3 vbp.n6 8.08368
R2078 vbp.n3 vbp.n5 8.21681
R2079 vbp.t17 vbp.n4 16.1817
R2080 vbp vbp.n2 8.77241
R2081 vbp vbp.t2 40.0025
R2082 vbp.t6 vbp 21.3013
R2083 vbp vbp.t16 21.3065
R2084 vbp.t3 vbp.n7 21.3313
R2085 vbp.n6 vbp.t14 21.0504
R2086 vbp.t4 vbp.n6 21.0498
R2087 vbp.n5 vbp.t7 20.9537
R2088 vbp.t11 vbp.n4 33.1891
R2089 vbp.t0 vbp.n2 21.7234
R2090 vbp.t9 vbp.n2 21.1857
R2091 vbp.t8 vbp.n1 20.9537
R2092 vbp.n0 vbp.t15 33.1158
R2093 vbp.n7 vbp 17.5035
R2094 vbp.n3 vbp 12.5283
R2095 vbp.n0 vbp.t5 16.2176
R2096 vbp vbp.n1 13.871
R2097 tail.n2 tail.t3 113.688
R2098 tail tail.t4 113.688
R2099 tail tail.t6 113.624
R2100 tail.n0 tail.t2 113.562
R2101 tail.n0 tail.t7 113.562
R2102 tail.n1 tail.t5 113.562
R2103 tail.n1 tail.t0 113.562
R2104 tail tail.t1 113.501
R2105 tail.n2 tail.t8 113.438
R2106 tail tail.t9 113.438
R2107 tail tail.n3 53.5531
R2108 tail.n3 tail.t10 6.92425
R2109 tail.n3 tail.t11 6.92425
R2110 tail tail.n1 1.9055
R2111 tail.n1 tail.n0 1.13844
R2112 tail tail.n2 1.13636
R2113 standby_b.n18 standby_b.t14 408.63
R2114 standby_b.n20 standby_b.t25 408.63
R2115 standby_b.n22 standby_b.t11 408.63
R2116 standby_b.n12 standby_b.t6 401.051
R2117 standby_b.t6 standby_b.n11 401.051
R2118 standby_b.t19 standby_b.n3 401.051
R2119 standby_b.n4 standby_b.t19 401.051
R2120 standby_b.n12 standby_b.t16 371.31
R2121 standby_b.t16 standby_b.n11 371.31
R2122 standby_b.t18 standby_b.n13 371.31
R2123 standby_b.n14 standby_b.t18 371.31
R2124 standby_b.t0 standby_b.n10 371.31
R2125 standby_b.n15 standby_b.t0 371.31
R2126 standby_b.n17 standby_b.t3 371.31
R2127 standby_b.t3 standby_b.n16 371.31
R2128 standby_b.n9 standby_b.t21 371.31
R2129 standby_b.t21 standby_b.n8 371.31
R2130 standby_b.t23 standby_b.n2 371.31
R2131 standby_b.n7 standby_b.t23 371.31
R2132 standby_b.t7 standby_b.n5 371.31
R2133 standby_b.n6 standby_b.t7 371.31
R2134 standby_b.n4 standby_b.t17 371.31
R2135 standby_b.t17 standby_b.n3 371.31
R2136 standby_b.n26 standby_b.t13 347.577
R2137 standby_b.n25 standby_b.t15 347.577
R2138 standby_b.n24 standby_b.t2 347.577
R2139 standby_b.n0 standby_b.t12 332.752
R2140 standby_b.t12 x4.in_b 332.752
R2141 standby_b.n0 standby_b.t4 332.411
R2142 standby_b.t4 x4.in_b 332.411
R2143 standby_b.n27 standby_b.t24 236.552
R2144 standby_b.n26 standby_b.t8 193.337
R2145 standby_b.n25 standby_b.t9 193.337
R2146 standby_b.n24 standby_b.t22 193.337
R2147 x7.x2.x4.RESET_B standby_b.n18 165.089
R2148 x7.x2.x4.RESET_B standby_b.n20 165.089
R2149 x7.x2.x4.RESET_B standby_b.n22 165.089
R2150 standby_b.n27 standby_b.t10 164.251
R2151 x7.x3.A1 standby_b.n27 154.47
R2152 x7.x2.x2.RESET_B standby_b.n26 152
R2153 x7.x2.x3.RESET_B standby_b.n25 152
R2154 x7.x2.x4.RESET_B standby_b.n24 152
R2155 standby_b.n18 standby_b.t1 132.282
R2156 standby_b.n20 standby_b.t5 132.282
R2157 standby_b.n22 standby_b.t20 132.282
R2158 standby_b.n6 standby_b.n3 29.7417
R2159 standby_b.n7 standby_b.n6 29.7417
R2160 standby_b.n8 standby_b.n7 29.7417
R2161 standby_b.n16 standby_b.n15 29.7417
R2162 standby_b.n15 standby_b.n14 29.7417
R2163 standby_b.n14 standby_b.n11 29.7417
R2164 standby_b.n5 standby_b.n4 29.7417
R2165 standby_b.n5 standby_b.n2 29.7417
R2166 standby_b.n9 standby_b.n2 29.7417
R2167 standby_b.n17 standby_b.n10 29.7417
R2168 standby_b.n13 standby_b.n10 29.7417
R2169 standby_b.n13 standby_b.n12 29.7417
R2170 standby_b.n8 standby_b.n1 17.6946
R2171 standby_b.n1 standby_b.n9 17.5064
R2172 standby_b.n19 x7.x2.x4.RESET_B 16.7098
R2173 standby_b.n1 x7.stby_b 15.0825
R2174 x7.x2.x2.RESET_B standby_b.n19 14.0185
R2175 x7.x2.x3.RESET_B standby_b.n21 14.0185
R2176 x7.x2.x4.RESET_B standby_b.n23 14.0185
R2177 x7.stby_b x7.x3.A1 13.8064
R2178 standby_b.n1 standby_b.n17 12.2358
R2179 standby_b.n16 standby_b.n1 12.0476
R2180 standby_b.n19 x7.x2.x2.RESET_B 11.4672
R2181 standby_b.n21 x7.x2.x3.RESET_B 11.4672
R2182 standby_b.n23 x7.x2.x4.RESET_B 11.4672
R2183 x4.in_b standby_b.n0 11.1417
R2184 x7.stby_b x7.x2.x4.RESET_B 10.5569
R2185 x4.in_b standby_b.n1 10.4718
R2186 standby_b.n23 x7.x2.x4.RESET_B 9.3005
R2187 x7.x2.x4.RESET_B x7.x2.x3.RESET_B 9.3005
R2188 standby_b.n21 x7.x2.x4.RESET_B 9.3005
R2189 x7.x2.x4.RESET_B x7.x2.x2.RESET_B 9.3005
R2190 a_9120_n9346.n1 a_9120_n9346.t3 649.659
R2191 a_9120_n9346.n0 a_9120_n9346.t1 227.685
R2192 a_9120_n9346.t4 a_9120_n9346.n2 44.6806
R2193 a_9120_n9346.n1 a_9120_n9346.t2 5.45407
R2194 a_9120_n9346.n0 a_9120_n9346.t0 5.07473
R2195 a_9120_n9346.n2 a_9120_n9346.n0 0.639781
R2196 a_9120_n9346.n2 a_9120_n9346.n1 0.0621233
R2197 x7.ena_done_b.n8 x7.ena_done_b.t1 373.866
R2198 x7.ena_done_b.n6 x7.ena_done_b.t5 333.651
R2199 x7.ena_done_b.n6 x7.ena_done_b.t6 297.233
R2200 x7.ena_done_b x7.ena_done_b.t0 247.159
R2201 x7.ena_done_b.n0 x7.ena_done_b.t3 241.536
R2202 x7.ena_done_b.n2 x7.ena_done_b.t4 207.423
R2203 x7.ena_done_b.n3 x7.ena_done_b.t7 202.133
R2204 x7.ena_done_b x7.ena_done_b.n6 195.701
R2205 x7.ena_done_b.n0 x7.ena_done_b.t2 169.237
R2206 x7.ena_done_b.n5 x7.ena_done_b.n2 159.758
R2207 x7.ena_done_b.n1 x7.ena_done_b.n0 155.84
R2208 x7.ena_done_b.n4 x7.ena_done_b.n3 152
R2209 x7.ena_done_b.n3 x7.ena_done_b.n2 36.8275
R2210 x7.ena_done_b x7.ena_done_b.n8 16.6907
R2211 x7.ena_done_b.n7 x7.ena_done_b 15.8995
R2212 x7.ena_done_b.n7 x7.ena_done_b 15.6656
R2213 x7.ena_done_b x7.ena_done_b.n5 13.8109
R2214 x7.ena_done_b x7.ena_done_b.n1 11.2245
R2215 x7.ena_done_b.n5 x7.ena_done_b.n4 5.4308
R2216 x7.ena_done_b.n4 x7.ena_done_b 3.68535
R2217 x7.ena_done_b.n1 x7.ena_done_b 3.2005
R2218 x7.ena_done_b.n8 x7.ena_done_b.n7 3.1005
R2219 standby_33.n0 standby_33.t0 227.886
R2220 standby_33 standby_33.t3 216.05
R2221 standby_33.n0 standby_33.n1 25.0903
R2222 standby_33.n0 standby_33.t4 12.7763
R2223 standby_33.n1 standby_33.t1 5.5105
R2224 standby_33.n1 standby_33.t2 5.5105
R2225 standby_33.n0 standby_33 1.67737
R2226 ibias.n7 ibias.n1 1544.9
R2227 ibias.n4 ibias.n3 1544.9
R2228 ibias.n2 ibias.n0 300.425
R2229 ibias.n8 ibias.n2 300.425
R2230 ibias.n9 ibias.n0 177.746
R2231 ibias.n9 ibias.n8 177.746
R2232 ibias.n5 ibias.n1 139.143
R2233 ibias.n6 ibias.n3 139.143
R2234 ibias.n9 ibias.t1 60.1061
R2235 ibias.n4 ibias.n0 46.2505
R2236 ibias.n8 ibias.n7 46.2505
R2237 ibias.n5 ibias.n4 40.8622
R2238 ibias.n7 ibias.n6 40.8622
R2239 ibias.n3 ibias.n2 12.3338
R2240 ibias.n9 ibias.n1 12.3338
R2241 ibias.n6 ibias.t0 4.16651
R2242 ibias.t0 ibias.n5 4.16651
R2243 ibias ibias.n9 1.58676
R2244 ibias_ip ibias_ip.t13 31.8332
R2245 ibias_ip.t12 ibias_ip 31.4808
R2246 ibias_ip ibias_ip.t10 61.7027
R2247 ibias_ip.t0 ibias_ip 31.3394
R2248 ibias_ip ibias_ip.t1 39.498
R2249 ibias_ip.n0 ibias_ip.t11 31.8633
R2250 ibias_ip ibias_ip.t6 31.1832
R2251 ibias_ip.n1 ibias_ip.t2 31.1727
R2252 ibias_ip.n0 ibias_ip.t8 31.193
R2253 ibias_ip.n0 ibias_ip.t4 31.1967
R2254 ibias_ip.t3 ibias_ip.n1 39.8957
R2255 ibias_ip ibias_ip.t7 39.8329
R2256 ibias_ip.t5 ibias_ip.n0 39.8506
R2257 ibias_ip.n0 ibias_ip.t9 39.8715
R2258 ibias_ip ibias_ip.n1 1.87886
R2259 ibias_ip ibias_ip.n0 1.34188
R2260 avdd_ip.n81 avdd_ip.n73 58547.9
R2261 avdd_ip.n81 avdd_ip.n80 58547.9
R2262 avdd_ip.n79 avdd_ip.n73 58547.9
R2263 avdd_ip.n80 avdd_ip.n79 58547.9
R2264 avdd_ip.n43 avdd_ip.n42 54381
R2265 avdd_ip.n82 avdd_ip.n71 28978.4
R2266 avdd_ip.n82 avdd_ip.n72 28978.4
R2267 avdd_ip.n78 avdd_ip.n71 28978.4
R2268 avdd_ip.n78 avdd_ip.n72 28978.4
R2269 avdd_ip.n93 avdd_ip.n26 7296
R2270 avdd_ip.n91 avdd_ip.n26 7296
R2271 avdd_ip.n93 avdd_ip.n27 7296
R2272 avdd_ip.n91 avdd_ip.n27 7296
R2273 avdd_ip.n77 avdd_ip.n75 5062.04
R2274 avdd_ip.n75 avdd_ip.n74 3209.98
R2275 avdd_ip.n76 avdd_ip.n62 1005.14
R2276 avdd_ip.n44 avdd_ip.n36 857.648
R2277 avdd_ip.n40 avdd_ip.n37 857.648
R2278 avdd_ip.n44 avdd_ip.n37 857.648
R2279 avdd_ip.n55 avdd_ip.n54 857.648
R2280 avdd_ip.n57 avdd_ip.n50 857.648
R2281 avdd_ip.n43 avdd_ip.t2 337.433
R2282 avdd_ip.n77 avdd_ip.n76 269.44
R2283 avdd_ip.n57 avdd_ip.n56 267.182
R2284 avdd_ip.n54 avdd_ip.n51 267.182
R2285 avdd_ip.n41 avdd_ip.n40 267.182
R2286 avdd_ip.n84 avdd_ip.n63 212.139
R2287 avdd_ip.n90 avdd_ip.n89 202.696
R2288 avdd_ip.n88 avdd_ip.n29 134.065
R2289 avdd_ip.n74 avdd_ip.n29 110.358
R2290 avdd_ip.t6 avdd_ip.n26 105.665
R2291 avdd_ip.t10 avdd_ip.n27 105.665
R2292 avdd_ip.n85 avdd_ip.n84 96.3051
R2293 avdd_ip.n58 avdd_ip.n57 92.5005
R2294 avdd_ip.n55 avdd_ip.n49 92.5005
R2295 avdd_ip.n54 avdd_ip.n53 92.5005
R2296 avdd_ip.n52 avdd_ip.n50 92.5005
R2297 avdd_ip.n45 avdd_ip.n44 92.5005
R2298 avdd_ip.n44 avdd_ip.n43 92.5005
R2299 avdd_ip.n38 avdd_ip.n37 92.5005
R2300 avdd_ip.t2 avdd_ip.n37 92.5005
R2301 avdd_ip.n40 avdd_ip.n39 92.5005
R2302 avdd_ip.n36 avdd_ip.n35 92.5005
R2303 avdd_ip.n39 avdd_ip.n35 91.4862
R2304 avdd_ip.n53 avdd_ip.n49 91.4829
R2305 avdd_ip.n92 avdd_ip.t6 79.5673
R2306 avdd_ip.n92 avdd_ip.t10 79.5673
R2307 avdd_ip.n85 avdd_ip.n62 73.3959
R2308 avdd_ip.n39 avdd_ip.n38 66.8321
R2309 avdd_ip.n53 avdd_ip.n52 66.3131
R2310 avdd_ip.n59 avdd_ip.n49 63.936
R2311 avdd_ip.n46 avdd_ip.n35 63.936
R2312 avdd_ip.n2 avdd_ip.t1 62.0945
R2313 avdd_ip.n17 avdd_ip.t23 61.1041
R2314 avdd_ip.n15 avdd_ip.t24 60.1061
R2315 avdd_ip.n14 avdd_ip.t20 60.1061
R2316 avdd_ip.n21 avdd_ip.t21 60.1061
R2317 avdd_ip.n24 avdd_ip.t19 60.1061
R2318 avdd_ip.n89 avdd_ip.t14 60.1061
R2319 avdd_ip.n89 avdd_ip.t11 60.1061
R2320 avdd_ip.n89 avdd_ip.t12 60.1061
R2321 avdd_ip.n63 avdd_ip.t9 60.1061
R2322 avdd_ip.n63 avdd_ip.t7 60.1061
R2323 avdd_ip.n63 avdd_ip.t8 60.1061
R2324 avdd_ip.n31 avdd_ip.t15 60.1061
R2325 avdd_ip.n31 avdd_ip.t13 60.1061
R2326 avdd_ip.n30 avdd_ip.t17 60.1061
R2327 avdd_ip.n30 avdd_ip.t16 60.1061
R2328 avdd_ip.n65 avdd_ip.t26 60.1061
R2329 avdd_ip.n65 avdd_ip.t18 60.1061
R2330 avdd_ip.n64 avdd_ip.t27 60.1061
R2331 avdd_ip.n64 avdd_ip.t22 60.1061
R2332 avdd_ip.n16 avdd_ip.t25 60.1061
R2333 avdd_ip.n41 avdd_ip.n36 57.4849
R2334 avdd_ip.n56 avdd_ip.n55 57.4849
R2335 avdd_ip.n51 avdd_ip.n50 57.4849
R2336 avdd_ip.n2 avdd_ip.n1 55.1707
R2337 avdd_ip.n2 avdd_ip.n0 54.9038
R2338 avdd_ip.n69 avdd_ip.n13 44.6614
R2339 avdd_ip.n58 avdd_ip.n48 43.3376
R2340 avdd_ip.n45 avdd_ip.n34 43.3376
R2341 avdd_ip.n83 avdd_ip.n70 30.1747
R2342 avdd_ip.n51 avdd_ip.t5 28.8172
R2343 avdd_ip.n56 avdd_ip.t5 28.8172
R2344 avdd_ip.t2 avdd_ip.n41 28.8172
R2345 avdd_ip.n90 avdd_ip.n28 10.6324
R2346 avdd_ip.n74 avdd_ip.n25 8.37369
R2347 avdd_ip.n16 avdd_ip.n15 7.25561
R2348 avdd_ip.n0 avdd_ip.t3 6.92425
R2349 avdd_ip.n0 avdd_ip.t0 6.92425
R2350 avdd_ip.n1 avdd_ip.t28 6.92425
R2351 avdd_ip.n1 avdd_ip.t4 6.92425
R2352 avdd_ip.n91 avdd_ip.n90 6.37981
R2353 avdd_ip.n92 avdd_ip.n91 6.37981
R2354 avdd_ip.n94 avdd_ip.n93 6.37981
R2355 avdd_ip.n93 avdd_ip.n92 6.37981
R2356 avdd_ip.n24 avdd_ip.n23 6.17839
R2357 avdd_ip.n78 avdd_ip.n77 6.15262
R2358 avdd_ip.n94 avdd_ip.n25 5.31953
R2359 avdd_ip.n52 avdd_ip.n48 4.38907
R2360 avdd_ip.n38 avdd_ip.n34 4.38907
R2361 avdd_ip.n95 avdd_ip.n94 3.87825
R2362 avdd_ip.n84 avdd_ip.n83 3.6009
R2363 avdd_ip.n60 avdd_ip.n48 2.4925
R2364 avdd_ip.n47 avdd_ip.n34 2.44611
R2365 avdd_ip.n29 avdd_ip.n27 2.43471
R2366 avdd_ip.n70 avdd_ip.n26 2.43471
R2367 avdd_ip.n59 avdd_ip.n58 2.37764
R2368 avdd_ip.n46 avdd_ip.n45 2.37764
R2369 avdd_ip.n60 avdd_ip.n59 2.3255
R2370 avdd_ip.n47 avdd_ip.n46 2.3255
R2371 avdd_ip.n22 avdd_ip.n21 1.87566
R2372 avdd_ip.n95 avdd_ip.n13 1.41891
R2373 avdd_ip.n4 avdd_ip.n3 1.18871
R2374 avdd_ip.n23 avdd_ip.n14 1.07773
R2375 avdd_ip.n79 avdd_ip.n78 1.05764
R2376 avdd_ip.n83 avdd_ip.n82 1.05764
R2377 avdd_ip.n82 avdd_ip.n81 1.05764
R2378 avdd_ip.n86 avdd_ip.n85 1.02375
R2379 avdd_ip.n21 avdd_ip.n20 0.982678
R2380 avdd_ip.n20 avdd_ip.n14 0.919312
R2381 avdd_ip.n17 avdd_ip.n16 0.90347
R2382 avdd_ip.n23 avdd_ip.n22 0.845955
R2383 avdd_ip.n11 avdd_ip.n4 0.827286
R2384 avdd_ip avdd_ip.n11 0.808179
R2385 avdd_ip.n66 avdd_ip.n64 0.65712
R2386 avdd_ip.n32 avdd_ip.n30 0.652725
R2387 avdd_ip.n88 avdd_ip.n87 0.613954
R2388 avdd_ip.n76 avdd_ip.n72 0.530586
R2389 avdd_ip.n80 avdd_ip.n72 0.530586
R2390 avdd_ip.n75 avdd_ip.n71 0.530586
R2391 avdd_ip.n73 avdd_ip.n71 0.530586
R2392 avdd_ip.n3 avdd_ip.n2 0.507794
R2393 avdd_ip.n70 avdd_ip.n69 0.448948
R2394 avdd_ip.n19 avdd_ip.n18 0.402976
R2395 avdd_ip.n33 avdd_ip.n32 0.319749
R2396 avdd_ip.n87 avdd_ip.n86 0.319015
R2397 avdd_ip.n67 avdd_ip.n66 0.319015
R2398 avdd_ip.n18 avdd_ip.n12 0.319015
R2399 avdd_ip.n20 avdd_ip.n19 0.282318
R2400 avdd_ip.n11 avdd_ip.n10 0.255087
R2401 avdd_ip.n32 avdd_ip.n31 0.25137
R2402 avdd_ip.n66 avdd_ip.n65 0.25137
R2403 avdd_ip.n96 avdd_ip.n12 0.243945
R2404 avdd_ip avdd_ip.n97 0.213307
R2405 avdd_ip.n87 avdd_ip.n28 0.211864
R2406 avdd_ip.n18 avdd_ip.n17 0.211864
R2407 avdd_ip.n97 avdd_ip 0.18211
R2408 avdd_ip.n25 avdd_ip.n24 0.174542
R2409 avdd_ip.n15 avdd_ip.n13 0.174542
R2410 avdd_ip.n62 avdd_ip.n61 0.166571
R2411 avdd_ip.n67 avdd_ip.n12 0.150396
R2412 avdd_ip.n86 avdd_ip.n33 0.150396
R2413 avdd_ip.n3 avdd_ip.t33 0.125045
R2414 avdd_ip.n7 avdd_ip.n4 0.123905
R2415 avdd_ip.n68 avdd_ip.n33 0.117461
R2416 avdd_ip.n10 avdd_ip.n9 0.111971
R2417 avdd_ip.n8 avdd_ip.n7 0.110265
R2418 avdd_ip.n68 avdd_ip.n67 0.108384
R2419 avdd_ip.n6 avdd_ip.n5 0.106696
R2420 avdd_ip.n9 avdd_ip.n8 0.106696
R2421 avdd_ip.n61 avdd_ip.n47 0.0839309
R2422 avdd_ip.n61 avdd_ip.n60 0.0812962
R2423 avdd_ip.n5 avdd_ip.t30 0.0180781
R2424 avdd_ip.n9 avdd_ip.t32 0.0180781
R2425 avdd_ip.n8 avdd_ip.t29 0.0180781
R2426 avdd_ip.n6 avdd_ip.t31 0.0180781
R2427 avdd_ip.n10 avdd_ip.n5 0.0174228
R2428 avdd_ip.n96 avdd_ip.n95 0.0173478
R2429 avdd_ip.n63 avdd_ip.n28 0.0154184
R2430 avdd_ip.n89 avdd_ip.n88 0.0154184
R2431 avdd_ip.n7 avdd_ip.n6 0.0150053
R2432 avdd_ip.n69 avdd_ip.n68 0.0108333
R2433 avdd_ip.n97 avdd_ip.n96 0.00292843
R2434 avdd_ip.n22 avdd_ip.n19 0.000885802
R2435 xout.n29 xout.t26 594.784
R2436 xout.n29 xout.t24 194.649
R2437 xout.n25 xout.t23 124.457
R2438 xout.n25 xout.t25 106.793
R2439 xout.t23 xout.n24 86.3125
R2440 xout.t25 xout.n23 86.3125
R2441 xout.n3 xout.t14 62.0071
R2442 xout.n4 xout.t12 62.0071
R2443 xout.n3 xout.t19 60.1061
R2444 xout.n4 xout.t20 60.1061
R2445 xout.n8 xout.t10 60.1061
R2446 xout.n8 xout.t9 60.1061
R2447 xout.n10 xout.t13 60.1061
R2448 xout.n10 xout.t11 60.1061
R2449 xout.n0 xout.t16 60.1061
R2450 xout.n0 xout.t18 60.1061
R2451 xout.n1 xout.t15 60.1061
R2452 xout.n1 xout.t17 60.1061
R2453 xout.n24 xout.n23 58.6245
R2454 xout.n22 xout.t7 43.5339
R2455 xout.n28 xout.n27 21.3269
R2456 xout.n16 xout.n15 18.5533
R2457 xout.n20 xout.n13 18.553
R2458 xout.n19 xout.n18 18.4723
R2459 xout.n19 xout.n17 18.4564
R2460 xout.n16 xout.n14 18.4564
R2461 xout.n27 xout.n23 12.2455
R2462 xout.n18 xout.t4 4.133
R2463 xout.n18 xout.t2 4.133
R2464 xout.n17 xout.t6 4.133
R2465 xout.n17 xout.t5 4.133
R2466 xout.n15 xout.t21 4.133
R2467 xout.n15 xout.t8 4.133
R2468 xout.n14 xout.t3 4.133
R2469 xout.n14 xout.t0 4.133
R2470 xout.n13 xout.t1 4.133
R2471 xout.n13 xout.t22 4.133
R2472 xout.n5 xout.n4 3.64406
R2473 xout.n5 xout.n3 3.61238
R2474 xout.n26 xout.n24 3.56553
R2475 xout.n22 xout.n21 2.24362
R2476 xout.n29 xout.n28 2.18092
R2477 xout.n28 xout.n22 1.03102
R2478 xout.n27 xout.n26 0.742745
R2479 xout.n26 xout.n25 0.715885
R2480 xout.n21 xout.n12 0.464586
R2481 xout.n2 xout.n0 0.424187
R2482 xout.n11 xout.n9 0.402558
R2483 xout xout.n29 0.377063
R2484 xout.n6 xout.n2 0.316998
R2485 xout.n2 xout.n1 0.310571
R2486 xout.n12 xout.n7 0.273717
R2487 xout.n7 xout.n6 0.261913
R2488 xout.n9 xout.n8 0.254998
R2489 xout.n11 xout.n10 0.25137
R2490 xout.n6 xout.n5 0.143668
R2491 xout.n9 xout.n7 0.126918
R2492 xout.n12 xout.n11 0.125886
R2493 xout.n21 xout.n20 0.0947164
R2494 xout.n20 xout.n16 0.0657574
R2495 xout.n20 xout.n19 0.0480746
R2496 inv_in.n19 inv_in.t0 47.4896
R2497 inv_in.n18 inv_in.t3 6.48745
R2498 inv_in.n19 inv_in.t1 6.24255
R2499 inv_in inv_in.n17 2.2182
R2500 inv_in.n18 inv_in 0.342687
R2501 inv_in inv_in.n18 0.217687
R2502 inv_in.n5 inv_in.n4 0.110198
R2503 inv_in.n7 inv_in.n6 0.110101
R2504 inv_in.n10 inv_in.n9 0.110101
R2505 inv_in.n8 inv_in.n2 0.110101
R2506 inv_in.n16 inv_in.n15 0.109734
R2507 inv_in.n14 inv_in.n0 0.109734
R2508 inv_in.n13 inv_in.n12 0.109709
R2509 inv_in.n11 inv_in.n1 0.109709
R2510 inv_in.n9 inv_in.n7 0.109325
R2511 inv_in.n9 inv_in.n8 0.109325
R2512 inv_in.n12 inv_in.n11 0.109325
R2513 inv_in.n11 inv_in.n3 0.109325
R2514 inv_in.n15 inv_in.n14 0.1086
R2515 inv_in.n16 inv_in.n0 0.1086
R2516 inv_in.n4 inv_in.n3 0.10222
R2517 inv_in.n7 inv_in.n5 0.101755
R2518 inv_in inv_in.n19 0.09425
R2519 inv_in.n18 inv_in 0.063
R2520 inv_in.n0 inv_in.t11 0.00880157
R2521 inv_in.n7 inv_in.t9 0.00848368
R2522 inv_in.n9 inv_in.t10 0.00848368
R2523 inv_in.n8 inv_in.t2 0.00848368
R2524 inv_in.n5 inv_in.t12 0.00838586
R2525 inv_in.n4 inv_in.t14 0.0083125
R2526 inv_in.n6 inv_in.t13 0.0083125
R2527 inv_in.n2 inv_in.t6 0.0083125
R2528 inv_in.n10 inv_in.t4 0.0083125
R2529 inv_in.n1 inv_in.t5 0.0083125
R2530 inv_in.n13 inv_in.t8 0.0083125
R2531 inv_in.n17 inv_in.t7 0.0083125
R2532 inv_in.n6 inv_in.n3 0.00106244
R2533 inv_in.n12 inv_in.n2 0.00106244
R2534 inv_in.n11 inv_in.n10 0.00106244
R2535 inv_in.n17 inv_in.n16 0.000989074
R2536 inv_in.n15 inv_in.n1 0.000548907
R2537 inv_in.n14 inv_in.n13 0.000548907
R2538 dout_ip.n0 dout_ip.t2 651.692
R2539 dout_ip.n0 dout_ip.t3 651.431
R2540 dout_ip.n1 dout_ip.t9 288.204
R2541 dout_ip.n5 dout_ip.t5 264.103
R2542 dout_ip.n2 dout_ip.t6 264.103
R2543 dout_ip.n0 dout_ip.t1 229.352
R2544 dout_ip.n0 dout_ip.t0 229.101
R2545 dout_ip.n1 dout_ip.t7 195.017
R2546 x7.x2.clkin dout_ip.n5 159.236
R2547 x7.x1.clkin dout_ip.n2 159.236
R2548 x7.x5.A dout_ip.n1 153.153
R2549 dout_ip.n4 x7.x2.x1.A 152
R2550 x7.x1.x1.A dout_ip.n3 152
R2551 dout_ip.n4 dout_ip.t8 145.209
R2552 dout_ip.n3 dout_ip.t4 145.209
R2553 dout_ip.n7 dout_ip.n6 117.519
R2554 dout_ip.n6 x7.x1.clkin 68.1959
R2555 dout_ip.n5 dout_ip.n4 37.6741
R2556 dout_ip.n3 dout_ip.n2 37.6741
R2557 x7.clkin dout_ip.n7 31.6505
R2558 dout_ip.n7 x7.x5.A 24.4485
R2559 x7.clkin dout_ip.n0 11.4719
R2560 x7.x2.clkin x7.x2.x1.A 10.3444
R2561 x7.x1.clkin x7.x1.x1.A 10.3444
R2562 dout_ip.n6 x7.x2.clkin 9.3005
R2563 avss.n20 avss.n19 18580.7
R2564 avss.n38 avss.n37 15308.7
R2565 avss.n76 avss.n20 12246.6
R2566 avss.n40 avss.n35 3599.36
R2567 avss.n41 avss.n35 3599.36
R2568 avss.n41 avss.n34 3599.36
R2569 avss.n40 avss.n34 3599.36
R2570 avss.n67 avss.n25 2489.59
R2571 avss.n67 avss.n26 2489.59
R2572 avss.n69 avss.n26 2489.59
R2573 avss.n69 avss.n25 2489.59
R2574 avss.n28 avss.n21 2489.59
R2575 avss.n28 avss.n22 2489.59
R2576 avss.n74 avss.n22 2489.59
R2577 avss.n74 avss.n21 2489.59
R2578 avss.n78 avss.n13 2489.59
R2579 avss.n78 avss.n14 2489.59
R2580 avss.n16 avss.n14 2489.59
R2581 avss.n16 avss.n13 2489.59
R2582 avss.n88 avss.n6 2489.59
R2583 avss.n90 avss.n6 2489.59
R2584 avss.n90 avss.n5 2489.59
R2585 avss.n88 avss.n5 2489.59
R2586 avss.n36 avss.n20 2342.14
R2587 avss.n77 avss.n76 930.542
R2588 avss.n76 avss.n75 930.542
R2589 avss.n43 avss.n42 881.42
R2590 avss.n19 avss.t16 633.244
R2591 avss.n15 avss.t14 633.244
R2592 avss.t0 avss.n17 633.244
R2593 avss.n77 avss.t2 633.244
R2594 avss.n75 avss.t4 633.244
R2595 avss.n29 avss.t6 633.244
R2596 avss.t20 avss.n30 633.244
R2597 avss.n37 avss.t22 633.244
R2598 avss.t12 avss.n36 412.863
R2599 avss.t10 avss.n38 397.358
R2600 avss.n17 avss.n15 362.704
R2601 avss.n30 avss.n29 362.704
R2602 avss.t8 avss.t12 306.255
R2603 avss.t24 avss.t8 306.255
R2604 avss.t24 avss.t18 306.255
R2605 avss.t18 avss.t10 306.255
R2606 avss.n39 avss.n32 295.807
R2607 avss.n66 avss.n65 289.13
R2608 avss.n87 avss.n3 289.13
R2609 avss.n92 avss.n91 288.753
R2610 avss.n70 avss.n24 288.753
R2611 avss.n89 avss.t16 234.865
R2612 avss.n89 avss.t14 234.865
R2613 avss.n18 avss.t0 234.865
R2614 avss.t2 avss.n18 234.865
R2615 avss.n27 avss.t4 234.865
R2616 avss.t6 avss.n27 234.865
R2617 avss.n68 avss.t20 234.865
R2618 avss.n68 avss.t22 234.865
R2619 avss.n31 avss.n10 152.73
R2620 avss.n73 avss.n72 152.73
R2621 avss.n80 avss.n7 152.73
R2622 avss.n79 avss.n12 152.73
R2623 avss.n39 avss.n33 118.081
R2624 avss.n91 avss.n4 103.529
R2625 avss.n64 avss.n31 103.529
R2626 avss.n72 avss.n71 103.529
R2627 avss.n66 avss.n64 103.529
R2628 avss.n71 avss.n70 103.529
R2629 avss.n86 avss.n7 103.529
R2630 avss.n12 avss.n4 103.529
R2631 avss.n87 avss.n86 103.529
R2632 avss.n88 avss.n87 97.5005
R2633 avss.n89 avss.n88 97.5005
R2634 avss.n91 avss.n90 97.5005
R2635 avss.n90 avss.n89 97.5005
R2636 avss.n13 avss.n7 97.5005
R2637 avss.n18 avss.n13 97.5005
R2638 avss.n14 avss.n12 97.5005
R2639 avss.n18 avss.n14 97.5005
R2640 avss.n31 avss.n21 97.5005
R2641 avss.n27 avss.n21 97.5005
R2642 avss.n72 avss.n22 97.5005
R2643 avss.n27 avss.n22 97.5005
R2644 avss.n70 avss.n69 97.5005
R2645 avss.n69 avss.n68 97.5005
R2646 avss.n67 avss.n66 97.5005
R2647 avss.n68 avss.n67 97.5005
R2648 avss.n42 avss.n33 69.8003
R2649 avss.n38 avss.n35 54.5071
R2650 avss.n5 avss.n3 48.7505
R2651 avss.n19 avss.n5 48.7505
R2652 avss.n8 avss.n6 48.7505
R2653 avss.n15 avss.n6 48.7505
R2654 avss.n16 avss.n8 48.7505
R2655 avss.n17 avss.n16 48.7505
R2656 avss.n79 avss.n78 48.7505
R2657 avss.n78 avss.n77 48.7505
R2658 avss.n74 avss.n73 48.7505
R2659 avss.n75 avss.n74 48.7505
R2660 avss.n28 avss.n23 48.7505
R2661 avss.n29 avss.n28 48.7505
R2662 avss.n25 avss.n23 48.7505
R2663 avss.n30 avss.n25 48.7505
R2664 avss.n65 avss.n26 48.7505
R2665 avss.n37 avss.n26 48.7505
R2666 avss.n40 avss.n39 45.0005
R2667 avss.t24 avss.n40 45.0005
R2668 avss.n42 avss.n41 45.0005
R2669 avss.n41 avss.t24 45.0005
R2670 avss.n64 avss.n63 40.3697
R2671 avss.n71 avss.n23 40.3697
R2672 avss.n86 avss.n85 40.3697
R2673 avss.n8 avss.n4 40.3697
R2674 avss.n94 avss.n1 39.7977
R2675 avss.n34 avss.n33 39.0005
R2676 avss.n36 avss.n34 39.0005
R2677 avss.n35 avss.n32 39.0005
R2678 avss.n94 avss 33.7505
R2679 avss.n84 avss.t1 29.9199
R2680 avss.n62 avss.t21 29.9199
R2681 avss.n62 avss.t7 29.9199
R2682 avss.n84 avss.t15 29.9199
R2683 avss.n2 avss.t17 29.798
R2684 avss.n57 avss.t23 29.798
R2685 avss.n11 avss.t3 29.798
R2686 avss.n11 avss.t5 29.798
R2687 avss.n32 avss.t11 20.9512
R2688 avss.n46 avss.n45 18.8362
R2689 avss.n46 avss.n44 18.6458
R2690 avss.n44 avss.t25 4.133
R2691 avss.n44 avss.t19 4.133
R2692 avss.n45 avss.t13 4.133
R2693 avss.n45 avss.t9 4.133
R2694 avss.n47 avss.n43 1.61679
R2695 avss.n55 avss 1.33946
R2696 avss.n58 avss.n24 1.21803
R2697 avss.n93 avss.n92 1.21803
R2698 avss.n54 avss.n47 0.8655
R2699 avss.n63 avss.n62 0.664786
R2700 avss.n81 avss.n10 0.664786
R2701 avss.n81 avss.n80 0.664786
R2702 avss.n85 avss.n84 0.664786
R2703 avss.n55 avss.n54 0.53175
R2704 avss.n56 avss.n9 0.434977
R2705 avss.n95 avss.n0 0.433066
R2706 avss.n61 avss.n59 0.433066
R2707 avss.n61 avss.n60 0.433066
R2708 avss.n60 avss.n0 0.433066
R2709 avss.n65 avss.n24 0.376971
R2710 avss.n92 avss.n3 0.376971
R2711 avss.n84 avss.n0 0.299413
R2712 avss.n62 avss.n61 0.299413
R2713 avss.n62 avss.n9 0.247783
R2714 avss.n84 avss.n83 0.247783
R2715 avss.n83 avss 0.245943
R2716 avss.n59 avss.n58 0.231236
R2717 avss.n82 avss.n9 0.201672
R2718 avss.n83 avss.n82 0.201672
R2719 avss.n2 avss.n1 0.2005
R2720 avss.n95 avss.n94 0.2005
R2721 avss.n47 avss.n46 0.1855
R2722 avss.n49 avss.n48 0.122162
R2723 avss.n82 avss.n81 0.120904
R2724 avss.n50 avss.n49 0.105544
R2725 avss.n51 avss.n50 0.101695
R2726 avss.n73 avss.n10 0.1005
R2727 avss.n80 avss.n79 0.1005
R2728 avss.n60 avss.n11 0.0997647
R2729 avss.n53 avss.n48 0.0989292
R2730 avss.n56 avss.n55 0.096886
R2731 avss.n54 avss.n53 0.0847138
R2732 avss.n63 avss.n23 0.0825513
R2733 avss.n85 avss.n8 0.0825513
R2734 avss.n51 avss.n48 0.0586846
R2735 avss.n57 avss.n56 0.0480171
R2736 avss avss.n95 0.0332586
R2737 avss.n59 avss 0.0330342
R2738 avss.n94 avss.n93 0.0328276
R2739 avss.n43 avss.n32 0.0328232
R2740 avss.n53 avss.n52 0.0277801
R2741 avss.n50 avss.t28 0.0083125
R2742 avss.n49 avss.t29 0.0083125
R2743 avss.n48 avss.t26 0.0083125
R2744 avss.n52 avss.t27 0.0083125
R2745 avss avss.n1 0.00342969
R2746 avss.n93 avss.n2 0.000931034
R2747 avss.n58 avss.n57 0.000928082
R2748 avss.n81 avss.n11 0.000683824
R2749 avss.n52 avss.n51 0.000622332
R2750 avdd.n92 avdd.n91 15807.9
R2751 avdd.n93 avdd.n92 15807.9
R2752 avdd.n93 avdd.n28 15807.9
R2753 avdd.n91 avdd.n28 15807.9
R2754 avdd.n90 avdd.n27 8112.97
R2755 avdd.n94 avdd.n27 8112.97
R2756 avdd.n94 avdd.n26 8112.97
R2757 avdd.n90 avdd.n26 8112.97
R2758 avdd.n98 avdd.n6 2166
R2759 avdd.n97 avdd.n6 2166
R2760 avdd.n98 avdd.n7 2166
R2761 avdd.n97 avdd.n7 2166
R2762 avdd.n78 avdd.n77 1643.17
R2763 avdd.n77 avdd.n76 1643.17
R2764 avdd.n74 avdd.n69 1643.17
R2765 avdd.n80 avdd.n69 1643.17
R2766 avdd.n52 avdd.n37 1643.17
R2767 avdd.n60 avdd.n37 1643.17
R2768 avdd.n55 avdd.n54 1643.17
R2769 avdd.n58 avdd.n55 1643.17
R2770 avdd.n89 avdd.n88 1439.4
R2771 avdd.n89 avdd.n29 1352.37
R2772 avdd.n66 avdd.n25 1313.54
R2773 avdd.n71 avdd.n70 1106.59
R2774 avdd.n70 avdd.n68 1106.59
R2775 avdd.n40 avdd.n39 1106.59
R2776 avdd.n39 avdd.n36 1106.59
R2777 avdd.n78 avdd.n68 536.587
R2778 avdd.n76 avdd.n71 536.587
R2779 avdd.n74 avdd.n71 536.587
R2780 avdd.n80 avdd.n68 536.587
R2781 avdd.n52 avdd.n40 536.587
R2782 avdd.n54 avdd.n40 536.587
R2783 avdd.n58 avdd.n36 536.587
R2784 avdd.n60 avdd.n36 536.587
R2785 avdd.n75 avdd.t6 382.582
R2786 avdd.n79 avdd.t6 382.582
R2787 avdd.n53 avdd.t2 382.582
R2788 avdd.n59 avdd.t2 382.582
R2789 avdd.n73 avdd.n30 319.248
R2790 avdd.n57 avdd.n56 319.248
R2791 avdd.n88 avdd.n31 287.265
R2792 avdd.n38 avdd.n29 287.265
R2793 avdd.n88 avdd.n30 276.295
R2794 avdd.n56 avdd.n29 276.295
R2795 avdd.n86 avdd.t7 227.377
R2796 avdd.n1 avdd.t19 227.377
R2797 avdd.n34 avdd.t3 227.377
R2798 avdd.n43 avdd.t8 227.377
R2799 avdd.n66 avdd.n3 205.554
R2800 avdd.n72 avdd.n31 189.742
R2801 avdd.n38 avdd.n35 189.742
R2802 avdd.n101 avdd.n3 186.73
R2803 avdd.t17 avdd.n6 157.492
R2804 avdd.t4 avdd.n7 157.492
R2805 avdd.n25 avdd.n4 118.862
R2806 avdd.n100 avdd.n4 115.031
R2807 avdd.n73 avdd.n72 108.569
R2808 avdd.n57 avdd.n35 108.569
R2809 avdd.t11 avdd.t17 107.677
R2810 avdd.t9 avdd.t11 107.677
R2811 avdd.t9 avdd.t0 107.677
R2812 avdd.t0 avdd.t4 107.677
R2813 avdd.n62 avdd.n5 63.4672
R2814 avdd.n23 avdd.t18 60.1061
R2815 avdd.n21 avdd.n20 54.9038
R2816 avdd.n21 avdd.n19 54.9038
R2817 avdd.n72 avdd.n2 32.2138
R2818 avdd.n61 avdd.n35 32.2138
R2819 avdd.n101 avdd.n100 31.7005
R2820 avdd.n102 avdd.n101 30.3938
R2821 avdd.n76 avdd.n73 26.4291
R2822 avdd.n76 avdd.n75 26.4291
R2823 avdd.n74 avdd.n2 26.4291
R2824 avdd.n75 avdd.n74 26.4291
R2825 avdd.n78 avdd.n32 26.4291
R2826 avdd.n79 avdd.n78 26.4291
R2827 avdd.n81 avdd.n80 26.4291
R2828 avdd.n80 avdd.n79 26.4291
R2829 avdd.n58 avdd.n57 26.4291
R2830 avdd.n59 avdd.n58 26.4291
R2831 avdd.n61 avdd.n60 26.4291
R2832 avdd.n60 avdd.n59 26.4291
R2833 avdd.n54 avdd.n41 26.4291
R2834 avdd.n54 avdd.n53 26.4291
R2835 avdd.n52 avdd.n51 26.4291
R2836 avdd.n53 avdd.n52 26.4291
R2837 avdd.n96 avdd.n24 15.6997
R2838 avdd.n97 avdd.n96 14.2313
R2839 avdd.t9 avdd.n97 14.2313
R2840 avdd.n99 avdd.n98 14.2313
R2841 avdd.n98 avdd.t9 14.2313
R2842 avdd.n77 avdd.n30 13.2148
R2843 avdd.n77 avdd.t6 13.2148
R2844 avdd.n70 avdd.n31 13.2148
R2845 avdd.n70 avdd.t6 13.2148
R2846 avdd.n69 avdd.n3 13.2148
R2847 avdd.t6 avdd.n69 13.2148
R2848 avdd.n39 avdd.n38 13.2148
R2849 avdd.n39 avdd.t2 13.2148
R2850 avdd.n56 avdd.n55 13.2148
R2851 avdd.n55 avdd.t2 13.2148
R2852 avdd.n49 avdd.n37 13.2148
R2853 avdd.t2 avdd.n37 13.2148
R2854 avdd.n7 avdd.n4 12.3338
R2855 avdd.n47 avdd.n6 12.3338
R2856 avdd.n100 avdd.n99 8.13132
R2857 avdd.n95 avdd.n25 7.54184
R2858 avdd.n82 avdd.n32 7.30037
R2859 avdd.n46 avdd.n41 7.22016
R2860 avdd.n20 avdd.t12 6.92425
R2861 avdd.n20 avdd.t10 6.92425
R2862 avdd.n19 avdd.t1 6.92425
R2863 avdd.n19 avdd.t5 6.92425
R2864 avdd.n48 avdd.n47 6.88003
R2865 avdd.n99 avdd.n5 6.16704
R2866 avdd.n67 avdd.n66 3.51587
R2867 avdd.n50 avdd.n49 3.30818
R2868 avdd.n82 avdd.n81 2.8599
R2869 avdd.n90 avdd.n89 2.84665
R2870 avdd.n91 avdd.n90 2.84665
R2871 avdd.n95 avdd.n94 2.84665
R2872 avdd.n94 avdd.n93 2.84665
R2873 avdd.n51 avdd.n46 2.78239
R2874 avdd.n48 avdd.n5 2.51338
R2875 avdd.n49 avdd.n48 2.33395
R2876 avdd.n67 avdd.n27 2.28445
R2877 avdd.n92 avdd.n27 2.28445
R2878 avdd.n50 avdd.n26 2.28445
R2879 avdd.n28 avdd.n26 2.28445
R2880 avdd.n84 avdd 1.89829
R2881 avdd.n23 avdd.n22 1.87575
R2882 avdd.n102 avdd.n2 1.70717
R2883 avdd.n62 avdd.n61 1.70717
R2884 avdd.n81 avdd.n67 1.56476
R2885 avdd.n51 avdd.n50 1.54047
R2886 avdd.n85 avdd.n1 1.11161
R2887 avdd.n96 avdd.n95 1.03878
R2888 avdd.n65 avdd.n33 0.909856
R2889 avdd.n87 avdd.n65 0.871595
R2890 avdd.n42 avdd.n29 0.517167
R2891 avdd.n63 avdd.n62 0.517167
R2892 avdd.n103 avdd.n102 0.517167
R2893 avdd.n88 avdd.n87 0.517167
R2894 avdd.n83 avdd.n1 0.457832
R2895 avdd.n88 avdd.n32 0.30326
R2896 avdd.n41 avdd.n29 0.29856
R2897 avdd.n44 avdd.n34 0.277965
R2898 avdd.n44 avdd.n43 0.242141
R2899 avdd.n13 avdd.n12 0.221624
R2900 avdd.n45 avdd.n44 0.191202
R2901 avdd.n15 avdd.n8 0.171
R2902 avdd.n64 avdd 0.165618
R2903 avdd.n18 avdd.n8 0.158572
R2904 avdd.n45 avdd.n33 0.155105
R2905 avdd.n22 avdd.n18 0.129984
R2906 avdd.n65 avdd.n64 0.124867
R2907 avdd.n24 avdd.n23 0.0960224
R2908 avdd.n18 avdd.n17 0.0860931
R2909 avdd.n16 avdd.n15 0.0718577
R2910 avdd.n15 avdd.n14 0.0677409
R2911 avdd.n46 avdd.n45 0.058264
R2912 avdd.n83 avdd.n82 0.058264
R2913 avdd.n86 avdd.n85 0.0482015
R2914 avdd avdd.n63 0.0421667
R2915 avdd avdd.n0 0.035342
R2916 avdd.n12 avdd.n0 0.0293462
R2917 avdd.n22 avdd.n21 0.0285269
R2918 avdd.n17 avdd.n16 0.0255438
R2919 avdd.n14 avdd.n13 0.0253723
R2920 avdd.n12 avdd.n8 0.0246031
R2921 avdd.n85 avdd.n84 0.0240664
R2922 avdd.n11 avdd.t15 0.0122401
R2923 avdd avdd.n103 0.0122337
R2924 avdd.n17 avdd.t13 0.0122173
R2925 avdd.n10 avdd.t16 0.0113908
R2926 avdd.n9 avdd.t14 0.011362
R2927 avdd.n63 avdd.n34 0.0105575
R2928 avdd.n103 avdd.n1 0.0105575
R2929 avdd.n17 avdd.n9 0.00991802
R2930 avdd.n11 avdd.n10 0.00930403
R2931 avdd.n47 avdd.n24 0.00805162
R2932 avdd.n64 avdd 0.00600766
R2933 avdd.n43 avdd.n42 0.00573256
R2934 avdd.n42 avdd.n33 0.00515116
R2935 avdd.n87 avdd.n86 0.00333375
R2936 avdd.n14 avdd.n9 0.00220261
R2937 avdd.n16 avdd.n10 0.00176706
R2938 avdd.n84 avdd.n83 0.00111075
R2939 avdd.n64 avdd.n0 0.00109866
R2940 avdd.n13 avdd.n11 0.000671533
R2941 standby.n1 standby.t0 260.322
R2942 standby.n0 standby.t1 194.635
R2943 standby.n1 standby.t2 175.169
R2944 standby.n2 standby.n1 152
R2945 standby.n2 standby.n0 69.674
R2946 standby standby.n2 1.55726
R2947 standby.n0 standby 0.748625
R2948 x3.out_b.n5 x3.out_b.t8 397.163
R2949 x3.out_b.n3 x3.out_b.t4 397.163
R2950 x3.out_b.n6 x3.out_b.t8 396.286
R2951 x3.out_b.n4 x3.out_b.t4 396.286
R2952 x3.out_b.t3 x3.out_b.n5 375.649
R2953 x3.out_b.n6 x3.out_b.t3 375.649
R2954 x3.out_b.n0 x3.out_b.t6 375.649
R2955 x3.out_b.n7 x3.out_b.t6 375.649
R2956 x3.out_b.t7 x3.out_b.n3 375.649
R2957 x3.out_b.n4 x3.out_b.t7 375.649
R2958 x3.out_b.n2 x3.out_b.t2 227.887
R2959 x3.out_b.n2 x3.out_b.n8 25.0905
R2960 x3.out_b.n5 x3.out_b.n0 21.5154
R2961 x3.out_b.n3 x3.out_b.n0 21.1069
R2962 x3.out_b.n7 x3.out_b.n4 20.6372
R2963 x3.out_b.n7 x3.out_b.n6 20.6372
R2964 x3.out_b.n2 x3.out_b.t5 12.777
R2965 x3.out_b.n8 x3.out_b.t0 5.5105
R2966 x3.out_b.n8 x3.out_b.t1 5.5105
R2967 x3.out_b.n1 x3.out_b.n0 5.32901
R2968 x3.out_b.n1 x3.out_b.n7 2.74252
R2969 x3.out_b.n2 x3.out_b.n1 1.06508
R2970 ena.n0 ena.t2 260.322
R2971 ena.n2 ena.t0 194.63
R2972 ena.n0 ena.t1 175.169
R2973 ena.n1 ena.n0 152
R2974 ena.n3 ena.n2 51.6747
R2975 ena ena.n3 4.94983
R2976 ena.n3 ena.n1 3.45996
R2977 ena.n1 ena 1.55726
R2978 ena.n2 ena 0.746125
R2979 vg1.n10 vg1.t0 85.228
R2980 vg1.n0 vg1.t3 61.1305
R2981 vg1.n7 vg1.t5 54.828
R2982 vg1.n7 vg1.t0 54.828
R2983 vg1.n5 vg1.t2 42.6599
R2984 vg1.n8 vg1.n7 32.9015
R2985 vg1.n10 vg1.n9 30.9745
R2986 vg1.n9 vg1.t1 20.9512
R2987 vg1.n6 vg1.n5 3.63479
R2988 vg1.n11 vg1.n10 2.3255
R2989 vg1.n12 vg1.n0 0.471594
R2990 vg1.n5 vg1.n4 0.390524
R2991 vg1.n9 vg1.n8 0.238607
R2992 vg1.n11 vg1.n6 0.176742
R2993 vg1 vg1.n12 0.133236
R2994 vg1.n1 vg1.t9 0.0767969
R2995 vg1.n2 vg1.n1 0.0752537
R2996 vg1.n3 vg1.n2 0.0752537
R2997 vg1.n4 vg1.t8 0.0717511
R2998 vg1.n0 vg1 0.0387813
R2999 vg1.n12 vg1.n11 0.0257152
R3000 vg1.n8 vg1.n6 0.0123355
R3001 vg1.n4 vg1.n3 0.00554581
R3002 vg1.n1 vg1.t4 0.00204321
R3003 vg1.n2 vg1.t7 0.00204321
R3004 vg1.n3 vg1.t6 0.00204321
R3005 xin.n36 xin.t8 594.832
R3006 xin.t18 xin.n5 380.808
R3007 xin.n6 xin.t18 380.808
R3008 xin.n6 xin.t15 380.611
R3009 xin.t15 xin.n5 380.611
R3010 xin.t13 xin.n7 380.611
R3011 xin.n8 xin.t13 380.611
R3012 xin.t19 xin.n4 380.611
R3013 xin.n9 xin.t19 380.611
R3014 xin.n11 xin.t16 380.611
R3015 xin.t16 xin.n10 380.611
R3016 xin.n12 xin.t11 380.611
R3017 xin.t11 xin.n3 380.611
R3018 xin.t10 xin.n13 380.611
R3019 xin.n14 xin.t10 380.611
R3020 xin.t17 xin.n2 380.611
R3021 xin.n15 xin.t17 380.611
R3022 xin.n17 xin.t14 380.611
R3023 xin.t14 xin.n16 380.611
R3024 xin.n18 xin.t12 380.611
R3025 xin.t12 xin.n1 380.611
R3026 xin.t9 xin.n19 380.611
R3027 xin.n20 xin.t9 380.611
R3028 xin.n21 xin.t6 380.611
R3029 xin.t6 xin.n0 380.611
R3030 xin.n36 xin.t21 194.639
R3031 xin.n25 xin.t20 124.457
R3032 xin.n25 xin.t7 106.793
R3033 xin.t7 xin.n23 86.3125
R3034 xin.t20 xin.n24 86.3125
R3035 xin.n24 xin.n23 58.6245
R3036 xin.n30 xin.t5 45.927
R3037 xin.n28 xin.n27 20.1298
R3038 xin.n27 xin.n23 12.2455
R3039 xin.n35 xin.n34 4.04311
R3040 xin.n26 xin.n24 3.56553
R3041 xin.n34 xin.n29 3.51336
R3042 xin.n30 xin.n29 3.51061
R3043 xin.n28 xin.n22 1.95915
R3044 xin.n35 xin.n28 1.1106
R3045 xin.n22 xin.n21 0.8105
R3046 xin.n22 xin.n0 0.7905
R3047 xin.n27 xin.n26 0.741791
R3048 xin.n26 xin.n25 0.715885
R3049 xin.n36 xin.n35 0.4755
R3050 xin xin.n36 0.377063
R3051 xin.n8 xin.n5 0.198
R3052 xin.n9 xin.n8 0.198
R3053 xin.n10 xin.n9 0.198
R3054 xin.n10 xin.n3 0.198
R3055 xin.n14 xin.n3 0.198
R3056 xin.n15 xin.n14 0.198
R3057 xin.n16 xin.n15 0.198
R3058 xin.n16 xin.n1 0.198
R3059 xin.n20 xin.n1 0.198
R3060 xin.n21 xin.n20 0.198
R3061 xin.n7 xin.n6 0.198
R3062 xin.n7 xin.n4 0.198
R3063 xin.n11 xin.n4 0.198
R3064 xin.n12 xin.n11 0.198
R3065 xin.n13 xin.n12 0.198
R3066 xin.n13 xin.n2 0.198
R3067 xin.n17 xin.n2 0.198
R3068 xin.n18 xin.n17 0.198
R3069 xin.n19 xin.n18 0.198
R3070 xin.n19 xin.n0 0.198
R3071 xin.t3 xin.t1 0.0760058
R3072 xin.n31 xin.n30 0.0410952
R3073 xin.n32 xin.n29 0.0410952
R3074 xin.n34 xin.n33 0.0410952
R3075 xin.n32 xin.t4 0.0264927
R3076 xin.n31 xin.t0 0.0264885
R3077 xin.n33 xin.t3 0.0264703
R3078 xin.n33 xin.t2 0.0264296
R3079 xin.t2 xin.n32 0.0264114
R3080 xin.t4 xin.n31 0.0264072
R3081 vg2.n2 vg2.t9 87.8852
R3082 vg2.n9 vg2.t5 87.8852
R3083 vg2.n5 vg2.t6 85.228
R3084 vg2.n12 vg2.t7 85.228
R3085 vg2.n15 vg2.t8 67.0783
R3086 vg2.n4 vg2.t9 54.828
R3087 vg2.t6 vg2.n4 54.828
R3088 vg2.n11 vg2.t5 54.828
R3089 vg2.t7 vg2.n11 54.828
R3090 vg2.n16 vg2.t0 42.6015
R3091 vg2.n4 vg2.n3 30.4005
R3092 vg2.n11 vg2.n10 30.4005
R3093 vg2.n3 vg2.n1 29.1205
R3094 vg2.n5 vg2.n1 29.1205
R3095 vg2.n10 vg2.n8 29.1205
R3096 vg2.n12 vg2.n8 29.1205
R3097 vg2.n6 vg2.n5 2.3255
R3098 vg2.n13 vg2.n12 2.3255
R3099 vg2.n3 vg2.n2 2.13477
R3100 vg2.n10 vg2.n9 2.13477
R3101 vg2 vg2.n14 0.742464
R3102 vg2.n16 vg2.n15 0.714193
R3103 vg2.n14 vg2.n6 0.474719
R3104 vg2.n14 vg2.n13 0.474719
R3105 vg2.n1 vg2.n0 0.423227
R3106 vg2.n8 vg2.n7 0.423227
R3107 vg2.n2 vg2.n0 0.308459
R3108 vg2.n9 vg2.n7 0.308459
R3109 vg2.n6 vg2.n0 0.284875
R3110 vg2.n13 vg2.n7 0.284875
R3111 vg2.n15 vg2.t3 0.170134
R3112 vg2 vg2.n16 0.119455
R3113 vg2.t1 vg2.t2 0.0652716
R3114 vg2.t4 vg2.t1 0.0652716
R3115 vg2.t3 vg2.t4 0.0652716
R3116 vrb.n2 vrb.t0 43.1048
R3117 vrb.n0 vrb.t4 22.3777
R3118 vrb.n1 vrb.t1 22.1989
R3119 vrb.n1 vrb.t3 21.3671
R3120 vrb.n0 vrb.t2 21.3663
R3121 vrb.n3 vrb.n2 1.11856
R3122 vrb.n3 vrb.n0 0.759192
R3123 vrb.n2 vrb.n1 0.758408
R3124 vrb vrb.n3 0.0491111
R3125 vn.t9 vn.n4 182.935
R3126 vn.t5 vn.n1 144.126
R3127 vn.n9 vn.n6 97.2442
R3128 vn.n10 vn.n4 97.2442
R3129 vn.n5 vn.t9 88.2031
R3130 vn.t8 vn.n4 85.228
R3131 vn.n6 vn.t8 85.228
R3132 vn.n10 vn.t3 85.228
R3133 vn.t3 vn.n9 85.228
R3134 vn.n2 vn.t5 85.228
R3135 vn.n0 vn.t2 64.2147
R3136 vn.n8 vn.n2 58.8987
R3137 vn.n0 vn.n3 56.3112
R3138 vn vn.t7 21.1687
R3139 vn.n9 vn.n8 17.975
R3140 vn.n10 vn.n1 17.975
R3141 vn vn.n7 16.8187
R3142 vn.n3 vn.t0 6.92425
R3143 vn.n3 vn.t1 6.92425
R3144 vn.n7 vn.t4 4.3505
R3145 vn.n7 vn.t6 4.3505
R3146 vn vn.n2 2.80102
R3147 vn.n9 vn 2.44682
R3148 vn.n4 vn 2.3255
R3149 vn vn.n10 2.3255
R3150 vn.n6 vn.n5 2.20282
R3151 vn.n5 vn 1.25668
R3152 vn.n8 vn 2.69718
R3153 vn vn.n1 2.67028
R3154 vn vn.n0 2.03836
R3155 x3.out.n3 x3.out.t6 393.144
R3156 x3.out.n5 x3.out.t7 393.144
R3157 x3.out.n4 x3.out.t6 391.815
R3158 x3.out.t7 x3.out.n2 391.815
R3159 x3.out.n5 x3.out.t4 371.31
R3160 x3.out.t4 x3.out.n2 371.31
R3161 x3.out.t3 x3.out.n1 371.31
R3162 x3.out.n6 x3.out.t3 371.31
R3163 x3.out.n4 x3.out.t8 371.31
R3164 x3.out.t8 x3.out.n3 371.31
R3165 x3.out.n0 x3.out.t0 227.886
R3166 x3.out.n0 x3.out.n9 25.0903
R3167 x3.out.n1 x3.out.n5 21.8335
R3168 x3.out.n3 x3.out.n1 21.6959
R3169 x3.out.n6 x3.out.n4 20.5053
R3170 x3.out.n7 x3.out.n2 19.6003
R3171 x3.out.n0 x3.out.t5 12.7763
R3172 x3.out.n9 x3.out.t1 5.5105
R3173 x3.out.n9 x3.out.t2 5.5105
R3174 x3.out.n8 x3.out.n1 5.0449
R3175 x3.out.n8 x3.out.n7 2.71826
R3176 x3.out.n7 x3.out.n6 0.90555
R3177 x3.out x3.out.n8 0.88175
R3178 x3.out x3.out.n0 0.794875
R3179 x4.out_b.n0 x4.out_b.t2 227.887
R3180 x4.out_b.n0 x4.out_b.n1 25.0905
R3181 x4.out_b.n0 x4.out_b.t3 12.777
R3182 x4.out_b.n1 x4.out_b.t0 5.5105
R3183 x4.out_b.n1 x4.out_b.t1 5.5105
R3184 x4.out_b x4.out_b.n0 0.83175
R3185 dout.n0 dout.t0 120.561
R3186 dout.n0 dout.t1 61.4115
R3187 dout dout.n0 3.88384
R3188 a_22601_n15524.t0 a_22601_n15524.t1 120.212
R3189 a_8268_n12482.t0 a_8268_n12482.t1 193.599
C0 vn inv_in 0.137437f
C1 ibias_ip vbp 1.36181f
C2 x4.out_b avss 1.60462f
C3 inv_in dvdd 0.696511f
C4 a_2132_n14926# a_2132_n15258# 0.299356f
C5 a_15539_n2241# a_16620_n1869# 0.102355f
C6 a_21775_n2791# dvdd 0.235866f
C7 a_4857_n1521# standby_ip 0.144556f
C8 avss_ip x3.out 2.42141f
C9 dvdd_ip vbp 26.197498f
C10 a_21211_n1943# a_21036_n1869# 0.251137f
C11 a_19955_n2241# dvdd 0.844484f
C12 a_17747_n2241# a_18263_n1869# 0.104035f
C13 a_4857_n1521# dvdd 0.264852f
C14 ena_ip a_16273_n2273# 0.183844f
C15 a_14009_n2701# dvdd 0.136733f
C16 avss_ip a_2132_n17582# 0.229847f
C17 a_24530_n21010# a_24530_n21342# 0.306038f
C18 a_15705_n2791# dvdd 0.631528f
C19 x3.in_b avdd 1.00629f
C20 avss_ip a_2130_n20180# 0.234105f
C21 x7.stby_done_b a_20376_n2791# 0.179696f
C22 a_14009_n2404# x7.ena_done_b 0.173521f
C23 x7.x2.Qb2 a_19567_n2791# 0.127083f
C24 avss_ip a_2132_n15258# 0.245921f
C25 a_2130_n21176# xin 0.159603f
C26 a_17359_n2247# x7.x1.x2.Q 0.161495f
C27 a_18932_n16088# a_18932_n16420# 0.299356f
C28 ena_ip x3.in_b 0.676051f
C29 vg2 a_2132_n17582# 0.155259f
C30 a_19003_n1943# a_19567_n2247# 0.106826f
C31 xin_buf xin 1.99369f
C32 ena_ip a_18481_n2273# 0.183839f
C33 avss_ip a_24530_n21342# 0.187124f
C34 a_14009_n2404# x7.clk_disable 0.122842f
C35 dvss_ip a_10620_n9334# 0.174627f
C36 avss_ip a_18932_n16420# 0.690377f
C37 vg2 a_2132_n15258# 0.154162f
C38 xin_buf inv_in 0.113575p
C39 x7.x1.Qb1 a_17359_n2247# 0.127083f
C40 a_24530_n22338# xin 0.168028f
C41 a_20579_n2425# dvdd 0.144018f
C42 avss_ip a_24530_n19018# 0.187516f
C43 a_20689_n2273# dvdd 0.225909f
C44 a_17747_n2241# a_18828_n1869# 0.102355f
C45 avss_ip avdd 2.34938f
C46 ena_ip a_16795_n1943# 0.357273f
C47 a_24530_n20014# xin 0.159204f
C48 standby_ip ibias 0.288163f
C49 a_2130_n21176# a_2130_n21508# 0.306949f
C50 dvdd_ip vn 1.05192f
C51 a_16055_n2791# dvdd 0.234f
C52 dvdd_ip standby_ip 3.44007f
C53 a_15539_n2791# x7.x2.Qb1 0.630684f
C54 a_10620_n7674# a_10620_n8006# 0.306784f
C55 a_21211_n2817# a_21775_n2791# 0.106826f
C56 dvss_ip a_24220_n8172# 0.412162f
C57 x7.x1.x4.Q dvdd 0.118427f
C58 dvdd_ip dvdd 14.0307f
C59 xin_buf a_10620_n8006# 0.166951f
C60 a_14009_n2404# x7.stby_done_b 0.245503f
C61 dvss_ip a_18932_n16752# 0.11359f
C62 a_2132_n16254# a_2132_n16586# 0.299336f
C63 ena_ip a_19003_n1943# 0.357273f
C64 a_2130_n18852# a_2130_n19184# 0.307023f
C65 dvss_ip a_18932_n14428# 0.117297f
C66 x3.out avdd 9.26841f
C67 a_2971_n1521# ena 0.188898f
C68 inv_in xin 0.302115f
C69 xin_buf xout 3.51791f
C70 a_21211_n1943# dvdd 0.467188f
C71 x7.x1.Qb2 a_19567_n2247# 0.127083f
C72 a_24220_n8836# a_24220_n9168# 0.309571f
C73 vbp tail 10.143401f
C74 standby_33 ibias_ip 0.621612f
C75 avss_ip a_2132_n17914# 0.528436f
C76 a_16620_n2791# dvdd 0.320791f
C77 standby_33 ibias 1.10533f
C78 ibias_ip xin_buf 1.72895f
C79 x7.ena_done_b a_15000_n1881# 0.263497f
C80 avss_ip a_2130_n20512# 0.234105f
C81 dvdd_ip dout 1.66314f
C82 a_18932_n17416# a_18932_n17748# 0.299356f
C83 x7.ena_done_b a_15705_n2241# 0.195776f
C84 dvdd_ip a_10620_n7674# 0.100908f
C85 standby_ip avss 1.86774f
C86 dvdd_ip standby_33 3.26892f
C87 avss_ip a_2132_n15590# 0.241841f
C88 a_24530_n20014# a_24530_n20346# 0.307948f
C89 ena_ip x7.x1.Qb1 0.347396f
C90 dvdd_ip vrb 0.182588f
C91 a_2130_n21508# xin 0.167748f
C92 dvss_ip vbp 1.28877f
C93 dvdd_ip xin_buf 19.1703f
C94 dvdd avss 0.230567f
C95 vg2 a_2132_n17914# 0.154785f
C96 a_15539_n2791# dvdd 0.651082f
C97 a_17913_n2791# a_18481_n2549# 0.174808f
C98 avss_ip a_24530_n21674# 0.194498f
C99 a_2971_n1521# ena_ip 0.142973f
C100 a_2130_n19184# xin 0.164971f
C101 x7.x1.Qb2 a_18168_n1881# 0.171293f
C102 dvss_ip a_10620_n9666# 0.193818f
C103 a_18932_n15092# a_18932_n15424# 0.299356f
C104 vg2 a_2132_n15590# 0.156683f
C105 avss_ip a_18932_n16752# 0.452744f
C106 a_15000_n1881# x7.x1.x2.CLK 0.134958f
C107 avss_ip a_24530_n19350# 0.193645f
C108 x7.x2.Qb1 a_15960_n2791# 0.171293f
C109 x7.ena_done_b a_17913_n2241# 0.193771f
C110 a_21775_n2247# dvdd 0.236037f
C111 xin xout 12.4168f
C112 a_19003_n2817# x7.x2.x3.Q 0.119961f
C113 a_15705_n2241# a_16273_n2273# 0.174808f
C114 ena_ip x7.x1.Qb2 0.347451f
C115 avss_ip a_18932_n14428# 0.151712f
C116 a_10620_n9002# a_10620_n9334# 0.307266f
C117 a_24530_n20346# xin 0.158905f
C118 x7.stby_done_b x7.x2.Qb1 0.111333f
C119 standby_ip x7.ena_done_b 0.121215f
C120 inv_in xout 1.1656f
C121 x7.stby_done_b a_15000_n2791# 0.263439f
C122 x7.stby_done_b a_17913_n2791# 0.193805f
C123 a_2132_n17582# a_2132_n17914# 0.299336f
C124 x7.ena_done_b dvdd 6.16668f
C125 ena_ip avdd 0.711014f
C126 dvss_ip a_24220_n8504# 0.435581f
C127 xin_buf a_10620_n8338# 0.166314f
C128 inv_in inv_m1 0.243271f
C129 vg2 a_18932_n14428# 0.5683f
C130 vn tail 0.670061f
C131 a_2130_n20180# a_2130_n20512# 0.308883f
C132 standby_33 avss 1.55853f
C133 dvdd_ip xin 4.32555f
C134 a_18481_n2549# a_18263_n2791# 0.209641f
C135 x7.clk_disable dvdd 0.383458f
C136 dvss_ip a_18932_n14760# 0.144339f
C137 x7.x1.x3.Q dvdd 0.112744f
C138 a_2132_n15258# a_2132_n15590# 0.29969f
C139 a_18481_n2549# dvdd 0.225643f
C140 avdd_ip xin_buf 9.05887f
C141 dvss_ip vn 6.6789f
C142 dvdd_ip inv_in 10.408401f
C143 x7.x2.x4.Q dvdd 0.118417f
C144 vrb vg1 0.454276f
C145 x7.x1.x2.CLK dvdd 0.406962f
C146 x7.stby_done_b a_19955_n2791# 0.648907f
C147 a_19955_n2791# a_20121_n2791# 0.608363f
C148 a_16273_n2273# dvdd 0.230873f
C149 a_19567_n2791# x7.x2.x3.Q 0.161495f
C150 dvss_ip dvdd 20.2555f
C151 a_16273_n2273# a_16055_n1869# 0.209641f
C152 a_15705_n2791# a_16055_n2791# 0.219472f
C153 a_24530_n21342# a_24530_n21674# 0.307869f
C154 a_17913_n2241# a_18481_n2273# 0.174808f
C155 avss_ip a_2130_n20844# 0.234274f
C156 a_24220_n7840# a_24220_n8172# 0.307266f
C157 avss_ip a_2132_n15922# 0.231212f
C158 a_2130_n21840# xin 0.172286f
C159 x4.out_b avdd 7.47205f
C160 x7.stby_done_b dvdd 5.41509f
C161 a_20121_n2791# dvdd 0.653362f
C162 x3.in_b dvdd 0.22553f
C163 a_18932_n16420# a_18932_n16752# 0.299356f
C164 a_18481_n2273# dvdd 0.225651f
C165 a_20121_n2241# a_20471_n1869# 0.219472f
C166 avss_ip a_24530_n22006# 0.186833f
C167 ena_ip a_20471_n1869# 0.196932f
C168 ena_ip a_14009_n2404# 0.156624f
C169 a_24530_n19018# a_24530_n19350# 0.307948f
C170 a_2130_n19516# xin 0.164971f
C171 xin_buf tail 4.40803f
C172 a_19003_n2817# dvdd 0.456345f
C173 vg2 a_2132_n15922# 0.154604f
C174 avss_ip a_18932_n17084# 0.726269f
C175 avss_ip a_24530_n19682# 0.193645f
C176 avdd_ip xin 6.74409f
C177 dvdd_ip xout 4.80514f
C178 dvss_ip dout 6.66227f
C179 inv_in avss 0.144174f
C180 a_19955_n2791# a_20471_n2791# 0.104035f
C181 a_16795_n1943# dvdd 0.461387f
C182 a_20121_n2791# a_20689_n2549# 0.174808f
C183 dvss_ip a_10620_n7674# 0.359271f
C184 vg1 xin 0.215332p
C185 dvss_ip standby_33 3.27772f
C186 avss_ip a_18932_n14760# 0.178926f
C187 x7.x2.Qb2 a_17913_n2791# 0.756617f
C188 dvss_ip vrb 1.20334f
C189 ibias_ip ibias 0.846688f
C190 a_15705_n2791# a_16620_n2791# 0.125324f
C191 a_24530_n20678# xin 0.159253f
C192 dvdd_ip inv_m1 2.8465f
C193 avdd_ip inv_in 0.669037f
C194 dvss_ip xin_buf 27.955f
C195 a_2130_n21508# a_2130_n21840# 0.307948f
C196 a_18481_n2273# a_18263_n1869# 0.209641f
C197 dout_filt dvdd 1.76335f
C198 dvdd_ip ibias_ip 1.46921f
C199 a_10620_n8006# a_10620_n8338# 0.307266f
C200 x7.x1.x2.CLK a_15539_n2241# 0.240273f
C201 a_21211_n2817# x7.x2.x4.Q 0.119961f
C202 dvss_ip a_24220_n8836# 0.421193f
C203 xin_buf a_10620_n8670# 0.16582f
C204 x7.x1.Qb1 a_15705_n2241# 0.756617f
C205 a_20471_n2791# dvdd 0.234572f
C206 a_15539_n2791# a_15705_n2791# 0.608363f
C207 a_2132_n16586# a_2132_n16918# 0.298902f
C208 a_19003_n1943# dvdd 0.456365f
C209 a_20121_n2241# a_21036_n1869# 0.125324f
C210 a_19003_n2817# a_18828_n2791# 0.251137f
C211 ena_ip a_21036_n1869# 0.254262f
C212 a_2130_n19184# a_2130_n19516# 0.308883f
C213 x7.x2.Qb2 a_19955_n2791# 0.241144f
C214 dvss_ip a_18932_n15092# 0.147461f
C215 a_19567_n2791# dvdd 0.230807f
C216 tail xin 1.6128f
C217 x7.ena_done_b a_19955_n2241# 0.648846f
C218 a_20689_n2549# a_20471_n2791# 0.209641f
C219 a_19955_n2791# a_21036_n2791# 0.102355f
C220 a_17359_n2247# dvdd 0.234839f
C221 a_2132_n14262# a_2132_n14594# 0.299692f
C222 a_16795_n1943# a_16620_n1869# 0.251137f
C223 inv_m1 inv_m2 0.947856f
C224 inv_in tail 0.604094f
C225 a_21211_n1943# x7.x1.x4.Q 0.119961f
C226 x7.x1.x2.Q dvdd 0.116301f
C227 a_24220_n9168# a_24220_n9500# 0.30635f
C228 dout_filt dout 0.639323f
C229 x7.x2.Qb2 dvdd 1.2179f
C230 avdd_ip xout 7.21813f
C231 dvss_ip xin 1.63056f
C232 avss_ip a_2130_n21176# 0.242612f
C233 a_18932_n17748# vg1 0.408298f
C234 vg1 xout 0.637062f
C235 avss_ip vrb 6.48162f
C236 a_21775_n2791# x7.x2.x4.Q 0.161495f
C237 dvss_ip inv_in 14.9291f
C238 avss_ip xin_buf 10.8147f
C239 x7.x1.Qb1 dvdd 1.22948f
C240 dvdd_ip inv_m2 1.90217f
C241 avss_ip a_2132_n16254# 0.230757f
C242 a_24530_n20346# a_24530_n20678# 0.307948f
C243 a_2130_n22172# xin 0.581116f
C244 a_21036_n2791# dvdd 0.31454f
C245 a_15539_n2791# a_16055_n2791# 0.104035f
C246 x7.clk_disable a_14009_n2701# 0.419961f
C247 a_15000_n2791# x7.x2.x2.CLK 0.134958f
C248 avss_ip a_2130_n18852# 0.557241f
C249 a_18932_n15424# vg1 0.560332f
C250 a_19567_n2247# dvdd 0.230816f
C251 x7.x1.Qb2 a_17913_n2241# 0.756617f
C252 a_2971_n1521# dvdd 0.261493f
C253 avss_ip a_24530_n22338# 0.488441f
C254 a_2130_n19848# xin 0.165429f
C255 vg2 vrb 4.64006f
C256 a_18932_n15424# a_18932_n15756# 0.299356f
C257 a_18371_n2425# dvdd 0.143768f
C258 xin_buf vg2 3.5685f
C259 vg2 a_2132_n16254# 0.155116f
C260 dvdd_ip avdd_ip 3.59467f
C261 avss_ip a_18932_n17416# 0.56453f
C262 dvdd ena 0.377442f
C263 avss_ip a_24530_n20014# 0.193645f
C264 dvdd_ip vg1 0.707385f
C265 x7.stby_done_b a_21775_n2791# 0.160191f
C266 x7.x1.Qb2 dvdd 1.22125f
C267 dvss_ip a_10620_n8006# 0.203148f
C268 avss_ip a_18932_n15092# 0.193668f
C269 a_21775_n2247# x7.x1.x4.Q 0.161495f
C270 a_16795_n2817# a_17359_n2791# 0.106826f
C271 a_10620_n9334# a_10620_n9666# 0.310516f
C272 a_24530_n21010# xin 0.159641f
C273 standby_ip avdd 0.690112f
C274 tail xout 1.23159f
C275 a_19003_n1943# a_18828_n1869# 0.251137f
C276 avdd dvdd 0.106948f
C277 x7.stby_done_b a_15705_n2791# 0.20129f
C278 dvss_ip a_24220_n9168# 0.4382f
C279 xin_buf a_10620_n9002# 0.156922f
C280 a_17747_n2791# x7.x2.Qb2 0.630684f
C281 a_2130_n20512# a_2130_n20844# 0.307948f
C282 a_15539_n2791# a_16620_n2791# 0.102355f
C283 ena_ip standby_ip 4.63202f
C284 dvss_ip xout 14.2041f
C285 avss_ip xin 73.1079f
C286 a_20121_n2241# dvdd 0.655086f
C287 a_21211_n1943# a_21775_n2247# 0.106826f
C288 ena_ip dvdd 7.78413f
C289 ena_ip a_16055_n1869# 0.196968f
C290 dvdd_ip tail 3.21426f
C291 dvss_ip inv_m1 3.10099f
C292 avss_ip inv_in 1.9489f
C293 x7.x2.x2.CLK dvdd 0.367738f
C294 a_2132_n15590# a_2132_n15922# 0.298886f
C295 a_16273_n2549# dvdd 0.232251f
C296 dvss_ip ibias_ip 20.300303f
C297 a_15539_n2241# x7.x1.Qb1 0.630684f
C298 vg2 xin 6.28706f
C299 avdd_ip avss 0.574893f
C300 a_21211_n2817# a_21036_n2791# 0.251137f
C301 a_14009_n2701# dout_filt 0.140187f
C302 x7.x2.Qb2 a_18168_n2791# 0.171293f
C303 a_20579_n2247# dvdd 0.144024f
C304 inv_in vg2 0.137694f
C305 dvdd_ip dvss_ip 0.502455p
C306 a_24530_n21674# a_24530_n22006# 0.306949f
C307 avdd_ip vg1 1.99589f
C308 ena_ip a_18263_n1869# 0.196932f
C309 avss_ip a_2130_n21508# 0.234275f
C310 standby_33 avdd 9.00234f
C311 a_24220_n8172# a_24220_n8504# 0.310516f
C312 xin_buf avdd 0.176178f
C313 avss_ip a_2132_n16586# 0.229609f
C314 x7.x1.Qb1 a_17747_n2241# 0.241144f
C315 x7.x2.Qb1 a_17359_n2791# 0.127083f
C316 avss_ip a_2130_n19184# 0.234105f
C317 a_18932_n15756# vg1 0.267005f
C318 a_18932_n16752# a_18932_n17084# 0.299356f
C319 a_20471_n1869# dvdd 0.234574f
C320 standby_ip x4.out_b 0.931668f
C321 a_14009_n2404# a_14285_n2281# 0.143754f
C322 a_14009_n2404# dvdd 0.221473f
C323 ena_ip a_16620_n1869# 0.25803f
C324 avss_ip a_2132_n14262# 1.08299f
C325 a_24530_n19350# a_24530_n19682# 0.307948f
C326 a_2130_n20180# xin 0.1652f
C327 a_16795_n2817# x7.x2.x2.Q 0.119961f
C328 avss_ip a_18932_n17748# 0.633601f
C329 vg2 a_2132_n16586# 0.154861f
C330 avss_ip xout 26.396301f
C331 a_16795_n2817# dvdd 0.462729f
C332 avss_ip a_24530_n20346# 0.193441f
C333 x7.ena_done_b a_21775_n2247# 0.160065f
C334 dvss_ip a_10620_n8338# 0.203056f
C335 dvss_ip inv_m2 1.69963f
C336 a_18932_n14428# a_18932_n14760# 0.299356f
C337 a_17747_n2241# x7.x1.Qb2 0.630684f
C338 avss_ip a_18932_n15424# 0.222697f
C339 ena_ip a_15539_n2241# 0.611445f
C340 a_24530_n21342# xin 0.166712f
C341 vg2 xout 0.938912f
C342 a_2130_n21840# a_2130_n22172# 0.306949f
C343 ena_ip a_18828_n1869# 0.25803f
C344 dvdd_ip dout_filt 2.6369f
C345 a_10620_n8338# a_10620_n8670# 0.307266f
C346 a_24530_n19018# xin 0.126575f
C347 inv_in a_24220_n7840# 0.423473f
C348 dvss_ip a_24220_n9500# 0.412902f
C349 dvdd_ip avss_ip 2.2865f
C350 avdd_ip dvss_ip 20.735699f
C351 xin_buf a_10620_n9334# 0.138691f
C352 dvss_ip vg1 6.37401f
C353 a_2132_n16918# a_2132_n17250# 0.299677f
C354 a_21036_n1869# dvdd 0.31455f
C355 x7.x1.Qb2 a_19955_n2241# 0.241144f
C356 dvdd standby 0.386478f
C357 ena_ip a_17747_n2241# 0.61356f
C358 a_2130_n19516# a_2130_n19848# 0.307948f
C359 x3.in_b avss 1.85499f
C360 dvss_ip a_18932_n15756# 0.124217f
C361 a_17359_n2791# x7.x2.x2.Q 0.161495f
C362 standby_33 x4.out_b 0.696369f
C363 dvdd_ip vg2 0.10449f
C364 x7.x2.x3.Q dvdd 0.112734f
C365 a_17359_n2791# dvdd 0.236098f
C366 dvss_ip x7.ena_done_b 1.48709f
C367 a_2132_n14594# a_2132_n14926# 0.298902f
C368 a_24220_n9500# a_24220_n9832# 0.307266f
C369 a_19955_n2241# a_20121_n2241# 0.608363f
C370 a_17913_n2791# a_18263_n2791# 0.219472f
C371 x7.x2.Qb1 dvdd 1.15446f
C372 avss_ip a_2130_n21840# 0.234358f
C373 ena_ip a_19955_n2241# 0.613409f
C374 dvss_ip tail 0.416372f
C375 a_15000_n2791# dvdd 0.238886f
C376 a_18371_n2247# dvdd 0.143775f
C377 a_17913_n2791# dvdd 0.653627f
C378 x7.ena_done_b x7.stby_done_b 1.61077f
C379 avss_ip a_2132_n16918# 0.236584f
C380 a_24530_n20678# a_24530_n21010# 0.307948f
C381 avss_ip a_2130_n19516# 0.234105f
C382 a_15000_n1881# dvdd 0.25026f
C383 avss_ip avss 7.31391f
C384 a_14285_n2079# dvdd 0.149051f
C385 a_15705_n2241# dvdd 0.668389f
C386 a_24530_n19018# xout 0.377144f
C387 a_15705_n2241# a_16055_n1869# 0.219472f
C388 avss_ip a_2132_n14594# 0.792432f
C389 a_2130_n20512# xin 0.164971f
C390 a_15705_n2791# a_16273_n2549# 0.174808f
C391 avdd_ip avss_ip 0.856941p
C392 a_18932_n15756# a_18932_n16088# 0.299356f
C393 vg2 a_2132_n16918# 0.156129f
C394 avss_ip vg1 20.7774f
C395 x7.stby_done_b x7.clk_disable 0.724301f
C396 avss_ip a_24530_n20678# 0.193645f
C397 dvss_ip a_10620_n8670# 0.203056f
C398 x7.ena_done_b a_20376_n1881# 0.179696f
C399 avss_ip a_18932_n15756# 0.237057f
C400 a_24530_n21674# xin 0.159429f
C401 avdd_ip vg2 0.488655f
C402 a_19955_n2791# dvdd 0.843855f
C403 dvss_ip x7.stby_done_b 1.50194f
C404 vbp xin_buf 3.4756f
C405 vg2 vg1 1.36272f
C406 a_19955_n2241# a_20471_n1869# 0.104035f
C407 a_17913_n2241# dvdd 0.655351f
C408 a_20121_n2241# a_20689_n2273# 0.174808f
C409 a_17913_n2791# a_18828_n2791# 0.125324f
C410 ena_ip a_20689_n2273# 0.183839f
C411 a_24530_n19350# xin 0.159253f
C412 x3.out avss 5.85073f
C413 dvss_ip a_24220_n9832# 0.676369f
C414 a_18263_n2791# dvdd 0.23444f
C415 xin_buf a_10620_n9666# 0.140848f
C416 standby_ip dvdd 10.280701f
C417 a_2130_n20844# a_2130_n21176# 0.306949f
C418 x7.x2.Qb1 a_17747_n2791# 0.241144f
C419 x7.x1.Qb1 a_15960_n1881# 0.171293f
C420 x7.x2.x2.Q dvdd 0.11753f
C421 ena_ip ibias 0.171255f
C422 x7.stby_done_b a_20121_n2791# 0.953635f
C423 x7.clk_disable dout_filt 0.71038f
C424 a_14285_n2281# dvdd 0.170927f
C425 a_16055_n1869# dvdd 0.237126f
C426 a_15705_n2241# a_16620_n1869# 0.125324f
C427 a_17747_n2791# a_17913_n2791# 0.608363f
C428 a_16273_n2549# a_16055_n2791# 0.209641f
C429 a_2132_n15922# a_2132_n16254# 0.300147f
C430 a_17913_n2241# a_18263_n1869# 0.219472f
C431 a_16163_n2425# dvdd 0.147354f
C432 dvss_ip dout_filt 7.440259f
C433 a_19003_n1943# x7.x1.x3.Q 0.119961f
C434 avss_ip a_3134_n13324# 1.13338f
C435 dvss_ip avss_ip 23.869501f
C436 a_15539_n2241# a_15705_n2241# 0.608363f
C437 a_20689_n2549# dvdd 0.225901f
C438 a_18263_n1869# dvdd 0.234443f
C439 a_19955_n2241# a_21036_n1869# 0.102355f
C440 a_20689_n2273# a_20471_n1869# 0.209641f
C441 a_24530_n22006# a_24530_n22338# 0.307023f
C442 avss_ip a_2130_n22172# 0.237164f
C443 ena_ip a_21211_n1943# 0.305293f
C444 a_24220_n8504# a_24220_n8836# 0.309571f
C445 a_4857_n1521# standby 0.18913f
C446 x7.stby_done_b dout_filt 0.19319f
C447 dvss_ip vg2 3.9276f
C448 avss_ip a_2132_n17250# 0.236693f
C449 a_18828_n2791# dvdd 0.312702f
C450 vbp inv_in 0.265485f
C451 dvdd dout 0.550876f
C452 vn xin_buf 4.74796f
C453 avdd avss 0.110507p
C454 avss_ip a_2130_n19848# 0.234105f
C455 a_18932_n17084# a_18932_n17416# 0.299356f
C456 a_20121_n2791# a_20471_n2791# 0.219472f
C457 a_16620_n1869# dvdd 0.318883f
C458 a_17747_n2791# a_18263_n2791# 0.104035f
C459 avdd_ip avdd 9.33419f
C460 avss_ip a_2132_n14926# 0.652798f
C461 a_16163_n2247# dvdd 0.146808f
C462 a_24530_n19682# a_24530_n20014# 0.307948f
C463 a_2130_n20844# xin 0.166057f
C464 vg2 a_2132_n17250# 0.155881f
C465 ena_ip avss 1.87755f
C466 a_17747_n2791# dvdd 0.843691f
C467 a_17913_n2241# a_18828_n1869# 0.125324f
C468 avss_ip a_24530_n21010# 0.193969f
C469 a_19567_n2247# x7.x1.x3.Q 0.161495f
C470 x7.x2.x2.CLK a_15539_n2791# 0.240273f
C471 dvss_ip a_10620_n9002# 0.19184f
C472 a_18932_n14760# a_18932_n15092# 0.299356f
C473 a_15539_n2241# dvdd 0.844577f
C474 avss_ip a_18932_n16088# 0.544237f
C475 a_15539_n2241# a_16055_n1869# 0.104035f
C476 a_24530_n22006# xin 0.166657f
C477 a_21211_n2817# dvdd 0.467216f
C478 x7.x2.Qb1 a_15705_n2791# 0.756617f
C479 a_18828_n1869# dvdd 0.312712f
C480 a_17747_n2241# a_17913_n2241# 0.608363f
C481 a_19003_n2817# a_19567_n2791# 0.106826f
C482 a_24530_n19682# xin 0.159253f
C483 a_10620_n8670# a_10620_n9002# 0.307266f
C484 x3.in_b x3.out 0.933643f
C485 vn xin 3.09633f
C486 a_2132_n17250# a_2132_n17582# 0.299692f
C487 x7.ena_done_b a_20121_n2241# 0.953602f
C488 ena_ip x7.ena_done_b 0.702741f
C489 a_20121_n2791# a_21036_n2791# 0.125324f
C490 a_17747_n2241# dvdd 0.844319f
C491 dvss_ip a_24220_n7840# 0.402598f
C492 a_16795_n1943# a_17359_n2247# 0.106826f
C493 a_17747_n2791# a_18828_n2791# 0.102355f
C494 xin_buf a_10620_n7674# 0.173169f
C495 standby_33 xin_buf 2.34818f
C496 a_2130_n19848# a_2130_n20180# 0.307023f
C497 a_16795_n2817# a_16620_n2791# 0.251137f
C498 avss_ip vg2 0.156017p
C499 a_16795_n1943# x7.x1.x2.Q 0.119961f
C500 xout dvss 4.260475f
C501 xin dvss 11.878201f
C502 dout dvss 6.13496f
C503 standby dvss 1.31628f
C504 ena dvss 1.29685f
C505 avss dvss 11.55251f
C506 ibias dvss 6.38685f
C507 dvdd dvss 0.140297p
C508 avdd dvss 95.102425f
C509 a_24530_n22338# dvss 0.197063f
C510 a_2130_n22172# dvss 0.199586f
C511 a_24530_n22006# dvss 0.197123f
C512 a_2130_n21840# dvss 0.205689f
C513 a_24530_n21674# dvss 0.191047f
C514 a_2130_n21508# dvss 0.205669f
C515 a_24530_n21342# dvss 0.197488f
C516 a_2130_n21176# dvss 0.199691f
C517 a_24530_n21010# dvss 0.191047f
C518 a_2130_n20844# dvss 0.20567f
C519 a_24530_n20678# dvss 0.191047f
C520 a_2130_n20512# dvss 0.205512f
C521 a_24530_n20346# dvss 0.190888f
C522 a_2130_n20180# dvss 0.205515f
C523 a_24530_n20014# dvss 0.190952f
C524 a_2130_n19848# dvss 0.205518f
C525 a_24530_n19682# dvss 0.191047f
C526 a_2130_n19516# dvss 0.205512f
C527 a_24530_n19350# dvss 0.191047f
C528 a_2130_n19184# dvss 0.205515f
C529 a_24530_n19018# dvss 0.191047f
C530 a_2130_n18852# dvss 0.205518f
C531 vg1 dvss -0.243245f
C532 a_2132_n17914# dvss 0.204459f
C533 a_18932_n17748# dvss 0.183093f
C534 a_2132_n17582# dvss 0.204591f
C535 a_18932_n17416# dvss 0.183093f
C536 a_2132_n17250# dvss 0.199339f
C537 a_18932_n17084# dvss 0.183093f
C538 a_2132_n16918# dvss 0.199339f
C539 a_18932_n16752# dvss 0.183093f
C540 a_2132_n16586# dvss 0.204459f
C541 a_18932_n16420# dvss 0.183093f
C542 a_2132_n16254# dvss 0.204591f
C543 a_18932_n16088# dvss 0.183093f
C544 a_2132_n15922# dvss 0.204459f
C545 a_18932_n15756# dvss 0.182956f
C546 a_2132_n15590# dvss 0.199472f
C547 a_18932_n15424# dvss 0.182179f
C548 a_2132_n15258# dvss 0.204459f
C549 a_18932_n15092# dvss 0.207654f
C550 a_2132_n14926# dvss 0.204459f
C551 a_18932_n14760# dvss 0.204459f
C552 a_2132_n14594# dvss 0.205118f
C553 a_18932_n14428# dvss 0.179624f
C554 a_2132_n14262# dvss 0.204591f
C555 vrb dvss 0.16284f
C556 a_3134_n13324# dvss 0.190586f
C557 vg2 dvss 4.397135f
C558 a_24220_n9832# dvss 0.206087f
C559 a_10620_n9666# dvss 0.186956f
C560 a_24220_n9500# dvss 0.206087f
C561 a_10620_n9334# dvss 0.205627f
C562 a_24220_n9168# dvss 0.187048f
C563 a_10620_n9002# dvss 0.205994f
C564 a_24220_n8836# dvss 0.186681f
C565 a_10620_n8670# dvss 0.205994f
C566 a_24220_n8504# dvss 0.186681f
C567 a_10620_n8338# dvss 0.205994f
C568 a_24220_n8172# dvss 0.20572f
C569 a_10620_n8006# dvss 0.205994f
C570 a_24220_n7840# dvss 0.206087f
C571 a_10620_n7674# dvss 0.200388f
C572 tail dvss 12.477897f
C573 inv_m2 dvss 0.562228f
C574 inv_m1 dvss 0.704134f
C575 inv_in dvss 6.596221f
C576 xin_buf dvss 7.43464f
C577 vn dvss 4.91315f
C578 vbp dvss 19.58865f
C579 x4.out_b dvss 1.061455f
C580 x3.out dvss 2.07027f
C581 a_21775_n2791# dvss 0.2255f
C582 a_21036_n2791# dvss 0.266719f
C583 a_21211_n2817# dvss 0.721269f
C584 a_20471_n2791# dvss 0.269124f
C585 a_20689_n2549# dvss 0.185767f
C586 a_20121_n2791# dvss 0.307225f
C587 a_19955_n2791# dvss 0.565683f
C588 a_19567_n2791# dvss 0.198301f
C589 a_18828_n2791# dvss 0.263274f
C590 a_19003_n2817# dvss 0.699257f
C591 a_18263_n2791# dvss 0.269103f
C592 a_18481_n2549# dvss 0.18572f
C593 a_17913_n2791# dvss 0.307195f
C594 x7.x2.Qb2 dvss 0.510929f
C595 a_17747_n2791# dvss 0.56557f
C596 dout_filt dvss 5.8975f
C597 a_17359_n2791# dvss 0.198798f
C598 a_16620_n2791# dvss 0.264546f
C599 a_16795_n2817# dvss 0.700156f
C600 a_16055_n2791# dvss 0.276301f
C601 a_16273_n2549# dvss 0.187951f
C602 a_15705_n2791# dvss 0.351701f
C603 x7.x2.Qb1 dvss 0.540099f
C604 a_15539_n2791# dvss 0.620802f
C605 x7.x2.x2.CLK dvss 0.389657f
C606 a_14009_n2701# dvss 0.233987f
C607 x7.clk_disable dvss 4.60726f
C608 a_15000_n2791# dvss 0.342356f
C609 x7.stby_done_b dvss 2.67735f
C610 ibias_ip dvss 13.1769f
C611 standby_33 dvss 13.62504f
C612 a_21775_n2247# dvss 0.225515f
C613 a_21036_n1869# dvss 0.266723f
C614 a_21211_n1943# dvss 0.721243f
C615 a_20471_n1869# dvss 0.269077f
C616 a_20689_n2273# dvss 0.185771f
C617 a_20121_n2241# dvss 0.307238f
C618 a_19955_n2241# dvss 0.56568f
C619 a_19567_n2247# dvss 0.198316f
C620 a_18828_n1869# dvss 0.263277f
C621 a_19003_n1943# dvss 0.699232f
C622 a_18263_n1869# dvss 0.269056f
C623 a_18481_n2273# dvss 0.185724f
C624 a_17913_n2241# dvss 0.307208f
C625 x7.x1.Qb2 dvss 0.510897f
C626 a_17747_n2241# dvss 0.565567f
C627 a_17359_n2247# dvss 0.198813f
C628 a_16620_n1869# dvss 0.264549f
C629 a_16795_n1943# dvss 0.70013f
C630 a_16055_n1869# dvss 0.271684f
C631 a_16273_n2273# dvss 0.187955f
C632 a_15705_n2241# dvss 0.341334f
C633 x7.x1.Qb1 dvss 0.528095f
C634 a_15539_n2241# dvss 0.580494f
C635 x7.x1.x2.CLK dvss 0.38222f
C636 a_15000_n1881# dvss 0.351108f
C637 x7.ena_done_b dvss 5.912164f
C638 a_14009_n2404# dvss 0.605583f
C639 x3.in_b dvss 1.85375f
C640 standby_ip dvss 20.4485f
C641 ena_ip dvss 14.4202f
C642 a_4857_n1521# dvss 0.293752f
C643 a_2971_n1521# dvss 0.292633f
C644 avss_ip dvss 29.749199f
C645 dvss_ip dvss 41.9846f
C646 avdd_ip dvss 0.98484p
C647 dvdd_ip dvss 0.352295p
C648 a_8268_n12482.t1 dvss 3.56607f
C649 a_22601_n15524.t1 dvss 1.2f
C650 a_22601_n15524.t0 dvss 1.2f
C651 dout.t1 dvss 0.223213f
C652 dout.n0 dvss 3.29562f
C653 x4.out_b.n0 dvss 5.53652f
C654 x4.out_b.t3 dvss 1.30743f
C655 x4.out_b.n1 dvss 0.140668f
C656 x3.out.n0 dvss 7.39524f
C657 x3.out.n1 dvss 0.893601f
C658 x3.out.n2 dvss 0.392503f
C659 x3.out.t6 dvss 0.479128f
C660 x3.out.n3 dvss 0.382459f
C661 x3.out.t8 dvss 0.458669f
C662 x3.out.n4 dvss 0.394877f
C663 x3.out.t7 dvss 0.479113f
C664 x3.out.t4 dvss 0.458669f
C665 x3.out.n5 dvss 0.382543f
C666 x3.out.t3 dvss 0.458669f
C667 x3.out.n6 dvss 0.161457f
C668 x3.out.n7 dvss 0.521199f
C669 x3.out.n8 dvss 1.69978f
C670 x3.out.t5 dvss 1.7568f
C671 x3.out.n9 dvss 0.188953f
C672 vn.n0 dvss 2.86008f
C673 vn.n1 dvss 0.636215f
C674 vn.n2 dvss 0.311146f
C675 vn.n3 dvss 0.106375f
C676 vn.t2 dvss 0.171883f
C677 vn.n4 dvss 0.444704f
C678 vn.t8 dvss 0.871134f
C679 vn.t9 dvss 1.02426f
C680 vn.n5 dvss 0.591267f
C681 vn.n6 dvss 0.320978f
C682 vn.t5 dvss 0.973785f
C683 vn.t7 dvss 0.133384f
C684 vn.n8 dvss 0.489753f
C685 vn.n9 dvss 0.299827f
C686 vn.t3 dvss 0.871134f
C687 vn.n10 dvss 0.296493f
C688 vrb.t2 dvss 0.274519f
C689 vrb.t4 dvss 0.33602f
C690 vrb.n0 dvss 3.02505f
C691 vrb.t3 dvss 0.274548f
C692 vrb.t1 dvss 0.333171f
C693 vrb.n1 dvss 3.02989f
C694 vrb.n2 dvss 2.40037f
C695 vrb.n3 dvss 1.30448f
C696 vg2.n0 dvss 0.282949f
C697 vg2.n1 dvss 0.261019f
C698 vg2.t9 dvss 0.640509f
C699 vg2.n2 dvss 1.17147f
C700 vg2.n3 dvss 0.244906f
C701 vg2.n4 dvss 0.522037f
C702 vg2.t6 dvss 0.628646f
C703 vg2.n5 dvss 0.314177f
C704 vg2.n6 dvss 0.32051f
C705 vg2.n7 dvss 0.282949f
C706 vg2.n8 dvss 0.261019f
C707 vg2.t5 dvss 0.640544f
C708 vg2.n9 dvss 1.17258f
C709 vg2.n10 dvss 0.244906f
C710 vg2.n11 dvss 0.522037f
C711 vg2.t7 dvss 0.628646f
C712 vg2.n12 dvss 0.313029f
C713 vg2.n13 dvss 0.32051f
C714 vg2.t8 dvss 0.505469f
C715 vg2.t2 dvss 39.125f
C716 vg2.t1 dvss 39.3426f
C717 vg2.t4 dvss 39.3426f
C718 vg2.t3 dvss 39.11f
C719 vg2.n15 dvss 9.00528f
C720 vg2.n16 dvss 2.91513f
C721 xin.n0 dvss 0.172822f
C722 xin.n5 dvss 0.184148f
C723 xin.t18 dvss 0.1922f
C724 xin.t15 dvss 0.19211f
C725 xin.n6 dvss 0.184148f
C726 xin.t13 dvss 0.19211f
C727 xin.t19 dvss 0.19211f
C728 xin.t16 dvss 0.19211f
C729 xin.t11 dvss 0.19211f
C730 xin.t10 dvss 0.19211f
C731 xin.t17 dvss 0.19211f
C732 xin.t14 dvss 0.19211f
C733 xin.t12 dvss 0.19211f
C734 xin.t9 dvss 0.19211f
C735 xin.t6 dvss 0.19211f
C736 xin.n21 dvss 0.175223f
C737 xin.n22 dvss 0.784969f
C738 xin.n23 dvss 0.308623f
C739 xin.n24 dvss 0.374761f
C740 xin.t20 dvss 0.828066f
C741 xin.t7 dvss 0.796281f
C742 xin.n25 dvss 0.514f
C743 xin.n26 dvss 0.386948f
C744 xin.n27 dvss 3.79487f
C745 xin.n28 dvss 4.5191f
C746 xin.n29 dvss 3.61279f
C747 xin.t1 dvss 57.0239f
C748 xin.t3 dvss 44.1862f
C749 xin.t0 dvss 44.012f
C750 xin.t5 dvss 0.124226f
C751 xin.n30 dvss 4.7746f
C752 xin.n31 dvss 27.2736f
C753 xin.t4 dvss 31.1925f
C754 xin.n32 dvss 27.266699f
C755 xin.t2 dvss 31.1614f
C756 xin.n33 dvss 27.270199f
C757 xin.n34 dvss 3.77704f
C758 xin.n35 dvss 1.85671f
C759 xin.n36 dvss 0.500575f
C760 vg1.n0 dvss 0.44953f
C761 vg1.t8 dvss 46.057503f
C762 vg1.t9 dvss 46.8352f
C763 vg1.t4 dvss 23.996801f
C764 vg1.n1 dvss 23.9575f
C765 vg1.t7 dvss 23.996801f
C766 vg1.n2 dvss 23.4861f
C767 vg1.t6 dvss 23.996801f
C768 vg1.n3 dvss 12.9859f
C769 vg1.n4 dvss 15.228601f
C770 vg1.n5 dvss 3.04049f
C771 vg1.n6 dvss 1.50262f
C772 vg1.t0 dvss 0.271659f
C773 vg1.t5 dvss 0.353472f
C774 vg1.n7 dvss 0.229145f
C775 vg1.n9 dvss 0.281876f
C776 vg1.n10 dvss 0.146945f
C777 vg1.n11 dvss 0.153437f
C778 vg1.n12 dvss 0.372304f
C779 x3.out_b.t6 dvss 0.402581f
C780 x3.out_b.n0 dvss 0.790285f
C781 x3.out_b.n1 dvss 1.5584f
C782 x3.out_b.n2 dvss 6.60541f
C783 x3.out_b.t4 dvss 0.420289f
C784 x3.out_b.n3 dvss 0.339622f
C785 x3.out_b.t7 dvss 0.402581f
C786 x3.out_b.n4 dvss 0.342378f
C787 x3.out_b.t8 dvss 0.420331f
C788 x3.out_b.n5 dvss 0.338349f
C789 x3.out_b.t3 dvss 0.402581f
C790 x3.out_b.n6 dvss 0.345348f
C791 x3.out_b.n7 dvss 0.58218f
C792 x3.out_b.t5 dvss 1.5189f
C793 x3.out_b.n8 dvss 0.163419f
C794 avdd.n0 dvss 0.492818f
C795 avdd.n1 dvss 1.6981f
C796 avdd.n4 dvss 0.266474f
C797 avdd.n5 dvss 0.585389f
C798 avdd.n6 dvss 1.03476f
C799 avdd.n7 dvss 1.03476f
C800 avdd.t17 dvss 0.894926f
C801 avdd.t11 dvss 0.702496f
C802 avdd.t4 dvss 0.894926f
C803 avdd.t0 dvss 0.702496f
C804 avdd.n8 dvss 0.46232f
C805 avdd.t14 dvss 7.53658f
C806 avdd.n9 dvss 7.5153f
C807 avdd.t13 dvss 9.12027f
C808 avdd.t16 dvss 7.25381f
C809 avdd.n10 dvss 7.71793f
C810 avdd.t15 dvss 9.163919f
C811 avdd.n11 dvss 3.68652f
C812 avdd.n12 dvss 0.768588f
C813 avdd.n13 dvss 0.579746f
C814 avdd.n14 dvss 0.560241f
C815 avdd.n15 dvss 0.353066f
C816 avdd.n16 dvss 0.487874f
C817 avdd.n17 dvss 3.7478f
C818 avdd.n18 dvss 0.731215f
C819 avdd.n21 dvss 1.93441f
C820 avdd.n22 dvss 0.967373f
C821 avdd.t18 dvss 0.135207f
C822 avdd.n23 dvss 0.34342f
C823 avdd.n24 dvss 5.68989f
C824 avdd.n25 dvss 1.05169f
C825 avdd.n26 dvss 1.1887f
C826 avdd.n27 dvss 1.1887f
C827 avdd.n28 dvss 4.46094f
C828 avdd.n29 dvss 1.35368f
C829 avdd.n32 dvss 0.548551f
C830 avdd.n33 dvss 1.56238f
C831 avdd.n34 dvss 1.46595f
C832 avdd.n35 dvss 0.107384f
C833 avdd.n36 dvss 0.107943f
C834 avdd.n37 dvss 0.158157f
C835 avdd.t2 dvss 2.51038f
C836 avdd.n39 dvss 0.10415f
C837 avdd.n40 dvss 0.107943f
C838 avdd.n41 dvss 0.559667f
C839 avdd.n43 dvss 0.687088f
C840 avdd.n44 dvss 1.48367f
C841 avdd.n45 dvss 1.13727f
C842 avdd.n46 dvss 0.744579f
C843 avdd.n47 dvss 2.46523f
C844 avdd.n48 dvss 3.43088f
C845 avdd.n49 dvss 1.15288f
C846 avdd.n50 dvss 0.362301f
C847 avdd.n51 dvss 0.321745f
C848 avdd.n52 dvss 0.106191f
C849 avdd.n53 dvss 1.67879f
C850 avdd.n54 dvss 0.106191f
C851 avdd.n55 dvss 0.158157f
C852 avdd.n58 dvss 0.106191f
C853 avdd.n59 dvss 1.67879f
C854 avdd.n60 dvss 0.106191f
C855 avdd.n62 dvss 0.116928f
C856 avdd.n63 dvss 0.719248f
C857 avdd.n64 dvss 1.37927f
C858 avdd.n65 dvss 1.47231f
C859 avdd.n66 dvss 1.45902f
C860 avdd.n67 dvss 0.366507f
C861 avdd.n68 dvss 0.107943f
C862 avdd.n69 dvss 0.158157f
C863 avdd.t6 dvss 2.51038f
C864 avdd.n70 dvss 0.10415f
C865 avdd.n71 dvss 0.107943f
C866 avdd.n72 dvss 0.107384f
C867 avdd.n74 dvss 0.106191f
C868 avdd.n75 dvss 1.67879f
C869 avdd.n76 dvss 0.106191f
C870 avdd.n77 dvss 0.158157f
C871 avdd.n78 dvss 0.106191f
C872 avdd.n79 dvss 1.67879f
C873 avdd.n80 dvss 0.106191f
C874 avdd.n81 dvss 0.319178f
C875 avdd.n82 dvss 0.73302f
C876 avdd.n83 dvss 1.95073f
C877 avdd.n84 dvss 4.13419f
C878 avdd.n85 dvss 0.707422f
C879 avdd.n86 dvss 0.479606f
C880 avdd.n87 dvss 1.32047f
C881 avdd.n88 dvss 1.35617f
C882 avdd.n89 dvss 0.536684f
C883 avdd.n90 dvss 1.19042f
C884 avdd.n91 dvss 4.48227f
C885 avdd.n92 dvss 4.46094f
C886 avdd.n93 dvss 4.48227f
C887 avdd.n94 dvss 1.19042f
C888 avdd.n95 dvss 0.66577f
C889 avdd.n96 dvss 3.27742f
C890 avdd.n97 dvss 0.20944f
C891 avdd.t9 dvss 0.702496f
C892 avdd.n98 dvss 0.20944f
C893 avdd.n99 dvss 0.731637f
C894 avdd.n100 dvss 0.757787f
C895 avdd.n101 dvss 0.146948f
C896 avdd.n103 dvss 0.303016f
C897 avss.n0 dvss 0.274689f
C898 avss.n1 dvss 0.256432f
C899 avss.n2 dvss 0.199691f
C900 avss.n4 dvss 0.10291f
C901 avss.t16 dvss 0.441575f
C902 avss.t14 dvss 0.441575f
C903 avss.n9 dvss 0.832446f
C904 avss.n10 dvss 0.117588f
C905 avss.n11 dvss 0.501337f
C906 avss.n15 dvss 0.506602f
C907 avss.n17 dvss 0.506602f
C908 avss.t0 dvss 0.441575f
C909 avss.n18 dvss 0.238935f
C910 avss.t2 dvss 0.441575f
C911 avss.n19 dvss 3.28532f
C912 avss.n20 dvss 7.3481f
C913 avss.t4 dvss 0.441575f
C914 avss.n24 dvss 0.152326f
C915 avss.n27 dvss 0.238935f
C916 avss.t6 dvss 0.441575f
C917 avss.n29 dvss 0.506602f
C918 avss.n30 dvss 0.506602f
C919 avss.t20 dvss 0.441575f
C920 avss.t22 dvss 0.441575f
C921 avss.n32 dvss 0.370586f
C922 avss.n33 dvss 0.325025f
C923 avss.n34 dvss 0.132878f
C924 avss.n35 dvss 0.404741f
C925 avss.n36 dvss 2.98049f
C926 avss.t12 dvss 0.860518f
C927 avss.t8 dvss 0.732948f
C928 avss.n37 dvss 2.16357f
C929 avss.n38 dvss 1.84584f
C930 avss.t10 dvss 0.841962f
C931 avss.t18 dvss 0.732948f
C932 avss.n39 dvss 0.3741f
C933 avss.n40 dvss 0.133098f
C934 avss.t24 dvss 0.732948f
C935 avss.n41 dvss 0.133098f
C936 avss.n42 dvss 1.68799f
C937 avss.n43 dvss 0.462717f
C938 avss.n46 dvss 1.36147f
C939 avss.n47 dvss 1.03577f
C940 avss.t26 dvss 8.17429f
C941 avss.n48 dvss 7.701231f
C942 avss.t29 dvss 8.17429f
C943 avss.n49 dvss 8.01034f
C944 avss.t28 dvss 8.17429f
C945 avss.n50 dvss 7.90618f
C946 avss.n51 dvss 4.01706f
C947 avss.t27 dvss 8.17429f
C948 avss.n52 dvss 2.18128f
C949 avss.n53 dvss 4.97729f
C950 avss.n54 dvss 1.85282f
C951 avss.n55 dvss 1.94389f
C952 avss.n56 dvss 1.85115f
C953 avss.n58 dvss 0.227287f
C954 avss.n59 dvss 0.265186f
C955 avss.n60 dvss 0.643717f
C956 avss.n61 dvss 0.274689f
C957 avss.n62 dvss 0.354568f
C958 avss.n64 dvss 0.102951f
C959 avss.n68 dvss 0.238935f
C960 avss.n71 dvss 0.10291f
C961 avss.n73 dvss 0.117505f
C962 avss.n75 dvss 0.79544f
C963 avss.n76 dvss 1.9882f
C964 avss.n77 dvss 0.79544f
C965 avss.n79 dvss 0.117505f
C966 avss.n80 dvss 0.117588f
C967 avss.n81 dvss 0.455799f
C968 avss.n82 dvss 1.20688f
C969 avss.n83 dvss 0.606761f
C970 avss.n84 dvss 0.354568f
C971 avss.n86 dvss 0.102951f
C972 avss.n89 dvss 0.238935f
C973 avss.n92 dvss 0.152326f
C974 avss.n94 dvss 0.162188f
C975 avss.n95 dvss 0.241706f
C976 x7.x1.clkin dvss 0.290534f
C977 x7.x2.clkin dvss 0.174689f
C978 dout_ip.n0 dvss 3.72627f
C979 x7.clkin dvss 5.05976f
C980 dout_ip.n6 dvss 0.35872f
C981 dout_ip.n7 dvss 0.352547f
C982 inv_in.t3 dvss 0.657711f
C983 inv_in.t11 dvss 5.68012f
C984 inv_in.n0 dvss 5.17707f
C985 inv_in.t5 dvss 5.52894f
C986 inv_in.n1 dvss 2.62426f
C987 inv_in.t6 dvss 5.52894f
C988 inv_in.n2 dvss 2.66147f
C989 inv_in.n3 dvss 2.79669f
C990 inv_in.t14 dvss 5.52894f
C991 inv_in.n4 dvss 5.29306f
C992 inv_in.t12 dvss 5.55261f
C993 inv_in.n5 dvss 5.28615f
C994 inv_in.t13 dvss 5.52894f
C995 inv_in.n6 dvss 2.66147f
C996 inv_in.t9 dvss 5.5836f
C997 inv_in.n7 dvss 5.39875f
C998 inv_in.t10 dvss 5.5836f
C999 inv_in.t2 dvss 5.5836f
C1000 inv_in.n8 dvss 5.26653f
C1001 inv_in.n9 dvss 5.40864f
C1002 inv_in.t4 dvss 5.52894f
C1003 inv_in.n10 dvss 2.66147f
C1004 inv_in.n11 dvss 2.90209f
C1005 inv_in.n12 dvss 2.75998f
C1006 inv_in.t8 dvss 5.52894f
C1007 inv_in.n13 dvss 2.62426f
C1008 inv_in.n14 dvss 2.76492f
C1009 inv_in.n15 dvss 2.76492f
C1010 inv_in.n16 dvss 2.76201f
C1011 inv_in.t7 dvss 5.52894f
C1012 inv_in.n17 dvss 5.4592f
C1013 inv_in.n18 dvss 0.82306f
C1014 inv_in.t0 dvss 0.104143f
C1015 inv_in.t1 dvss 0.647866f
C1016 inv_in.n19 dvss 2.16816f
C1017 xout.t18 dvss 0.243993f
C1018 xout.t16 dvss 0.243993f
C1019 xout.n0 dvss 2.4243f
C1020 xout.t17 dvss 0.243993f
C1021 xout.t15 dvss 0.243993f
C1022 xout.n1 dvss 1.60432f
C1023 xout.n2 dvss 6.32987f
C1024 xout.t14 dvss 0.256529f
C1025 xout.t19 dvss 0.243993f
C1026 xout.n3 dvss 1.22843f
C1027 xout.t12 dvss 0.256529f
C1028 xout.t20 dvss 0.243993f
C1029 xout.n4 dvss 1.23308f
C1030 xout.n5 dvss 2.18555f
C1031 xout.n6 dvss 8.527769f
C1032 xout.n7 dvss 3.77761f
C1033 xout.t9 dvss 0.243993f
C1034 xout.t10 dvss 0.243993f
C1035 xout.n8 dvss 1.27442f
C1036 xout.n9 dvss 1.83376f
C1037 xout.t11 dvss 0.243993f
C1038 xout.t13 dvss 0.243993f
C1039 xout.n10 dvss 1.43377f
C1040 xout.n11 dvss 1.68066f
C1041 xout.n12 dvss 1.24537f
C1042 xout.n13 dvss 0.227228f
C1043 xout.n14 dvss 0.217681f
C1044 xout.n15 dvss 0.229174f
C1045 xout.n16 dvss 4.49086f
C1046 xout.n17 dvss 0.217681f
C1047 xout.n18 dvss 0.149204f
C1048 xout.n19 dvss 2.97025f
C1049 xout.n20 dvss 3.47714f
C1050 xout.n21 dvss 4.15788f
C1051 xout.n22 dvss 4.02374f
C1052 xout.n23 dvss 0.626416f
C1053 xout.n24 dvss 0.760656f
C1054 xout.t25 dvss 1.61622f
C1055 xout.t23 dvss 1.68073f
C1056 xout.n25 dvss 1.04327f
C1057 xout.n26 dvss 0.785936f
C1058 xout.n27 dvss 8.087669f
C1059 xout.n28 dvss 9.65943f
C1060 xout.n29 dvss 1.9924f
C1061 avdd_ip.n0 dvss 0.183001f
C1062 avdd_ip.n1 dvss 0.193101f
C1063 avdd_ip.t1 dvss 0.312571f
C1064 avdd_ip.n2 dvss 25.687199f
C1065 avdd_ip.t33 dvss 0.201546p
C1066 avdd_ip.n3 dvss 42.3367f
C1067 avdd_ip.n4 dvss 31.209301f
C1068 avdd_ip.t30 dvss 12.6155f
C1069 avdd_ip.n5 dvss 8.054391f
C1070 avdd_ip.t31 dvss 12.6155f
C1071 avdd_ip.n6 dvss 7.765079f
C1072 avdd_ip.n7 dvss 10.2323f
C1073 avdd_ip.t29 dvss 12.6155f
C1074 avdd_ip.n8 dvss 11.3223f
C1075 avdd_ip.t32 dvss 12.6155f
C1076 avdd_ip.n9 dvss 11.2988f
C1077 avdd_ip.n10 dvss 11.0453f
C1078 avdd_ip.n11 dvss 25.8585f
C1079 avdd_ip.n12 dvss 11.8125f
C1080 avdd_ip.n13 dvss 15.647901f
C1081 avdd_ip.t20 dvss 0.272851f
C1082 avdd_ip.n14 dvss 0.353227f
C1083 avdd_ip.t24 dvss 0.272851f
C1084 avdd_ip.n15 dvss 1.24555f
C1085 avdd_ip.t25 dvss 0.272851f
C1086 avdd_ip.n16 dvss 1.36471f
C1087 avdd_ip.t23 dvss 0.284354f
C1088 avdd_ip.n17 dvss 1.00481f
C1089 avdd_ip.n18 dvss 1.60279f
C1090 avdd_ip.n19 dvss 0.908877f
C1091 avdd_ip.n20 dvss 0.312041f
C1092 avdd_ip.t21 dvss 0.272851f
C1093 avdd_ip.n21 dvss 0.511759f
C1094 avdd_ip.n22 dvss 1.0293f
C1095 avdd_ip.n23 dvss 1.19091f
C1096 avdd_ip.t19 dvss 0.272851f
C1097 avdd_ip.n24 dvss 1.06873f
C1098 avdd_ip.n25 dvss 4.33929f
C1099 avdd_ip.n26 dvss 15.187299f
C1100 avdd_ip.n27 dvss 15.187299f
C1101 avdd_ip.t6 dvss 19.331099f
C1102 avdd_ip.n28 dvss 1.61496f
C1103 avdd_ip.t11 dvss 0.272851f
C1104 avdd_ip.n29 dvss 5.41016f
C1105 avdd_ip.t16 dvss 0.272851f
C1106 avdd_ip.t17 dvss 0.272851f
C1107 avdd_ip.n30 dvss 2.76186f
C1108 avdd_ip.t13 dvss 0.272851f
C1109 avdd_ip.t15 dvss 0.272851f
C1110 avdd_ip.n31 dvss 1.60468f
C1111 avdd_ip.n32 dvss 2.4602f
C1112 avdd_ip.n33 dvss 6.7614f
C1113 avdd_ip.n40 dvss 0.275331f
C1114 avdd_ip.t2 dvss 0.366056f
C1115 avdd_ip.n42 dvss -24.5529f
C1116 avdd_ip.n43 dvss 24.8309f
C1117 avdd_ip.n47 dvss 2.63147f
C1118 avdd_ip.t5 dvss 0.425863f
C1119 avdd_ip.n54 dvss 0.275331f
C1120 avdd_ip.n57 dvss 0.275331f
C1121 avdd_ip.n60 dvss 2.34174f
C1122 avdd_ip.n61 dvss 3.08369f
C1123 avdd_ip.n62 dvss 7.458549f
C1124 avdd_ip.t7 dvss 0.272851f
C1125 avdd_ip.t8 dvss 0.272851f
C1126 avdd_ip.t9 dvss 0.272851f
C1127 avdd_ip.n63 dvss 2.28083f
C1128 avdd_ip.t22 dvss 0.272851f
C1129 avdd_ip.t27 dvss 0.272851f
C1130 avdd_ip.n64 dvss 2.68748f
C1131 avdd_ip.t18 dvss 0.272851f
C1132 avdd_ip.t26 dvss 0.272851f
C1133 avdd_ip.n65 dvss 1.60335f
C1134 avdd_ip.n66 dvss 2.5326f
C1135 avdd_ip.n67 dvss 6.54556f
C1136 avdd_ip.n68 dvss 5.37955f
C1137 avdd_ip.n69 dvss 12.5401f
C1138 avdd_ip.n70 dvss 7.683919f
C1139 avdd_ip.n71 dvss 8.52327f
C1140 avdd_ip.n72 dvss 8.52327f
C1141 avdd_ip.n73 dvss 32.6198f
C1142 avdd_ip.n74 dvss 7.0648f
C1143 avdd_ip.n75 dvss 2.67542f
C1144 avdd_ip.n76 dvss 5.79729f
C1145 avdd_ip.n77 dvss 37.3139f
C1146 avdd_ip.n78 dvss 13.6449f
C1147 avdd_ip.n79 dvss 32.799896f
C1148 avdd_ip.n80 dvss 32.6198f
C1149 avdd_ip.n81 dvss 32.799896f
C1150 avdd_ip.n82 dvss 8.53496f
C1151 avdd_ip.n83 dvss 8.47481f
C1152 avdd_ip.n84 dvss 3.99638f
C1153 avdd_ip.n85 dvss 32.939102f
C1154 avdd_ip.n86 dvss 7.89575f
C1155 avdd_ip.n87 dvss 2.20457f
C1156 avdd_ip.n88 dvss 5.76955f
C1157 avdd_ip.t12 dvss 0.272851f
C1158 avdd_ip.t14 dvss 0.272851f
C1159 avdd_ip.n89 dvss 2.2737f
C1160 avdd_ip.n90 dvss 0.777352f
C1161 avdd_ip.n91 dvss 1.40119f
C1162 avdd_ip.t10 dvss 19.331099f
C1163 avdd_ip.n92 dvss 16.5454f
C1164 avdd_ip.n93 dvss 1.40119f
C1165 avdd_ip.n94 dvss 2.89537f
C1166 avdd_ip.n95 dvss 1.66736f
C1167 avdd_ip.n96 dvss 7.11433f
C1168 avdd_ip.n97 dvss 23.7224f
C1169 ibias_ip.n0 dvss 4.75326f
C1170 ibias_ip.n1 dvss 0.974101f
C1171 ibias_ip.t13 dvss 0.653909f
C1172 ibias_ip.t2 dvss 0.646782f
C1173 ibias_ip.t6 dvss 0.644915f
C1174 ibias_ip.t0 dvss 0.650434f
C1175 ibias_ip.t4 dvss 0.647233f
C1176 ibias_ip.t11 dvss 0.653916f
C1177 ibias_ip.t8 dvss 0.645067f
C1178 ibias_ip.t12 dvss 0.646314f
C1179 ibias_ip.t10 dvss 0.184945f
C1180 standby_33.n0 dvss 7.3102f
C1181 standby_33.t3 dvss 0.80334f
C1182 standby_33.t4 dvss 1.62318f
C1183 standby_33.n1 dvss 0.174581f
C1184 x7.ena_done_b.n7 dvss 1.96309f
C1185 a_9120_n9346.t0 dvss 1.47746f
C1186 a_9120_n9346.n0 dvss 3.32132f
C1187 a_9120_n9346.t2 dvss 1.67898f
C1188 a_9120_n9346.n1 dvss 2.97825f
C1189 a_9120_n9346.n2 dvss 1.80939f
C1190 x7.x2.x4.RESET_B dvss 1.471743f
C1191 standby_b.n0 dvss 0.153287f
C1192 x4.in_b dvss 2.69011f
C1193 standby_b.n1 dvss 3.12348f
C1194 x7.stby_b dvss 1.34845f
C1195 standby_b.t12 dvss 0.182513f
C1196 standby_b.t4 dvss 0.182371f
C1197 standby_b.n3 dvss 0.157601f
C1198 standby_b.t19 dvss 0.228815f
C1199 standby_b.t17 dvss 0.217171f
C1200 standby_b.n4 dvss 0.157601f
C1201 standby_b.t7 dvss 0.217171f
C1202 standby_b.t23 dvss 0.217171f
C1203 standby_b.t21 dvss 0.217171f
C1204 standby_b.n11 dvss 0.162102f
C1205 standby_b.t6 dvss 0.229503f
C1206 standby_b.t16 dvss 0.217171f
C1207 standby_b.n12 dvss 0.161693f
C1208 standby_b.t18 dvss 0.217171f
C1209 standby_b.t0 dvss 0.217171f
C1210 standby_b.t3 dvss 0.217171f
C1211 tail.n0 dvss 0.76343f
C1212 tail.n1 dvss 2.82244f
C1213 tail.n2 dvss 0.753923f
C1214 tail.n3 dvss 0.119757f
C1215 tail.t0 dvss 0.102772f
C1216 tail.t5 dvss 0.102893f
C1217 tail.t7 dvss 0.102832f
C1218 tail.t2 dvss 0.102832f
C1219 tail.t4 dvss 0.103102f
C1220 tail.t9 dvss 0.102562f
C1221 tail.t3 dvss 0.103102f
C1222 tail.t8 dvss 0.102562f
C1223 tail.t6 dvss 0.102998f
C1224 tail.t1 dvss 0.102668f
C1225 vbp.n0 dvss 0.179072f
C1226 vbp.n1 dvss 0.347213f
C1227 vbp.n2 dvss 0.361375f
C1228 vbp.n3 dvss 6.70539f
C1229 vbp.n4 dvss 0.178688f
C1230 vbp.n5 dvss 0.347213f
C1231 vbp.n6 dvss 0.345626f
C1232 vbp.n7 dvss 0.353693f
C1233 vbp.t13 dvss 0.876014f
C1234 vbp.t5 dvss 0.946258f
C1235 vbp.t1 dvss 0.114991f
C1236 vbp.t9 dvss 0.880979f
C1237 vbp.t7 dvss 0.853138f
C1238 vbp.t12 dvss 0.876026f
C1239 vbp.t17 dvss 0.946667f
C1240 vbp.t11 dvss 1.12602f
C1241 vbp.t14 dvss 0.854726f
C1242 vbp.t4 dvss 0.854724f
C1243 vbp.t0 dvss 0.908023f
C1244 vbp.t15 dvss 1.12462f
C1245 vbp.t8 dvss 0.853138f
C1246 vbp.t16 dvss 0.891507f
C1247 vbp.t6 dvss 0.891734f
C1248 vbp.t10 dvss 0.871833f
C1249 vbp.t3 dvss 0.8852f
C1250 vbp.t2 dvss 0.123277f
C1251 vbreg.n0 dvss 3.5606f
C1252 vbreg.n1 dvss 0.713612f
C1253 vbreg.n2 dvss 0.583542f
C1254 vbreg.n3 dvss 3.65749f
C1255 vbreg.n4 dvss 1.34473f
C1256 vbreg.n5 dvss 3.556f
C1257 vbreg.n6 dvss 0.687636f
C1258 vbreg.n7 dvss 0.582626f
C1259 vbreg.n8 dvss 1.213f
C1260 vbreg.n9 dvss 2.841f
C1261 vbreg.n10 dvss 0.583359f
C1262 vbreg.n11 dvss 2.61721f
C1263 vbreg.n12 dvss 0.592924f
C1264 vbreg.n14 dvss 0.594449f
C1265 vbreg.n15 dvss 0.931401f
C1266 vbreg.n16 dvss 0.933049f
C1267 vbreg.n17 dvss 0.404251f
C1268 vbreg.n18 dvss 0.933049f
C1269 vbreg.t11 dvss 1.20117f
C1270 vbreg.n19 dvss 0.931401f
C1271 vbreg.t2 dvss 0.23921f
C1272 vbreg.n20 dvss 1.79539f
C1273 vbreg.n21 dvss 12.184299f
C1274 vbreg.t4 dvss 0.228907f
C1275 vbreg.n22 dvss 1.25884f
C1276 vbreg.n23 dvss 0.616431f
C1277 vbreg.t7 dvss 1.20117f
C1278 vbreg.n24 dvss 0.662505f
C1279 vbreg.t19 dvss 1.20117f
C1280 vbreg.n25 dvss 0.404251f
C1281 vbreg.n26 dvss 0.400957f
C1282 vbreg.t20 dvss 1.20117f
C1283 vbreg.t18 dvss 1.20117f
C1284 vbreg.t15 dvss 1.20117f
C1285 vbreg.n27 dvss 1.00001f
C1286 vbreg.t16 dvss 1.20117f
C1287 vbreg.n28 dvss 0.685977f
C1288 vbreg.n29 dvss 0.530447f
C1289 vbreg.n30 dvss 0.404251f
C1290 vbreg.n31 dvss 0.710975f
C1291 vbreg.t10 dvss 1.21612f
C1292 vbreg.t13 dvss 1.20117f
C1293 vbreg.n32 dvss 1.00001f
C1294 vbreg.t12 dvss 1.20117f
C1295 vbreg.n34 dvss 1.00001f
C1296 vbreg.t14 dvss 1.20117f
C1297 vbreg.n35 dvss 0.692695f
C1298 vbreg.n36 dvss 1.00001f
C1299 vbreg.t9 dvss 1.20117f
C1300 vbreg.n37 dvss 0.530447f
C1301 vbreg.n38 dvss 0.661796f
C1302 vbreg.t17 dvss 1.20117f
C1303 vbreg.n39 dvss 1.00001f
C1304 vbreg.n40 dvss 0.168268f
C1305 vbreg.n41 dvss 1.00001f
C1306 vbreg.t8 dvss 0.228404f
C1307 vbreg.n42 dvss 0.81533f
C1308 vbreg.n43 dvss 0.528798f
C1309 vbreg.n44 dvss 0.404251f
C1310 vbreg.n45 dvss 1.00001f
C1311 vbreg.t22 dvss 1.20117f
C1312 vbreg.t24 dvss 1.20117f
C1313 vbreg.t25 dvss 1.20117f
C1314 vbreg.n46 dvss 1.00001f
C1315 vbreg.t21 dvss 1.20117f
C1316 vbreg.n47 dvss 0.531546f
C1317 vbreg.t23 dvss 1.21618f
C1318 vbreg.n48 dvss 1.00001f
C1319 vbreg.n50 dvss 1.30967f
C1320 vbreg.n51 dvss 0.705365f
C1321 vbreg.n52 dvss 0.531546f
C1322 vbreg.n53 dvss 0.404251f
C1323 vbreg.n54 dvss 0.527699f
C1324 vbreg.n55 dvss 0.527699f
C1325 vbreg.n56 dvss 0.404251f
C1326 vbreg.n57 dvss 0.55298f
C1327 vbreg.t6 dvss 0.214967f
C1328 vbreg.t3 dvss 0.228223f
C1329 vbreg.t1 dvss 0.268952f
C1330 vbreg.t5 dvss 0.218294f
C1331 vbreg.t0 dvss 0.138373f
C1332 icnode.t1 dvss 80.4574f
C1333 dvdd.n0 dvss 0.231928f
C1334 dvdd.n4 dvss 0.114981f
C1335 dvdd.n5 dvss 0.114981f
C1336 dvdd.n27 dvss 0.114981f
C1337 dvdd.n29 dvss 0.114981f
C1338 dvdd.t12 dvss 0.165457f
C1339 dvdd.n38 dvss 0.47343f
C1340 dvdd.n39 dvss 0.249961f
C1341 dvdd.t48 dvss 0.165457f
C1342 dvdd.n49 dvss 1.8472f
C1343 dvdd.t175 dvss 3.83628f
C1344 dvdd.n50 dvss 3.2293f
C1345 dvdd.n51 dvss 1.13209f
C1346 dvdd.t134 dvss 0.103953f
C1347 dvdd.t56 dvss 0.103953f
C1348 dvdd.t157 dvss 0.103953f
C1349 dvdd.n275 dvss 6.53977f
C1350 dvdd.n276 dvss 9.40408f
C1351 dvdd.t178 dvss 3.83628f
C1352 dvdd.n277 dvss 6.79779f
C1353 dvdd.t177 dvss 3.83628f
C1354 dvdd.n278 dvss 3.72992f
C1355 dvdd.t176 dvss 3.83628f
C1356 dvdd.n279 dvss 3.60793f
C1357 dvdd.n280 dvss 2.57602f
C1358 dvdd.n281 dvss 0.390563f
C1359 dvdd.n290 dvss 0.466107f
C1360 dvdd.n291 dvss 0.869136f
C1361 dvdd.n292 dvss 0.243102f
C1362 dvdd.n293 dvss 0.211035f
C1363 dvdd.t14 dvss 0.222917f
C1364 dvdd.t20 dvss 0.187598f
C1365 dvdd.t22 dvss 0.187598f
C1366 dvdd.t16 dvss 0.187598f
C1367 dvdd.t18 dvss 0.140698f
C1368 dvdd.t26 dvss 0.140698f
C1369 dvdd.t8 dvss 0.187598f
C1370 dvdd.t10 dvss 0.187598f
C1371 dvdd.t24 dvss 0.187598f
C1372 dvdd.t28 dvss 0.222917f
C1373 dvdd.n295 dvss 0.211035f
C1374 dvdd.n296 dvss 0.255981f
C1375 dvdd.n297 dvss 0.773905f
C1376 dvdd.n298 dvss 0.37474f
.ends

