magic
tech sky130A
magscale 1 2
timestamp 1712203273
<< dnwell >>
rect 2208 -2310 5968 238
<< nwell >>
rect 2128 32 6048 318
rect 2128 -2104 2414 32
rect 5762 -2104 6048 32
rect 2128 -2390 6048 -2104
<< nsubdiff >>
rect 2165 261 6011 281
rect 2165 227 2245 261
rect 5931 227 6011 261
rect 2165 207 6011 227
rect 2165 201 2239 207
rect 2165 -2273 2185 201
rect 2219 -2273 2239 201
rect 2165 -2279 2239 -2273
rect 5937 201 6011 207
rect 5937 -2273 5957 201
rect 5991 -2273 6011 201
rect 5937 -2279 6011 -2273
rect 2165 -2299 6011 -2279
rect 2165 -2333 2245 -2299
rect 5931 -2333 6011 -2299
rect 2165 -2353 6011 -2333
<< nsubdiffcont >>
rect 2245 227 5931 261
rect 2185 -2273 2219 201
rect 5957 -2273 5991 201
rect 2245 -2333 5931 -2299
<< locali >>
rect 2185 227 2245 261
rect 5931 227 5991 261
rect 2185 201 2219 227
rect 2185 -2299 2219 -2273
rect 5957 201 5991 227
rect 5957 -2299 5991 -2273
rect 2185 -2333 2245 -2299
rect 5931 -2333 5991 -2299
<< metal1 >>
rect 4538 110 4738 310
rect 920 -302 1120 -102
rect 5846 -306 6046 -106
rect 590 -1134 790 -934
rect 958 -1548 1060 -534
rect 1136 -1014 1192 -614
rect 1136 -1082 1396 -1014
rect 1136 -1472 1192 -1082
rect 898 -2018 1098 -1818
rect 5848 -2000 6048 -1800
rect 1744 -2360 1944 -2160
rect 3112 -2358 3312 -2158
use sky130_fd_pr__nfet_01v8_69TQ3K  XM1
timestamp 1712071977
transform -1 0 1010 0 -1 -1374
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_3HMWVM  XM2
timestamp 1712071977
transform -1 0 1010 0 -1 -715
box -296 -319 296 319
use sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B  XM3
timestamp 1712071977
transform 0 1 3236 -1 0 -687
box -357 -558 357 558
use sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B  XM4
timestamp 1712071977
transform 0 1 3236 -1 0 -1393
box -357 -558 357 558
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM5
timestamp 1712071977
transform 0 1 4339 -1 0 -1040
box -658 -397 658 397
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM6
timestamp 1712071977
transform 0 1 4943 -1 0 -1040
box -658 -397 658 397
<< labels >>
flabel metal1 5848 -2000 6048 -1800 0 FreeSans 128 0 0 0 out
port 2 nsew
flabel metal1 5846 -306 6046 -106 0 FreeSans 128 0 0 0 out_b
port 3 nsew
flabel metal1 4538 110 4738 310 0 FreeSans 128 0 0 0 avdd
port 0 nsew
flabel metal1 3112 -2358 3312 -2158 0 FreeSans 128 0 0 0 avss
port 6 nsew
flabel metal1 1744 -2360 1944 -2160 0 FreeSans 128 0 0 0 in_b
port 7 nsew
flabel metal1 590 -1134 790 -934 0 FreeSans 128 0 0 0 in
port 4 nsew
flabel metal1 920 -302 1120 -102 0 FreeSans 128 0 0 0 dvdd
port 1 nsew
flabel metal1 898 -2018 1098 -1818 0 FreeSans 128 0 0 0 dvss
port 5 nsew
<< end >>
