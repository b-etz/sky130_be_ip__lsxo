magic
tech sky130A
magscale 1 2
timestamp 1712851378
<< metal3 >>
rect -1492 4172 -120 4200
rect -1492 148 -204 4172
rect -140 148 -120 4172
rect -1492 120 -120 148
rect 120 4172 1492 4200
rect 120 148 1408 4172
rect 1472 148 1492 4172
rect 120 120 1492 148
rect -1492 -148 -120 -120
rect -1492 -4172 -204 -148
rect -140 -4172 -120 -148
rect -1492 -4200 -120 -4172
rect 120 -148 1492 -120
rect 120 -4172 1408 -148
rect 1472 -4172 1492 -148
rect 120 -4200 1492 -4172
<< via3 >>
rect -204 148 -140 4172
rect 1408 148 1472 4172
rect -204 -4172 -140 -148
rect 1408 -4172 1472 -148
<< mimcap >>
rect -1452 4120 -452 4160
rect -1452 200 -1412 4120
rect -492 200 -452 4120
rect -1452 160 -452 200
rect 160 4120 1160 4160
rect 160 200 200 4120
rect 1120 200 1160 4120
rect 160 160 1160 200
rect -1452 -200 -452 -160
rect -1452 -4120 -1412 -200
rect -492 -4120 -452 -200
rect -1452 -4160 -452 -4120
rect 160 -200 1160 -160
rect 160 -4120 200 -200
rect 1120 -4120 1160 -200
rect 160 -4160 1160 -4120
<< mimcapcontact >>
rect -1412 200 -492 4120
rect 200 200 1120 4120
rect -1412 -4120 -492 -200
rect 200 -4120 1120 -200
<< metal4 >>
rect -1004 4121 -900 4320
rect -224 4172 -120 4320
rect -1413 4120 -491 4121
rect -1413 200 -1412 4120
rect -492 200 -491 4120
rect -1413 199 -491 200
rect -1004 -199 -900 199
rect -224 148 -204 4172
rect -140 148 -120 4172
rect 608 4121 712 4320
rect 1388 4172 1492 4320
rect 199 4120 1121 4121
rect 199 200 200 4120
rect 1120 200 1121 4120
rect 199 199 1121 200
rect -224 -148 -120 148
rect -1413 -200 -491 -199
rect -1413 -4120 -1412 -200
rect -492 -4120 -491 -200
rect -1413 -4121 -491 -4120
rect -1004 -4320 -900 -4121
rect -224 -4172 -204 -148
rect -140 -4172 -120 -148
rect 608 -199 712 199
rect 1388 148 1408 4172
rect 1472 148 1492 4172
rect 1388 -148 1492 148
rect 199 -200 1121 -199
rect 199 -4120 200 -200
rect 1120 -4120 1121 -200
rect 199 -4121 1121 -4120
rect -224 -4320 -120 -4172
rect 608 -4320 712 -4121
rect 1388 -4172 1408 -148
rect 1472 -4172 1492 -148
rect 1388 -4320 1492 -4172
<< properties >>
string FIXED_BBOX 120 120 1200 4200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5 l 20 val 209.5 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
