magic
tech sky130A
magscale 1 2
timestamp 1712073863
<< metal3 >>
rect -7398 4572 -2626 4600
rect -7398 148 -2710 4572
rect -2646 148 -2626 4572
rect -7398 120 -2626 148
rect -2386 4572 2386 4600
rect -2386 148 2302 4572
rect 2366 148 2386 4572
rect -2386 120 2386 148
rect 2626 4572 7398 4600
rect 2626 148 7314 4572
rect 7378 148 7398 4572
rect 2626 120 7398 148
rect -7398 -148 -2626 -120
rect -7398 -4572 -2710 -148
rect -2646 -4572 -2626 -148
rect -7398 -4600 -2626 -4572
rect -2386 -148 2386 -120
rect -2386 -4572 2302 -148
rect 2366 -4572 2386 -148
rect -2386 -4600 2386 -4572
rect 2626 -148 7398 -120
rect 2626 -4572 7314 -148
rect 7378 -4572 7398 -148
rect 2626 -4600 7398 -4572
<< via3 >>
rect -2710 148 -2646 4572
rect 2302 148 2366 4572
rect 7314 148 7378 4572
rect -2710 -4572 -2646 -148
rect 2302 -4572 2366 -148
rect 7314 -4572 7378 -148
<< mimcap >>
rect -7358 4520 -2958 4560
rect -7358 200 -7318 4520
rect -2998 200 -2958 4520
rect -7358 160 -2958 200
rect -2346 4520 2054 4560
rect -2346 200 -2306 4520
rect 2014 200 2054 4520
rect -2346 160 2054 200
rect 2666 4520 7066 4560
rect 2666 200 2706 4520
rect 7026 200 7066 4520
rect 2666 160 7066 200
rect -7358 -200 -2958 -160
rect -7358 -4520 -7318 -200
rect -2998 -4520 -2958 -200
rect -7358 -4560 -2958 -4520
rect -2346 -200 2054 -160
rect -2346 -4520 -2306 -200
rect 2014 -4520 2054 -200
rect -2346 -4560 2054 -4520
rect 2666 -200 7066 -160
rect 2666 -4520 2706 -200
rect 7026 -4520 7066 -200
rect 2666 -4560 7066 -4520
<< mimcapcontact >>
rect -7318 200 -2998 4520
rect -2306 200 2014 4520
rect 2706 200 7026 4520
rect -7318 -4520 -2998 -200
rect -2306 -4520 2014 -200
rect 2706 -4520 7026 -200
<< metal4 >>
rect -5210 4521 -5106 4720
rect -2730 4572 -2626 4720
rect -7319 4520 -2997 4521
rect -7319 200 -7318 4520
rect -2998 200 -2997 4520
rect -7319 199 -2997 200
rect -5210 -199 -5106 199
rect -2730 148 -2710 4572
rect -2646 148 -2626 4572
rect -198 4521 -94 4720
rect 2282 4572 2386 4720
rect -2307 4520 2015 4521
rect -2307 200 -2306 4520
rect 2014 200 2015 4520
rect -2307 199 2015 200
rect -2730 -148 -2626 148
rect -7319 -200 -2997 -199
rect -7319 -4520 -7318 -200
rect -2998 -4520 -2997 -200
rect -7319 -4521 -2997 -4520
rect -5210 -4720 -5106 -4521
rect -2730 -4572 -2710 -148
rect -2646 -4572 -2626 -148
rect -198 -199 -94 199
rect 2282 148 2302 4572
rect 2366 148 2386 4572
rect 4814 4521 4918 4720
rect 7294 4572 7398 4720
rect 2705 4520 7027 4521
rect 2705 200 2706 4520
rect 7026 200 7027 4520
rect 2705 199 7027 200
rect 2282 -148 2386 148
rect -2307 -200 2015 -199
rect -2307 -4520 -2306 -200
rect 2014 -4520 2015 -200
rect -2307 -4521 2015 -4520
rect -2730 -4720 -2626 -4572
rect -198 -4720 -94 -4521
rect 2282 -4572 2302 -148
rect 2366 -4572 2386 -148
rect 4814 -199 4918 199
rect 7294 148 7314 4572
rect 7378 148 7398 4572
rect 7294 -148 7398 148
rect 2705 -200 7027 -199
rect 2705 -4520 2706 -200
rect 7026 -4520 7027 -200
rect 2705 -4521 7027 -4520
rect 2282 -4720 2386 -4572
rect 4814 -4720 4918 -4521
rect 7294 -4572 7314 -148
rect 7378 -4572 7398 -148
rect 7294 -4720 7398 -4572
<< properties >>
string FIXED_BBOX 2626 120 7106 4600
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 22 l 22 val 984.72 carea 2.00 cperi 0.19 nx 3 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
