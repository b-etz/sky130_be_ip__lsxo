* PEX produced on Mon Apr 15 19:45:33 EDT 2024 using /home/brady/sources/osic-multitool-src/iic-pex.sh with m=3 and s=1
* NGSPICE file created from sky130_be_ip__lsxo.ext - technology: sky130A

.subckt sky130_be_ip__lsxo ibias dout xout xin ena avss avdd standby dvss dvdd
X0 a_16620_n1869.t1 a_15705_n2241.t2 a_16273_n2273.t1 dvss.t122 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1 a_20376_n2791.t1 x7.stby_done_b.t2 dvdd.t140 dvdd.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_21036_n1869.t3 a_19955_n2241.t2 a_20689_n2273.t2 dvdd.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3 a_10620_n8338.t0 a_24220_n8172.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X4 a_16795_n2817.t1 a_16620_n2791.t4 a_16974_n2791.t1 dvss.t152 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5 dvdd.t37 ena_ip.t2 x3.in_b.t0 dvdd.t36 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X6 dvdd.t87 a_21036_n1869.t4 a_21211_n1943.t2 dvdd.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_18828_n2791.t2 a_17913_n2791.t2 a_18481_n2549.t3 dvss.t135 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X8 a_2130_n19848.t1 a_24530_n20014.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X9 vbreg.t2 icnode.t1 a_11526_n12394.t1 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X10 x7.x2.x2.CLK.t1 a_15000_n2791.t3 dvss.t186 dvss.t185 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X11 a_18168_n1881.t1 x7.x1.Qb2.t2 dvss.t114 dvss.t113 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X12 tail.t11 vbp.t3 dvdd_ip.t52 dvdd_ip.t42 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X13 a_16317_n2791.t0 a_16273_n2549.t4 a_16151_n2791.t0 dvss.t21 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X14 dvss.t200 standby_b.t2 dvss_ip dvss.t199 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X15 a_9120_n9346.t0 a_24220_n9832.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X16 a_16795_n1943.t1 a_16620_n1869.t4 a_16974_n1881.t1 dvss.t167 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X17 x7.ena_done_b.t0 a_21775_n2247.t2 dvdd.t53 dvdd.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X18 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X19 a_20121_n2241.t0 a_19955_n2241.t3 dvdd.t162 dvdd.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_2130_n21176.t1 a_24530_n21342.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X21 ibias_ip.t0 standby_33.t3 ibias.t1 ibias.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X22 xout.t18 vbreg.t9 avdd_ip.t28 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X23 inv_m1.t0 inv_in.t1 dvdd_ip.t1 dvdd_ip.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X24 a_2132_n15590.t1 a_18932_n15756.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X25 dout_ip.t1 inv_m2.t2 dvdd_ip.t10 dvdd_ip.t9 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X26 a_20733_n2791.t1 a_20689_n2549.t4 a_20567_n2791.t1 dvss.t39 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X27 inv_in.t2 xin_buf.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X28 x7.x1.x2.CLK.t1 a_15000_n1881.t3 dvss.t23 dvss.t22 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X29 avdd_ip.t29 avss_ip sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X30 a_16317_n1881.t1 a_16273_n2273.t4 a_16151_n1869.t1 dvss.t150 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X31 x7.stby_done_b.t0 a_21775_n2791.t2 dvss.t147 dvss.t146 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X32 a_14009_n2701.t1 x7.clk_disable.t2 dvss.t153 dvss.t131 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.07665 ps=0.785 w=0.42 l=0.15
X33 dvss.t34 standby_ip.t2 standby_b.t1 dvss.t33 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X34 dvss.t171 a_2971_n1521.t2 ena_ip.t1 dvss.t170 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X35 dvss.t202 standby_b.t3 a_16317_n2791.t1 dvss.t201 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X36 avdd_ip.t30 avss_ip sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X37 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X38 dvss.t151 x7.ena_done_b.t2 a_14035_n1997.t0 dvss.t8 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X39 x7.stby_done_b.t1 a_21775_n2791.t3 dvdd.t161 dvdd.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X40 a_2132_n17582.t1 a_18932_n17416.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X41 inv_m1.t1 inv_in.t3 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X42 avss.t26 avdd.t16 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X43 a_10620_n9666.t0 a_24220_n9832.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X44 a_20733_n1881.t1 a_20689_n2273.t4 a_20567_n1869.t1 dvss.t83 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X45 dvdd.t30 x7.x2.x2.CLK.t2 a_15539_n2791.t0 dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X46 a_16782_n2425.t1 a_15705_n2791.t2 a_16620_n2791.t3 dvdd.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X47 dvdd_ip.t8 inv_m1.t2 inv_m2.t0 dvdd_ip.t7 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X48 a_4857_n1521.t0 standby.t0 dvdd.t115 dvdd.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X49 avdd_ip.t3 x3.out_b.t3 avdd.t10 avdd.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X50 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X51 a_20121_n2791.t1 a_19955_n2791.t2 dvss.t149 dvss.t148 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X52 dvss.t27 ena_ip.t3 a_16317_n1881.t0 dvss.t26 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X53 x7.x1.Qb2.t0 a_19567_n2247.t2 dvss.t77 dvss.t76 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X54 dvss.t72 ena.t0 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X55 dvdd.t136 a_19003_n2817.t3 a_19567_n2791.t0 dvdd.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X56 avss_ip vg1.t0 vg1.t1 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X57 a_21145_n1869.t1 a_19955_n2241.t4 a_21036_n1869.t2 dvss.t40 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X58 avdd_ip.t21 vbreg.t10 avdd_ip.t20 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X59 a_21211_n2817.t0 standby_b.t4 dvdd.t103 dvdd.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X60 avss_ip xin.t6 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=23.6118 ps=175.6 w=4 l=0.5
X61 a_19003_n2817.t1 a_18828_n2791.t4 a_19182_n2791.t1 dvss.t174 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X62 a_15000_n1881.t2 dout_ip.t4 dvdd.t144 dvdd.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
X63 a_2132_n17250.t0 a_18932_n17416.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X64 a_20121_n2241.t1 a_19955_n2241.t5 dvss.t42 dvss.t41 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X65 dvss_ip ibias_ip.t11 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=5.8 ps=45.8 w=2 l=2
X66 a_10620_n9666.t1 a_24220_n9500.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X67 a_18359_n1869.t1 a_17913_n2241.t2 a_18263_n1869.t0 dvss.t24 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X68 xout.t17 vbreg.t11 avdd_ip.t27 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X69 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=75
X70 vbreg.t4 vg2.t5 vrb.t3 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X71 a_18525_n2791.t1 a_18481_n2549.t4 a_18359_n2791.t0 dvss.t180 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X72 a_2130_n20844.t1 a_24530_n21010.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X73 a_15083_n2791.t0 dout_ip.t5 a_15000_n2791.t2 dvss.t172 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X74 a_21036_n1869.t0 a_20121_n2241.t2 a_20689_n2273.t1 dvss.t175 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X75 dvss_ip standby_b.t5 dvss.t134 dvss.t133 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X76 a_2132_n15590.t0 a_18932_n15424.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X77 a_14285_n2079.t0 x7.ena_done_b.t3 a_14285_n2281.t0 dvdd.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X78 a_19003_n1943.t0 a_18828_n1869.t4 a_19182_n1881.t0 dvss.t75 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X79 vn.t6 xin.t7 vn.t5 dvdd_ip.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X80 avss.t19 standby_b.t6 standby_33.t1 avss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X81 a_10620_n7674.t0 a_24220_n7840.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X82 ibias_ip.t10 ibias_ip.t9 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X83 avdd.t18 x3.out_b.t4 avdd_ip.t6 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X84 a_15960_n2791.t2 x7.x2.Qb1.t2 dvdd.t95 dvdd.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X85 a_2130_n19516.t0 a_24530_n19682.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X86 xin.t8 avdd_ip.t2 sky130_fd_pr__diode_pd2nw_05v5 perim=1.8e+06 area=2.025e+11
X87 a_20579_n2247.t0 ena_ip.t4 dvdd.t62 dvdd.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X88 dvdd.t109 a_2971_n1521.t3 ena_ip.t0 dvdd.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X89 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X90 a_15083_n1881.t1 dout_ip.t6 a_15000_n1881.t1 dvss.t192 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X91 a_18525_n1881.t0 a_18481_n2273.t4 a_18359_n1869.t0 dvss.t18 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X92 a_18168_n2791.t1 x7.x2.Qb2.t2 dvdd.t23 dvdd.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X93 dvss.t118 standby_b.t7 a_18525_n2791.t0 dvss.t117 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X94 xin_buf.t2 xout.t23 tail.t0 dvdd_ip.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X95 a_16273_n2549.t0 a_16055_n2791.t4 dvdd.t9 dvdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X96 dvss.t191 x7.stby_done_b.t3 a_15083_n2791.t1 dvss.t190 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X97 xout.t4 xin.t9 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X98 x7.x1.x4.Q.t1 a_21211_n1943.t3 dvss.t164 dvss.t163 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X99 dvdd.t139 x7.stby_done_b.t4 a_15000_n2791.t1 dvdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X100 a_14009_n2404.t1 standby_ip.t3 a_14285_n2079.t2 dvdd.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X101 dvss_ip standby_b.t8 dvss.t36 dvss.t35 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X102 avdd_ip.t26 vbreg.t12 xout.t16 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X103 tail.t10 vbp.t4 dvdd_ip.t51 dvdd_ip.t32 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X104 a_2130_n20844.t0 a_24530_n20678.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X105 a_16729_n1869.t1 a_15539_n2241.t2 a_16620_n1869.t0 dvss.t119 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X106 avss_ip vg2.t4 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X107 dvdd_ip.t50 vbp.t5 dvdd_ip.t49 dvdd_ip.t29 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X108 a_16273_n2273.t0 a_16055_n1869.t4 dvdd.t51 dvdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X109 a_2132_n15258.t0 a_18932_n15424.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X110 a_18990_n2425.t1 a_17913_n2791.t3 a_18828_n2791.t3 dvdd.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X111 a_14285_n2281.t3 x7.stby_done_b.t5 dvdd.t138 dvdd.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X112 avdd_ip.t25 vbreg.t13 avdd_ip.t24 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X113 dvss.t53 ena_ip.t5 a_18525_n1881.t1 dvss.t52 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X114 dvdd.t131 a_21211_n1943.t4 a_21775_n2247.t0 dvdd.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X115 dvss.t90 x7.ena_done_b.t4 a_15083_n1881.t0 dvss.t89 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X116 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X117 a_16795_n1943.t0 ena_ip.t6 dvdd.t105 dvdd.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X118 dvss.t173 standby.t1 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X119 dvss.t38 standby_b.t9 dvss_ip dvss.t37 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X120 a_2130_n19516.t1 a_24530_n19350.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X121 dvdd.t11 a_14009_n2404.t4 x7.clk_disable.t1 dvdd.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X122 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X123 dvdd_ip.t54 standby_ip.t4 dvdd.t170 dvdd.t169 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X124 a_16163_n2247.t1 ena_ip.t7 dvdd.t107 dvdd.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X125 a_2132_n16918.t0 a_18932_n17084.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X126 dvdd.t173 x7.x2.Qb2.t3 a_19955_n2791.t1 dvdd.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X127 a_19003_n1943.t2 ena_ip.t8 dvdd.t73 dvdd.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X128 inv_in.t4 xin_buf.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X129 a_10620_n9334.t0 a_24220_n9500.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X130 dvss.t66 a_21211_n2817.t3 a_21775_n2791.t0 dvss.t65 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X131 a_3134_n13324.t0 vrb.t4 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=75
X132 dvdd_ip.t55 standby_ip.t5 dvdd.t172 dvdd.t171 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X133 a_16974_n2791.t0 standby_b.t10 dvss.t94 dvss.t93 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X134 x7.x1.x2.Q.t1 a_16795_n1943.t3 dvss.t30 dvss.t29 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X135 a_2132_n17582.t0 a_18932_n17748.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X136 dvdd.t3 x7.x1.x2.CLK.t2 a_15539_n2241.t0 dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X137 dvdd_ip.t48 vbp.t6 tail.t9 dvdd_ip.t27 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X138 a_19182_n2791.t0 standby_b.t11 dvss.t96 dvss.t95 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X139 dvss.t197 a_19003_n2817.t4 a_18937_n2791.t1 dvss.t196 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X140 avss_ip avss_ip avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X141 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X142 dout_ip.t3 inv_m2.t3 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X143 a_15705_n2791.t0 a_15539_n2791.t2 dvdd.t132 dvdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X144 avdd.t19 x3.out_b.t5 x3.out.t0 avdd.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X145 dvdd.t118 a_16795_n2817.t3 a_16782_n2425.t0 dvdd.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X146 dvss.t85 a_21211_n1943.t5 a_21775_n2247.t1 dvss.t84 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X147 xout.t22 xin.t10 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X148 avss_ip avss_ip avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X149 a_16974_n1881.t0 ena_ip.t9 dvss.t64 dvss.t63 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X150 dvdd.t65 a_16795_n1943.t4 a_17359_n2247.t0 dvdd.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X151 xin.t5 a_24530_n22338.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X152 avss_ip x3.out.t3 avss.t3 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X153 dvss.t155 x7.clk_disable.t3 dout_filt.t0 dvss.t154 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X154 a_16055_n2791.t1 a_15539_n2791.t3 a_15960_n2791.t0 dvss.t120 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X155 dvdd.t71 standby_ip.t6 dvdd_ip.t6 dvdd.t70 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X156 standby_33.t0 x4.out_b.t3 avdd.t2 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X157 a_16055_n1869.t2 a_15705_n2241.t3 a_15960_n1881.t3 dvdd.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X158 dvdd_ip.t47 vbp.t7 tail.t8 dvdd_ip.t40 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X159 a_20471_n2791.t3 a_20121_n2791.t2 a_20376_n2791.t3 dvdd.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X160 avss_ip xout.t24 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
**devattr s=257843176,88584 d=257843176,88584
X161 tail.t7 vbp.t8 dvdd_ip.t46 dvdd_ip.t38 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X162 dvdd.t154 a_19003_n2817.t5 a_18990_n2425.t0 dvdd.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X163 a_10620_n9334.t1 a_24220_n9168.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X164 a_19182_n1881.t1 ena_ip.t10 dvss.t188 dvss.t187 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X165 avdd_ip.t23 vbreg.t14 xout.t15 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X166 avss_ip xin.t11 xout.t21 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X167 xin_buf.t1 xout.t25 xin_buf.t1 dvdd_ip.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0 ps=0 w=4 l=2
X168 a_3134_n13324.t1 avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=75
X169 a_21036_n2791.t1 a_19955_n2791.t3 a_20689_n2549.t2 dvdd.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X170 dvss.t145 a_19003_n1943.t3 a_18937_n1869.t1 dvss.t144 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X171 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X172 a_18937_n2791.t0 a_17747_n2791.t2 a_18828_n2791.t0 dvss.t4 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X173 dvss.t157 a_16795_n2817.t4 a_17359_n2791.t1 dvss.t156 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X174 a_16273_n2273.t3 a_16055_n1869.t5 dvss.t177 dvss.t176 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X175 dvdd.t141 a_16620_n1869.t5 a_16795_n1943.t2 dvdd.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X176 x7.x1.x2.Q.t0 a_16795_n1943.t5 dvdd.t67 dvdd.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X177 a_2130_n20512.t0 a_24530_n20678.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X178 avss_ip xin.t12 xout.t2 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X179 dvdd.t166 a_21036_n2791.t4 a_21211_n2817.t2 dvdd.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X180 x4.out_b.t2 standby_ip.t7 avss.t15 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X181 a_18481_n2549.t0 a_18263_n2791.t4 dvdd.t1 dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X182 dvss_ip inv_m1.t3 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=7.9025 ps=61.46 w=0.5 l=1
X183 ibias_ip.t8 ibias_ip.t7 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X184 dvss.t49 x7.x2.x2.CLK.t3 a_15539_n2791.t1 dvss.t48 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X185 xout.t7 xin.t13 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X186 a_2132_n14926.t1 a_18932_n15092.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X187 dvdd.t46 x7.clk_disable.t4 a_14357_n2743.t0 dvdd.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.005 as=0.0672 ps=0.85 w=0.64 l=0.15
X188 vn.t2 vn.t0 vn.t1 dvss_ip sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X189 a_20567_n2791.t0 a_20121_n2791.t3 a_20471_n2791.t2 dvss.t138 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X190 dvdd.t78 standby_ip.t8 dvdd_ip.t11 dvdd.t77 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X191 dvss_ip dout_filt.t3 dout.t1 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=1
X192 a_20471_n1869.t2 a_19955_n2241.t6 a_20376_n1881.t3 dvss.t198 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X193 a_18481_n2273.t2 a_18263_n1869.t4 dvdd.t116 dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X194 avss.t7 x3.out.t4 avss_ip avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X195 dvss.t212 a_16795_n1943.t6 a_17359_n2247.t1 dvss.t211 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X196 x7.x1.Qb1.t0 a_17359_n2247.t2 dvdd.t134 dvdd.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X197 dvdd_ip.t45 vbp.t9 tail.t6 dvdd_ip.t34 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X198 avss.t27 avdd.t15 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X199 x7.x2.x2.Q.t0 a_16795_n2817.t5 dvdd.t151 dvdd.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X200 a_14035_n2743.t0 dout_ip.t7 dout_filt.t1 dvss.t131 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X201 dvss.t3 x7.x1.x2.CLK.t3 a_15539_n2241.t1 dvss.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X202 dout_ip.t2 inv_m2.t4 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X203 xin_buf.t3 vn.t8 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X204 avdd_ip.t22 vbreg.t15 vg1.t3 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X205 a_2130_n19848.t0 a_24530_n19682.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X206 vrb.t2 vg2.t6 vbreg.t3 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X207 a_18828_n1869.t2 a_17913_n2241.t3 a_18481_n2273.t1 dvss.t79 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X208 x7.x2.Qb1.t0 a_17359_n2791.t2 dvss.t194 dvss.t193 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X209 a_2130_n20512.t1 a_24530_n20346.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X210 dvdd.t50 a_20689_n2273.t5 a_20579_n2247.t1 dvdd.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X211 x7.x1.x2.CLK.t0 a_15000_n1881.t4 dvdd.t34 dvdd.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X212 dvdd_ip.t12 standby_ip.t9 dvdd.t80 dvdd.t79 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X213 a_2132_n14926.t0 a_18932_n14760.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X214 x7.x2.Qb1.t1 a_17359_n2791.t3 dvdd.t165 dvdd.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X215 x7.x1.x3.Q.t1 a_19003_n1943.t4 dvss.t124 dvss.t123 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X216 xout.t6 xin.t14 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X217 avdd.t12 x3.out_b.t6 avdd_ip.t4 avdd.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X218 a_16273_n2549.t2 a_16055_n2791.t5 dvss.t74 dvss.t73 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X219 a_16151_n2791.t1 a_15705_n2791.t3 a_16055_n2791.t3 dvss.t78 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X220 vg1.t4 xin.t4 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X221 avss_ip xin.t15 xout.t5 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X222 dvss_ip inv_m1.t4 inv_m2.t1 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X223 a_2130_n19184.t0 a_24530_n19018.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X224 dvdd_ip.t44 vbp.t10 dvdd_ip.t43 dvdd_ip.t42 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X225 inv_in.t5 xin_buf.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X226 dvdd.t128 a_4857_n1521.t2 standby_ip.t0 dvdd.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X227 a_14035_n1997.t1 ena_ip.t11 a_14009_n2404.t0 dvss.t8 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X228 a_17913_n2791.t0 a_17747_n2791.t3 dvdd.t5 dvdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X229 a_4857_n1521.t1 standby.t2 dvss.t137 dvss.t136 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X230 a_10620_n9002.t1 a_24220_n9168.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X231 a_18263_n2791.t0 a_17747_n2791.t4 a_18168_n2791.t0 dvss.t5 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X232 a_14009_n2404.t3 standby_b.t12 a_14035_n2281.t0 dvss.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X233 a_16620_n1869.t3 a_15539_n2241.t3 a_16273_n2273.t2 dvdd.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X234 a_18263_n1869.t1 a_17913_n2241.t4 a_18168_n1881.t2 dvdd.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X235 a_10620_n9002.t0 a_24220_n8836.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X236 dvdd.t94 x7.x1.Qb2.t3 a_19955_n2241.t0 dvdd.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X237 a_2130_n20180.t0 a_24530_n20346.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X238 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X239 x3.out_b.t0 x3.out.t5 avdd.t8 avdd.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X240 xout.t8 xin.t16 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X241 avdd.t1 standby_33.t4 x4.out_b.t0 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X242 a_20579_n2247.t2 a_19955_n2241.t7 a_20471_n1869.t3 dvdd.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X243 dvdd.t119 a_16273_n2273.t5 a_16163_n2247.t2 dvdd.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X244 a_15000_n2791.t0 dout_ip.t8 dvdd.t75 dvdd.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
X245 dvdd.t112 a_18828_n1869.t5 a_19003_n1943.t1 dvdd.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X246 a_2130_n22172.t1 a_24530_n22006.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X247 avss_ip xin.t17 xout.t3 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X248 avdd_ip.t31 avss_ip sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X249 a_15705_n2241.t0 a_15539_n2241.t4 dvdd.t13 dvdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X250 a_2130_n21840.t0 a_24530_n22006.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X251 avdd_ip.t19 vbreg.t16 xout.t14 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X252 dvdd.t60 x7.x2.Qb1.t3 a_17747_n2791.t0 dvdd.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X253 a_2132_n16586.t1 a_18932_n16420.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X254 avss_ip xin.t18 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X255 a_10620_n8670.t0 a_24220_n8836.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X256 xin_buf.t4 vn.t9 xin_buf.t4 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0 ps=0 w=4 l=2
X257 x7.x1.Qb2.t1 a_19567_n2247.t3 dvdd.t164 dvdd.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X258 a_2132_n17250.t1 a_18932_n17084.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X259 a_14009_n2701.t0 x7.clk_disable.t5 dvdd.t48 dvdd.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.10855 ps=1.005 w=0.42 l=0.15
X260 dvss.t17 x7.x2.Qb2.t4 a_19955_n2791.t0 dvss.t16 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X261 dvss.t32 standby_ip.t10 x7.clkin dvss.t31 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X262 dvss_ip ibias_ip.t12 vbp.t0 dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X263 inv_in.t6 xin_buf.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X264 a_22601_n15524.t1 vbreg.t17 a_22601_n15524.t0 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X265 a_20579_n2425.t1 standby_b.t13 dvdd.t104 dvdd.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X266 a_16163_n2247.t0 a_15539_n2241.t5 a_16055_n1869.t1 dvdd.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X267 avss_ip xin.t19 xout.t1 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X268 x7.x2.Qb2.t1 a_19567_n2791.t2 dvss.t82 dvss.t81 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X269 vbreg.t6 vg1.t5 vbreg.t5 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X270 vg1.t6 xin.t3 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X271 avss_ip x3.out.t6 avss.t1 avss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X272 x3.in_b.t1 ena_ip.t12 dvss.t98 dvss.t97 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X273 x7.x2.Qb2.t0 a_19567_n2791.t3 dvdd.t130 dvdd.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X274 dvss.t143 x7.x1.Qb2.t4 a_19955_n2241.t1 dvss.t142 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X275 a_15705_n2791.t1 a_15539_n2791.t4 dvss.t71 dvss.t70 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X276 standby_33.t2 standby_b.t14 avss.t17 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X277 vbreg.t0 vg2.t7 vrb.t1 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X278 tail.t1 xin.t20 vn.t7 dvdd_ip.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X279 dout_ip.t0 inv_m2.t5 dvdd_ip.t15 dvdd_ip.t9 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X280 dvdd.t175 dvss.t61 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X281 dvdd.t85 a_21211_n1943.t6 a_21198_n2247.t1 dvdd.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X282 a_2130_n20180.t1 a_24530_n20014.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X283 dvdd_ip.t37 vbp.t11 dvdd_ip.t36 dvdd_ip.t24 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X284 a_20376_n2791.t2 x7.stby_done_b.t6 dvss.t140 dvss.t139 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X285 a_18828_n1869.t1 a_17747_n2241.t2 a_18481_n2273.t0 dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X286 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X287 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X288 a_16795_n2817.t0 standby_b.t15 dvdd.t91 dvdd.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X289 a_2132_n14594.t1 a_18932_n14428.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X290 a_15705_n2241.t1 a_15539_n2241.t6 dvss.t126 dvss.t125 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X291 x3.out.t2 x3.in_b.t2 avss.t23 avss.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X292 a_16163_n2425.t2 standby_b.t16 dvdd.t122 dvdd.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X293 inv_in.t7 xin_buf.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X294 a_2132_n15258.t1 a_18932_n15092.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X295 a_19003_n2817.t0 standby_b.t17 dvdd.t123 dvdd.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X296 dvdd.t174 a_18481_n2273.t5 a_18371_n2247.t1 dvdd.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X297 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X298 a_20376_n1881.t1 x7.ena_done_b.t5 dvss.t92 dvss.t91 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X299 dvdd_ip.t14 inv_m1.t5 dvdd_ip.t13 dvdd_ip.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=1
X300 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X301 dvss.t106 standby_b.t18 dvss_ip dvss.t105 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X302 vg1.t7 xin.t2 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X303 a_2130_n19184.t1 a_24530_n19350.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X304 a_10620_n8670.t1 a_24220_n8504.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X305 a_17913_n2241.t0 a_17747_n2241.t3 dvdd.t35 dvdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X306 x7.x2.x4.Q.t1 a_21211_n2817.t4 dvss.t160 dvss.t159 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X307 dvss_ip ibias_ip.t5 ibias_ip.t6 dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X308 a_21198_n2247.t0 a_20121_n2241.t3 a_21036_n1869.t1 dvdd.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X309 a_20689_n2273.t3 a_20471_n1869.t4 dvss.t205 dvss.t204 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X310 x7.x1.x4.Q.t0 a_21211_n1943.t7 dvdd.t89 dvdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X311 xout.t20 vbreg.t18 xout.t19 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X312 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X313 a_2132_n16918.t1 a_18932_n16752.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X314 avss_ip vg2.t3 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X315 a_16055_n2791.t2 a_15705_n2791.t4 a_15960_n2791.t1 dvdd.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X316 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=75
X317 avss.t21 x3.in_b.t3 x3.out.t1 avss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X318 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X319 dvss_ip standby_b.t19 dvss.t108 dvss.t107 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X320 a_18371_n2247.t2 ena_ip.t13 dvdd.t88 dvdd.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X321 a_2130_n21508.t1 a_24530_n21674.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X322 a_18371_n2247.t0 a_17747_n2241.t4 a_18263_n1869.t2 dvdd.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X323 vbreg.t8 vbreg.t7 avdd_ip.t18 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X324 a_16620_n2791.t0 a_15705_n2791.t5 a_16273_n2549.t1 dvss.t43 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X325 x7.x2.x4.Q.t0 a_21211_n2817.t5 dvdd.t59 dvdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X326 dvdd.t126 a_16620_n2791.t5 a_16795_n2817.t2 dvdd.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X327 dvss_ip standby_b.t20 dvss.t208 dvss.t207 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X328 a_2130_n22172.t0 a_24530_n22338.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X329 a_10620_n8338.t1 a_24220_n8504.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X330 dvdd.t21 x7.x1.Qb1.t2 a_17747_n2241.t0 dvdd.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X331 dvdd.t43 standby_ip.t11 dvdd_ip.t3 dvdd.t42 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X332 inv_in.t8 xin_buf.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X333 a_2132_n16586.t0 a_18932_n16752.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X334 a_17913_n2791.t1 a_17747_n2791.t5 dvss.t7 dvss.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X335 a_16055_n1869.t0 a_15539_n2241.t7 a_15960_n1881.t2 dvss.t189 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X336 x7.x2.x2.Q.t1 a_16795_n2817.t6 dvss.t179 dvss.t178 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X337 avdd_ip.t32 avss_ip sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X338 x7.ena_done_b.t1 a_21775_n2247.t3 dvss.t130 dvss.t129 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X339 avss_ip vg2.t2 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X340 avss_ip avss_ip avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X341 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X342 a_20689_n2549.t1 a_20471_n2791.t4 dvss.t20 dvss.t19 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X343 dvss.t210 standby_b.t21 dvss_ip dvss.t209 sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X344 dvdd.t163 a_19003_n1943.t5 a_19567_n2247.t1 dvdd.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X345 dvdd_ip.t17 a_9120_n9346.t1 a_9120_n9346.t2 dvdd_ip.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X346 dvdd.t101 a_21211_n2817.t6 a_21775_n2791.t1 dvdd.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X347 a_20376_n1881.t0 x7.ena_done_b.t6 dvdd.t25 dvdd.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X348 a_18937_n1869.t0 a_17747_n2241.t5 a_18828_n1869.t0 dvss.t80 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X349 avss_ip xin.t21 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
**devattr s=257843176,88584 d=257843176,88584
X350 dvdd_ip.t41 vbp.t12 tail.t5 dvdd_ip.t40 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X351 a_21211_n2817.t1 a_21036_n2791.t5 a_21390_n2791.t1 dvss.t203 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X352 tail.t4 vbp.t13 dvdd_ip.t39 dvdd_ip.t38 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X353 a_17913_n2241.t1 a_17747_n2241.t6 dvss.t69 dvss.t68 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X354 dvdd.t54 a_20689_n2549.t5 a_20579_n2425.t2 dvdd.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X355 dvdd_ip.t53 standby_ip.t12 dvdd.t168 dvdd.t167 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X356 a_20567_n1869.t0 a_20121_n2241.t4 a_20471_n1869.t0 dvss.t183 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X357 dvdd.t176 dvss.t62 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X358 dvss.t162 a_19003_n2817.t6 a_19567_n2791.t1 dvss.t161 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X359 a_18481_n2273.t3 a_18263_n1869.t5 dvss.t45 dvss.t44 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X360 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X361 dvss_ip vn.t3 vn.t4 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X362 a_2130_n18852.t1 a_24530_n19018.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X363 dvss.t59 x7.x2.Qb1.t4 a_17747_n2791.t1 dvss.t58 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X364 dvdd.t177 dvss.t87 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X365 avss.t28 avdd.t14 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X366 avss.t13 standby_ip.t13 x4.out_b.t1 avss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X367 icnode.t0 vg2.t8 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X368 avdd_ip.t17 vbreg.t19 xout.t13 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X369 a_21211_n1943.t1 a_21036_n1869.t5 a_21390_n1881.t1 dvss.t86 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X370 a_15960_n2791.t3 x7.x2.Qb1.t5 dvss.t116 dvss.t115 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X371 a_11526_n12394.t0 icnode.t1 a_8268_n12482.t1 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X372 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X373 dvss.t51 a_19003_n1943.t6 a_19567_n2247.t0 dvss.t50 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X374 xout.t12 vbreg.t20 avdd_ip.t16 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X375 dvss.t195 a_4857_n1521.t3 standby_ip.t1 dvss.t136 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X376 a_14009_n2404.t2 standby_ip.t14 dvss.t60 dvss.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X377 inv_in.t9 xin_buf.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X378 dvdd_ip.t35 vbp.t1 vbp.t2 dvdd_ip.t34 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X379 a_2132_n14594.t0 a_18932_n14760.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X380 a_16620_n2791.t1 a_15539_n2791.t5 a_16273_n2549.t3 dvdd.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X381 dvss.t13 x7.x1.Qb1.t3 a_17747_n2241.t1 dvss.t12 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X382 a_18263_n2791.t3 a_17913_n2791.t4 a_18168_n2791.t3 dvdd.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X383 dvdd.t156 a_16795_n2817.t7 a_17359_n2791.t0 dvdd.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X384 a_2971_n1521.t0 ena.t1 dvss.t110 dvss.t109 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X385 dvss.t100 standby_b.t22 a_20733_n2791.t0 dvss.t99 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X386 a_15960_n1881.t1 x7.x1.Qb1.t4 dvss.t11 dvss.t10 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X387 a_14035_n2281.t1 x7.stby_done_b.t7 dvss.t141 dvss.t8 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X388 a_20579_n2425.t0 a_19955_n2791.t4 a_20471_n2791.t1 dvdd.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X389 a_21145_n2791.t0 a_19955_n2791.t5 a_21036_n2791.t0 dvss.t25 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X390 dvdd.t32 a_16273_n2549.t5 a_16163_n2425.t0 dvdd.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X391 a_16151_n1869.t0 a_15705_n2241.t4 a_16055_n1869.t3 dvss.t121 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X392 a_2130_n18852.t0 xout.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X393 dvdd.t147 a_18828_n2791.t5 a_19003_n2817.t2 dvdd.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X394 a_16782_n2247.t1 a_15705_n2241.t5 a_16620_n1869.t2 dvdd.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X395 x3.out_b.t2 ena_ip.t14 avss.t11 avss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X396 dvss.t9 a_14009_n2404.t5 x7.clk_disable.t0 dvss.t8 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X397 avss.t29 avdd.t13 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X398 dvdd.t69 standby_ip.t15 dvdd_ip.t5 dvdd.t68 sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X399 a_18481_n2549.t1 a_18263_n2791.t5 dvss.t1 dvss.t0 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X400 a_18359_n2791.t1 a_17913_n2791.t5 a_18263_n2791.t2 dvss.t184 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X401 avdd_ip.t0 x3.out_b.t7 avdd.t4 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X402 a_18263_n1869.t3 a_17747_n2241.t7 a_18168_n1881.t3 dvss.t206 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X403 dvss.t47 ena_ip.t15 a_20733_n1881.t0 dvss.t46 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X404 x7.x2.x3.Q.t1 a_19003_n2817.t7 dvss.t169 dvss.t168 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X405 xout.t11 vbreg.t21 avdd_ip.t15 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X406 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X407 x7.x1.x3.Q.t0 a_19003_n1943.t7 dvdd.t146 dvdd.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X408 a_21036_n2791.t2 a_20121_n2791.t4 a_20689_n2549.t3 dvss.t67 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X409 dvss.t102 standby_b.t23 dvss_ip dvss.t101 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X410 avdd_ip.t33 icnode.t1 sky130_fd_pr__cap_mim_m3_1 l=20 w=20
X411 a_21211_n1943.t0 ena_ip.t16 dvdd.t157 dvdd.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X412 inv_in.t10 xin_buf.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X413 inv_in.t11 xin_buf.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X414 a_10620_n8006.t1 a_24220_n8172.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X415 avdd_ip.t14 vbreg.t22 xout.t10 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X416 a_2130_n21840.t1 a_24530_n21674.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X417 inv_in.t12 xin_buf.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X418 a_10620_n8006.t0 a_24220_n7840.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X419 avdd.t6 x3.out_b.t8 avdd_ip.t1 avdd.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X420 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X421 avss.t9 ena_ip.t17 x3.out_b.t1 avss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X422 a_2132_n16254.t0 a_18932_n16420.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X423 a_16163_n2425.t1 a_15539_n2791.t6 a_16055_n2791.t0 dvdd.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X424 tail.t3 vbp.t14 dvdd_ip.t33 dvdd_ip.t32 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X425 a_8268_n12482.t1 a_8268_n12482.t0 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X426 x7.x2.x3.Q.t0 a_19003_n2817.t8 dvdd.t150 dvdd.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X427 dvss.t132 a_14009_n2701.t2 a_14035_n2743.t1 dvss.t131 sky130_fd_pr__nfet_01v8 ad=0.07665 pd=0.785 as=0.0441 ps=0.63 w=0.42 l=0.15
X428 x7.x2.x2.CLK.t0 a_15000_n2791.t4 dvdd.t160 dvdd.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X429 dvdd_ip.t31 vbp.t15 dvdd_ip.t30 dvdd_ip.t29 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X430 a_21390_n2791.t0 standby_b.t24 dvss.t55 dvss.t54 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X431 dvss.t128 a_21211_n2817.t7 a_21145_n2791.t1 dvss.t127 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X432 vg1.t8 xin.t1 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X433 dvss_ip standby_b.t25 dvss.t57 dvss.t56 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X434 inv_in.t13 xin_buf.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X435 a_16729_n2791.t1 a_15539_n2791.t7 a_16620_n2791.t2 dvss.t158 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X436 a_9120_n9346.t4 a_9120_n9346.t3 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X437 a_2130_n21176.t0 a_24530_n21010.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X438 a_2132_n17914.t1 vg1.t2 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X439 a_15960_n1881.t0 x7.x1.Qb1.t5 dvdd.t19 dvdd.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X440 a_20121_n2791.t0 a_19955_n2791.t6 dvdd.t82 dvdd.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X441 dvdd.t143 a_21211_n2817.t8 a_21198_n2425.t0 dvdd.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X442 a_14357_n2743.t1 dout_ip.t9 dout_filt.t2 dvdd.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X443 a_2971_n1521.t1 ena.t2 dvdd.t149 dvdd.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X444 a_21390_n1881.t0 ena_ip.t18 dvss.t112 dvss.t111 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X445 standby_b.t0 standby_ip.t16 dvdd.t39 dvdd.t38 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X446 dvss_ip ibias_ip.t3 ibias_ip.t4 dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X447 avss_ip x3.out.t7 avss.t5 avss.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X448 a_18828_n2791.t1 a_17747_n2791.t6 a_18481_n2549.t2 dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X449 a_18168_n1881.t0 x7.x1.Qb2.t5 dvdd.t113 dvdd.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X450 dvdd.t178 dvss.t88 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X451 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X452 dvss.t104 a_21211_n1943.t8 a_21145_n1869.t0 dvss.t103 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X453 a_14285_n2281.t1 ena_ip.t19 a_14285_n2079.t1 dvdd.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X454 avdd_ip.t13 vbreg.t23 avdd_ip.t12 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X455 a_2132_n16254.t1 a_18932_n16088.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X456 a_20689_n2549.t0 a_20471_n2791.t5 dvdd.t29 dvdd.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X457 dvdd.t27 x7.ena_done_b.t7 a_15000_n1881.t0 dvdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X458 dvdd.t15 standby_b.t26 a_14285_n2281.t2 dvdd.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X459 dvdd.t153 a_18481_n2549.t5 a_18371_n2425.t2 dvdd.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X460 dvdd_ip.t28 vbp.t16 tail.t2 dvdd_ip.t27 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X461 xout.t9 vbreg.t24 avdd_ip.t10 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X462 a_18990_n2247.t1 a_17913_n2241.t5 a_18828_n1869.t3 dvdd.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X463 a_20689_n2273.t0 a_20471_n1869.t5 dvdd.t99 dvdd.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X464 dvss_ip ibias_ip.t13 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X465 vg1.t9 xin.t0 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X466 avss.t25 x3.out.t8 avss_ip avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X467 avss_ip avss_ip avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X468 a_2132_n17914.t0 a_18932_n17748.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X469 a_2132_n14262.t0 a_18932_n14428.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X470 a_21198_n2425.t1 a_20121_n2791.t5 a_21036_n2791.t3 dvdd.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X471 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X472 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X473 dvss.t182 a_16795_n2817.t8 a_16729_n2791.t0 dvss.t181 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X474 inv_in.t14 xin_buf.t0 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X475 dvdd_ip.t26 vbp.t17 dvdd_ip.t25 dvdd_ip.t24 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X476 dvdd_ip.t2 standby_ip.t17 dvdd.t41 dvdd.t40 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X477 avss_ip vg2.t1 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X478 a_2132_n15922.t1 a_18932_n16088.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X479 a_18371_n2425.t1 standby_b.t27 dvdd.t17 dvdd.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X480 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X481 a_18371_n2425.t0 a_17747_n2791.t7 a_18263_n2791.t1 dvdd.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X482 ibias_ip.t2 ibias_ip.t1 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X483 dvss.t214 a_16795_n1943.t7 a_16729_n1869.t0 dvss.t213 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X484 dout.t0 dout_filt.t4 dvdd_ip.t21 dvdd_ip.t20 sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X485 a_2132_n14262.t1 vg2.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X486 dvdd.t155 a_16795_n1943.t8 a_16782_n2247.t0 dvdd.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X487 avdd_ip.t9 vbreg.t25 avdd_ip.t8 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X488 xout.t26 avdd_ip.t5 sky130_fd_pr__diode_pd2nw_05v5 perim=1.8e+06 area=2.025e+11
X489 a_20471_n2791.t0 a_19955_n2791.t7 a_20376_n2791.t0 dvss.t28 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X490 x7.x1.Qb1.t1 a_17359_n2247.t3 dvss.t166 dvss.t165 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X491 a_20471_n1869.t1 a_20121_n2241.t5 a_20376_n1881.t2 dvdd.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X492 dvdd.t56 standby_ip.t18 dvdd_ip.t4 dvdd.t55 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X493 a_2130_n21508.t0 a_24530_n21342.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X494 a_10620_n7674.t1 inv_in.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X495 dvdd.t121 a_19003_n1943.t8 a_18990_n2247.t0 dvdd.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X496 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X497 a_18168_n2791.t2 x7.x2.Qb2.t5 dvss.t15 dvss.t14 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X498 vrb.t0 vg2.t9 vbreg.t1 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X499 a_2132_n15922.t0 a_18932_n15756.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
R0 a_15705_n2241.t0 a_15705_n2241.n3 370.026
R1 a_15705_n2241.n0 a_15705_n2241.t2 351.356
R2 a_15705_n2241.n1 a_15705_n2241.t4 334.717
R3 a_15705_n2241.n3 a_15705_n2241.t1 325.971
R4 a_15705_n2241.n1 a_15705_n2241.t3 309.935
R5 a_15705_n2241.n0 a_15705_n2241.t5 305.683
R6 a_15705_n2241.n2 a_15705_n2241.n0 16.879
R7 a_15705_n2241.n3 a_15705_n2241.n2 10.8867
R8 a_15705_n2241.n2 a_15705_n2241.n1 9.3005
R9 a_16273_n2273.n3 a_16273_n2273.n2 647.119
R10 a_16273_n2273.n1 a_16273_n2273.t4 350.253
R11 a_16273_n2273.n2 a_16273_n2273.n0 260.339
R12 a_16273_n2273.n2 a_16273_n2273.n1 246.119
R13 a_16273_n2273.n1 a_16273_n2273.t5 189.588
R14 a_16273_n2273.n3 a_16273_n2273.t2 89.1195
R15 a_16273_n2273.n0 a_16273_n2273.t1 63.3338
R16 a_16273_n2273.t0 a_16273_n2273.n3 41.0422
R17 a_16273_n2273.n0 a_16273_n2273.t3 31.9797
R18 a_16620_n1869.n3 a_16620_n1869.n2 636.953
R19 a_16620_n1869.n1 a_16620_n1869.t4 366.856
R20 a_16620_n1869.n2 a_16620_n1869.n0 300.2
R21 a_16620_n1869.n2 a_16620_n1869.n1 225.036
R22 a_16620_n1869.n1 a_16620_n1869.t5 174.056
R23 a_16620_n1869.n0 a_16620_n1869.t1 70.0005
R24 a_16620_n1869.n3 a_16620_n1869.t3 68.0124
R25 a_16620_n1869.t2 a_16620_n1869.n3 63.3219
R26 a_16620_n1869.n0 a_16620_n1869.t0 61.6672
R27 dvss.n525 dvss.n524 184282
R28 dvss.n526 dvss.n525 126661
R29 dvss.n525 dvss.n124 10977.5
R30 dvss.n51 dvss.n17 8366.71
R31 dvss.n51 dvss.n18 8366.71
R32 dvss.n47 dvss.n18 8366.71
R33 dvss.n47 dvss.n17 8366.71
R34 dvss.n114 dvss.n113 7092.07
R35 dvss.n113 dvss.n112 5700.48
R36 dvss.n36 dvss.n31 4247.09
R37 dvss.n43 dvss.n31 4247.09
R38 dvss.n36 dvss.n32 4247.09
R39 dvss.n43 dvss.n32 4247.09
R40 dvss.n192 dvss.n186 4247.09
R41 dvss.n197 dvss.n186 4247.09
R42 dvss.n192 dvss.n187 4247.09
R43 dvss.n197 dvss.n187 4247.09
R44 dvss.n85 dvss.n15 2798.56
R45 dvss.n528 dvss.n15 2798.56
R46 dvss.n85 dvss.n16 2798.56
R47 dvss.n528 dvss.n16 2798.56
R48 dvss.n122 dvss.n54 2798.56
R49 dvss.n115 dvss.n54 2798.56
R50 dvss.n122 dvss.n55 2798.56
R51 dvss.n115 dvss.n55 2798.56
R52 dvss.n46 dvss.n44 2575.49
R53 dvss.n391 dvss.n390 2387.64
R54 dvss.n124 dvss.n123 2028.39
R55 dvss.n124 dvss.n52 2022.88
R56 dvss.n113 dvss.n86 1748.54
R57 dvss.n392 dvss.n391 1680.95
R58 dvss.n93 dvss.n88 1407.97
R59 dvss.n110 dvss.n88 1407.97
R60 dvss.n110 dvss.n89 1407.97
R61 dvss.n66 dvss.n63 1407.97
R62 dvss.n66 dvss.n64 1407.97
R63 dvss.n67 dvss.n63 1407.97
R64 dvss.n67 dvss.n64 1407.97
R65 dvss.n557 dvss.n0 1212.38
R66 dvss.n82 dvss.n81 1198.25
R67 dvss.n199 dvss.n7 1198.25
R68 dvss.n390 dvss.n389 1198.25
R69 dvss.n377 dvss.n206 1198.25
R70 dvss.n337 dvss.n223 1198.25
R71 dvss.n297 dvss.n240 1198.25
R72 dvss.n257 dvss.n125 1198.25
R73 dvss.n523 dvss.n522 1198.25
R74 dvss.n189 dvss.n144 1198.25
R75 dvss.n190 dvss.n161 1198.25
R76 dvss.n403 dvss.n180 1198.25
R77 dvss.n393 dvss.n392 1198.25
R78 dvss.n105 dvss.n87 1198.25
R79 dvss.n557 dvss.n556 1175.19
R80 dvss.t41 dvss.t91 935.78
R81 dvss.t113 dvss.t68 935.78
R82 dvss.t10 dvss.t125 935.78
R83 dvss.n50 dvss.n49 784.03
R84 dvss.n25 dvss.n24 783.962
R85 dvss.n49 dvss.n48 783.75
R86 dvss.n30 dvss.n25 783.683
R87 dvss.n206 dvss.t22 748.625
R88 dvss.t148 dvss.t139 717.851
R89 dvss.t6 dvss.t14 717.851
R90 dvss.t115 dvss.t70 717.851
R91 dvss.t163 dvss.t84 689.909
R92 dvss.t86 dvss.t163 689.909
R93 dvss.t50 dvss.t123 689.909
R94 dvss.t123 dvss.t75 689.909
R95 dvss.t211 dvss.t29 689.909
R96 dvss.t29 dvss.t167 689.909
R97 dvss.n527 dvss.n526 639.12
R98 dvss.n86 dvss.t97 618.75
R99 dvss.n527 dvss.t97 618.75
R100 dvss.t183 dvss.t83 609.174
R101 dvss.t18 dvss.t24 609.174
R102 dvss.t150 dvss.t121 609.174
R103 dvss.t185 dvss.n180 574.28
R104 dvss.t129 dvss.n125 554.129
R105 dvss.n240 dvss.t76 554.129
R106 dvss.n223 dvss.t165 554.129
R107 dvss.t103 dvss.t111 546.789
R108 dvss.t187 dvss.t144 546.789
R109 dvss.t63 dvss.t213 546.789
R110 dvss.t159 dvss.t65 529.24
R111 dvss.t203 dvss.t159 529.24
R112 dvss.t168 dvss.t161 529.24
R113 dvss.t174 dvss.t168 529.24
R114 dvss.t178 dvss.t156 529.24
R115 dvss.t152 dvss.t178 529.24
R116 dvss.t46 dvss.t204 484.404
R117 dvss.t44 dvss.t52 484.404
R118 dvss.t176 dvss.t26 484.404
R119 dvss.t138 dvss.t39 467.307
R120 dvss.t184 dvss.t180 467.307
R121 dvss.t78 dvss.t21 467.307
R122 dvss.t22 dvss.t89 447.707
R123 dvss.n391 dvss.n199 426.382
R124 dvss.n523 dvss.t146 425.08
R125 dvss.t81 dvss.n189 425.08
R126 dvss.t193 dvss.n190 425.08
R127 dvss.t127 dvss.t54 419.45
R128 dvss.t196 dvss.t95 419.45
R129 dvss.t181 dvss.t93 419.45
R130 dvss.n111 dvss.n87 419.18
R131 dvss.t175 dvss.t40 400
R132 dvss.t80 dvss.t79 400
R133 dvss.t119 dvss.t122 400
R134 dvss.n93 dvss.n92 390.825
R135 dvss.t99 dvss.t19 371.594
R136 dvss.t117 dvss.t0 371.594
R137 dvss.t201 dvss.t73 371.594
R138 dvss.n526 dvss.t170 366.435
R139 dvss.t204 dvss.t175 363.303
R140 dvss.t79 dvss.t44 363.303
R141 dvss.t122 dvss.t176 363.303
R142 dvss.t84 dvss.t129 355.964
R143 dvss.t76 dvss.t50 355.964
R144 dvss.t165 dvss.t211 355.964
R145 dvss.t40 dvss.t103 352.295
R146 dvss.t198 dvss.t183 352.295
R147 dvss.t144 dvss.t80 352.295
R148 dvss.t24 dvss.t206 352.295
R149 dvss.t213 dvss.t119 352.295
R150 dvss.t121 dvss.t189 352.295
R151 dvss.t91 dvss.t198 348.625
R152 dvss.t206 dvss.t113 348.625
R153 dvss.t189 dvss.t10 348.625
R154 dvss.n112 dvss.n111 344.228
R155 dvss.t190 dvss.t185 343.442
R156 dvss.t111 dvss.t86 333.945
R157 dvss.t75 dvss.t187 333.945
R158 dvss.t167 dvss.t63 333.945
R159 dvss.n524 dvss.n125 308.257
R160 dvss.t142 dvss.t41 308.257
R161 dvss.t68 dvss.t12 308.257
R162 dvss.t125 dvss.t2 308.257
R163 dvss.n87 dvss 308.139
R164 dvss.n371 dvss.t11 307.536
R165 dvss.n331 dvss.t114 307.536
R166 dvss.n291 dvss.t92 307.536
R167 dvss.n141 dvss.t140 307.536
R168 dvss.n158 dvss.t15 307.536
R169 dvss.n409 dvss.t116 307.536
R170 dvss.t67 dvss.t25 306.846
R171 dvss.t135 dvss.t4 306.846
R172 dvss.t43 dvss.t158 306.846
R173 dvss.n64 dvss.n62 292.5
R174 dvss.n64 dvss.n59 292.5
R175 dvss.n68 dvss.n67 292.5
R176 dvss.n67 dvss.t173 292.5
R177 dvss.n63 dvss.n61 292.5
R178 dvss.n63 dvss.n53 292.5
R179 dvss.n66 dvss.n65 292.5
R180 dvss.t173 dvss.n66 292.5
R181 dvss.n91 dvss.n89 292.5
R182 dvss.n110 dvss.n109 292.5
R183 dvss.n111 dvss.n110 292.5
R184 dvss.n90 dvss.n88 292.5
R185 dvss.n88 dvss.t72 292.5
R186 dvss.n94 dvss.n93 292.5
R187 dvss.t192 dvss 289.909
R188 dvss.t19 dvss.t67 278.695
R189 dvss.t0 dvss.t135 278.695
R190 dvss.t73 dvss.t43 278.695
R191 dvss.n196 dvss.n194 276.286
R192 dvss.n240 dvss 275.229
R193 dvss dvss.n223 275.229
R194 dvss dvss.n206 275.229
R195 dvss.n390 dvss 275.229
R196 dvss.t31 dvss.n0 273.678
R197 dvss.n44 dvss.t31 273.678
R198 dvss.t65 dvss.t146 273.065
R199 dvss.t161 dvss.t81 273.065
R200 dvss.t156 dvss.t193 273.065
R201 dvss.t25 dvss.t127 270.25
R202 dvss.t28 dvss.t138 270.25
R203 dvss.t4 dvss.t196 270.25
R204 dvss.t5 dvss.t184 270.25
R205 dvss.t158 dvss.t181 270.25
R206 dvss.t139 dvss.t28 267.435
R207 dvss.t14 dvss.t5 267.435
R208 dvss.t120 dvss.t115 267.435
R209 dvss.t83 dvss.t46 264.221
R210 dvss.t52 dvss.t18 264.221
R211 dvss.t26 dvss.t150 264.221
R212 dvss.t89 dvss.t192 264.221
R213 dvss.t54 dvss.t203 256.175
R214 dvss.t95 dvss.t174 256.175
R215 dvss.t93 dvss.t152 256.175
R216 dvss.n46 dvss.t209 255.168
R217 dvss.n52 dvss.t35 255.168
R218 dvss.n344 dvss.t30 246.817
R219 dvss.n304 dvss.t124 246.817
R220 dvss.n264 dvss.t164 246.817
R221 dvss.n131 dvss.t160 246.817
R222 dvss.n474 dvss.t169 246.817
R223 dvss.n435 dvss.t179 246.817
R224 dvss.t109 dvss.t170 244.291
R225 dvss dvss.t142 238.532
R226 dvss.t12 dvss 238.532
R227 dvss.t2 dvss 238.532
R228 dvss.n524 dvss.n523 236.469
R229 dvss.t16 dvss.t148 236.469
R230 dvss.t58 dvss.t6 236.469
R231 dvss.t70 dvss.t48 236.469
R232 dvss.n123 dvss.n53 230.855
R233 dvss.n413 dvss.t155 229.185
R234 dvss.n33 dvss.t32 219.8
R235 dvss.n42 dvss.n34 217.329
R236 dvss.n194 dvss.n193 217.225
R237 dvss.n220 dvss.n219 214.742
R238 dvss.n237 dvss.n236 214.742
R239 dvss.n254 dvss.n253 214.742
R240 dvss.n130 dvss.n129 214.742
R241 dvss.n480 dvss.n146 214.742
R242 dvss.n441 dvss.n163 214.742
R243 dvss.n189 dvss 211.132
R244 dvss.n190 dvss 211.132
R245 dvss dvss.n180 211.132
R246 dvss.n392 dvss 211.132
R247 dvss.n351 dvss.n216 209.254
R248 dvss.n311 dvss.n233 209.254
R249 dvss.n271 dvss.n250 209.254
R250 dvss.n134 dvss.n133 209.254
R251 dvss.n152 dvss.n151 209.254
R252 dvss.n169 dvss.n168 209.254
R253 dvss.t209 dvss.t107 208.894
R254 dvss.t107 dvss.t37 208.894
R255 dvss.t37 dvss.t56 208.894
R256 dvss.t56 dvss.t101 208.894
R257 dvss.t133 dvss.t199 208.894
R258 dvss.t199 dvss.t207 208.894
R259 dvss.t207 dvss.t105 208.894
R260 dvss.t105 dvss.t35 208.894
R261 dvss.t39 dvss.t99 202.688
R262 dvss.t180 dvss.t117 202.688
R263 dvss.t21 dvss.t201 202.688
R264 dvss.t172 dvss.t190 202.688
R265 dvss.n542 dvss.n6 202.067
R266 dvss.n3 dvss.n2 200.516
R267 dvss.n77 dvss.n76 199.739
R268 dvss.n208 dvss.n207 199.739
R269 dvss.n359 dvss.n358 199.739
R270 dvss.n225 dvss.n224 199.739
R271 dvss.n319 dvss.n318 199.739
R272 dvss.n242 dvss.n241 199.739
R273 dvss.n279 dvss.n278 199.739
R274 dvss.n500 dvss.n138 199.739
R275 dvss.n487 dvss.n143 199.739
R276 dvss.n461 dvss.n155 199.739
R277 dvss.n448 dvss.n160 199.739
R278 dvss.n422 dvss.n172 199.739
R279 dvss.n179 dvss.n178 199.739
R280 dvss.n102 dvss.n101 199.739
R281 dvss.n42 dvss.n41 198.024
R282 dvss.t33 dvss.n53 187.785
R283 dvss.n383 dvss.n382 185
R284 dvss.n185 dvss.n184 185
R285 dvss.n555 dvss.n554 185
R286 dvss dvss.t16 182.982
R287 dvss dvss.t58 182.982
R288 dvss.n84 dvss.n12 181.835
R289 dvss.n84 dvss.n83 181.835
R290 dvss.n116 dvss.n58 181.835
R291 dvss.n117 dvss.n116 181.835
R292 dvss.n92 dvss.n89 174.962
R293 dvss.n191 dvss.t120 166.091
R294 dvss.n198 dvss.t172 154.831
R295 dvss.n34 dvss.n31 148.029
R296 dvss.n197 dvss.n196 146.25
R297 dvss.n198 dvss.n197 146.25
R298 dvss.n193 dvss.n192 146.25
R299 dvss.n192 dvss.n191 146.25
R300 dvss.n35 dvss.n32 146.25
R301 dvss.n32 dvss.t31 146.25
R302 dvss.n31 dvss.t31 146.25
R303 dvss.n37 dvss.n34 143.809
R304 dvss dvss.t136 141.269
R305 dvss.t48 dvss.t154 140.756
R306 dvss dvss.t131 140.144
R307 dvss.n196 dvss.n195 127.487
R308 dvss.n114 dvss.n82 122.319
R309 dvss.n116 dvss.n115 117.001
R310 dvss.n115 dvss.n114 117.001
R311 dvss.n117 dvss.n55 117.001
R312 dvss.t33 dvss.n55 117.001
R313 dvss.n122 dvss.n121 117.001
R314 dvss.n123 dvss.n122 117.001
R315 dvss.n58 dvss.n54 117.001
R316 dvss.t33 dvss.n54 117.001
R317 dvss.n529 dvss.n528 117.001
R318 dvss.n528 dvss.n527 117.001
R319 dvss.n16 dvss.n12 117.001
R320 dvss.t97 dvss.n16 117.001
R321 dvss.n85 dvss.n84 117.001
R322 dvss.n86 dvss.n85 117.001
R323 dvss.n83 dvss.n15 117.001
R324 dvss.t97 dvss.n15 117.001
R325 dvss.t101 dvss.n45 104.448
R326 dvss.n45 dvss.t133 104.448
R327 dvss.n191 dvss.t78 104.159
R328 dvss.n529 dvss.n13 102.025
R329 dvss.n530 dvss.n529 102.025
R330 dvss.n121 dvss.n56 102.025
R331 dvss.n121 dvss.n120 102.025
R332 dvss.n216 dvss.t64 100.001
R333 dvss.n233 dvss.t188 100.001
R334 dvss.n250 dvss.t112 100.001
R335 dvss.n133 dvss.t55 100.001
R336 dvss.n151 dvss.t96 100.001
R337 dvss.n168 dvss.t94 100.001
R338 dvss.n65 dvss.n62 91.4829
R339 dvss.n94 dvss.n90 91.4829
R340 dvss.n71 dvss.t34 83.7183
R341 dvss.n96 dvss.t98 83.7183
R342 dvss.n92 dvss.t72 81.1932
R343 dvss dvss.t109 80.5052
R344 dvss.n530 dvss.n12 79.8123
R345 dvss.n83 dvss.n13 79.8123
R346 dvss.n58 dvss.n56 79.8123
R347 dvss.n120 dvss.n117 79.8123
R348 dvss.n382 dvss.t23 72.8576
R349 dvss.n358 dvss.t27 72.8576
R350 dvss.n318 dvss.t53 72.8576
R351 dvss.n278 dvss.t47 72.8576
R352 dvss.n184 dvss.t186 72.8576
R353 dvss.n138 dvss.t100 72.8576
R354 dvss.n155 dvss.t118 72.8576
R355 dvss.n172 dvss.t202 72.8576
R356 dvss.n216 dvss.t214 70.0005
R357 dvss.n233 dvss.t145 70.0005
R358 dvss.n250 dvss.t104 70.0005
R359 dvss.n133 dvss.t128 70.0005
R360 dvss.n151 dvss.t197 70.0005
R361 dvss.n168 dvss.t182 70.0005
R362 dvss.n68 dvss.n62 69.6045
R363 dvss.n109 dvss.n90 69.0306
R364 dvss.t173 dvss 68.912
R365 dvss.n188 dvss.n176 68.8106
R366 dvss dvss.n198 67.5629
R367 dvss.n65 dvss.n61 66.3131
R368 dvss.n95 dvss.n94 65.475
R369 dvss.n358 dvss.t177 60.5809
R370 dvss.n318 dvss.t45 60.5809
R371 dvss.n278 dvss.t205 60.5809
R372 dvss.n138 dvss.t20 60.5809
R373 dvss.n155 dvss.t1 60.5809
R374 dvss.n172 dvss.t74 60.5809
R375 dvss.n382 dvss.t90 58.5719
R376 dvss.n184 dvss.t191 58.5719
R377 dvss.n219 dvss.t212 57.1434
R378 dvss.n236 dvss.t51 57.1434
R379 dvss.n253 dvss.t85 57.1434
R380 dvss.n129 dvss.t66 57.1434
R381 dvss.n146 dvss.t162 57.1434
R382 dvss.n163 dvss.t157 57.1434
R383 dvss.n554 dvss.t132 52.8576
R384 dvss.n554 dvss.t153 51.4291
R385 dvss.t154 dvss 42.227
R386 dvss.n195 dvss.n187 41.7862
R387 dvss.t154 dvss.n187 41.7862
R388 dvss.n194 dvss.n186 41.7862
R389 dvss.t154 dvss.n186 41.7862
R390 dvss.n43 dvss.n42 41.7862
R391 dvss.n44 dvss.n43 41.7862
R392 dvss.n37 dvss.n36 41.7862
R393 dvss.n36 dvss.n0 41.7862
R394 dvss.n51 dvss.n50 41.7862
R395 dvss.n52 dvss.n51 41.7862
R396 dvss.n48 dvss.n47 41.7862
R397 dvss.n47 dvss.n46 41.7862
R398 dvss.n553 dvss.n552 40.0735
R399 dvss.n207 dvss.t126 38.5719
R400 dvss.n207 dvss.t3 38.5719
R401 dvss.n224 dvss.t69 38.5719
R402 dvss.n224 dvss.t13 38.5719
R403 dvss.n241 dvss.t42 38.5719
R404 dvss.n241 dvss.t143 38.5719
R405 dvss.n143 dvss.t149 38.5719
R406 dvss.n143 dvss.t17 38.5719
R407 dvss.n160 dvss.t7 38.5719
R408 dvss.n160 dvss.t59 38.5719
R409 dvss.n178 dvss.t71 38.5719
R410 dvss.n178 dvss.t49 38.5719
R411 dvss.n108 dvss.n91 37.6894
R412 dvss.n70 dvss.n69 37.4862
R413 dvss.t173 dvss.t33 36.179
R414 dvss.n82 dvss.n59 36.179
R415 dvss.n6 dvss.t151 36.0005
R416 dvss.n546 dvss.n5 34.6358
R417 dvss.n547 dvss.n546 34.6358
R418 dvss.n548 dvss.n547 34.6358
R419 dvss.n388 dvss.n204 34.6358
R420 dvss.n381 dvss.n205 34.6358
R421 dvss.n364 dvss.n212 34.6358
R422 dvss.n365 dvss.n364 34.6358
R423 dvss.n366 dvss.n365 34.6358
R424 dvss.n366 dvss.n210 34.6358
R425 dvss.n370 dvss.n210 34.6358
R426 dvss.n352 dvss.n214 34.6358
R427 dvss.n356 dvss.n214 34.6358
R428 dvss.n357 dvss.n356 34.6358
R429 dvss.n360 dvss.n357 34.6358
R430 dvss.n339 dvss.n338 34.6358
R431 dvss.n343 dvss.n342 34.6358
R432 dvss.n345 dvss.n343 34.6358
R433 dvss.n349 dvss.n217 34.6358
R434 dvss.n350 dvss.n349 34.6358
R435 dvss.n324 dvss.n229 34.6358
R436 dvss.n325 dvss.n324 34.6358
R437 dvss.n326 dvss.n325 34.6358
R438 dvss.n326 dvss.n227 34.6358
R439 dvss.n330 dvss.n227 34.6358
R440 dvss.n312 dvss.n231 34.6358
R441 dvss.n316 dvss.n231 34.6358
R442 dvss.n317 dvss.n316 34.6358
R443 dvss.n320 dvss.n317 34.6358
R444 dvss.n299 dvss.n298 34.6358
R445 dvss.n303 dvss.n302 34.6358
R446 dvss.n305 dvss.n303 34.6358
R447 dvss.n309 dvss.n234 34.6358
R448 dvss.n310 dvss.n309 34.6358
R449 dvss.n284 dvss.n246 34.6358
R450 dvss.n285 dvss.n284 34.6358
R451 dvss.n286 dvss.n285 34.6358
R452 dvss.n286 dvss.n244 34.6358
R453 dvss.n290 dvss.n244 34.6358
R454 dvss.n272 dvss.n248 34.6358
R455 dvss.n276 dvss.n248 34.6358
R456 dvss.n277 dvss.n276 34.6358
R457 dvss.n280 dvss.n277 34.6358
R458 dvss.n259 dvss.n258 34.6358
R459 dvss.n263 dvss.n262 34.6358
R460 dvss.n265 dvss.n263 34.6358
R461 dvss.n269 dvss.n251 34.6358
R462 dvss.n270 dvss.n269 34.6358
R463 dvss.n521 dvss.n127 34.6358
R464 dvss.n517 dvss.n516 34.6358
R465 dvss.n516 dvss.n515 34.6358
R466 dvss.n512 dvss.n511 34.6358
R467 dvss.n511 dvss.n510 34.6358
R468 dvss.n507 dvss.n506 34.6358
R469 dvss.n506 dvss.n505 34.6358
R470 dvss.n505 dvss.n136 34.6358
R471 dvss.n501 dvss.n136 34.6358
R472 dvss.n499 dvss.n498 34.6358
R473 dvss.n498 dvss.n139 34.6358
R474 dvss.n494 dvss.n139 34.6358
R475 dvss.n494 dvss.n493 34.6358
R476 dvss.n493 dvss.n492 34.6358
R477 dvss.n482 dvss.n481 34.6358
R478 dvss.n479 dvss.n147 34.6358
R479 dvss.n475 dvss.n147 34.6358
R480 dvss.n473 dvss.n472 34.6358
R481 dvss.n472 dvss.n149 34.6358
R482 dvss.n468 dvss.n467 34.6358
R483 dvss.n467 dvss.n466 34.6358
R484 dvss.n466 dvss.n153 34.6358
R485 dvss.n462 dvss.n153 34.6358
R486 dvss.n460 dvss.n459 34.6358
R487 dvss.n459 dvss.n156 34.6358
R488 dvss.n455 dvss.n156 34.6358
R489 dvss.n455 dvss.n454 34.6358
R490 dvss.n454 dvss.n453 34.6358
R491 dvss.n443 dvss.n442 34.6358
R492 dvss.n440 dvss.n164 34.6358
R493 dvss.n436 dvss.n164 34.6358
R494 dvss.n434 dvss.n433 34.6358
R495 dvss.n433 dvss.n166 34.6358
R496 dvss.n429 dvss.n428 34.6358
R497 dvss.n428 dvss.n170 34.6358
R498 dvss.n424 dvss.n170 34.6358
R499 dvss.n424 dvss.n423 34.6358
R500 dvss.n421 dvss.n173 34.6358
R501 dvss.n417 dvss.n173 34.6358
R502 dvss.n417 dvss.n416 34.6358
R503 dvss.n416 dvss.n175 34.6358
R504 dvss.n410 dvss.n175 34.6358
R505 dvss.n402 dvss.n182 34.6358
R506 dvss.n397 dvss.n396 34.6358
R507 dvss.n76 dvss.t137 33.462
R508 dvss.n76 dvss.t195 33.462
R509 dvss.n101 dvss.t110 33.462
R510 dvss.n101 dvss.t171 33.462
R511 dvss.n2 dvss.t9 33.2313
R512 dvss.n342 dvss.n220 31.2476
R513 dvss.n302 dvss.n237 31.2476
R514 dvss.n262 dvss.n254 31.2476
R515 dvss.n517 dvss.n130 31.2476
R516 dvss.n480 dvss.n479 31.2476
R517 dvss.n441 dvss.n440 31.2476
R518 dvss.t8 dvss.t131 30.4092
R519 dvss dvss.n557 30.4092
R520 dvss.n372 dvss.n371 29.7417
R521 dvss.n332 dvss.n331 29.7417
R522 dvss.n292 dvss.n291 29.7417
R523 dvss.n488 dvss.n141 29.7417
R524 dvss.n449 dvss.n158 29.7417
R525 dvss.n409 dvss.n408 29.7417
R526 dvss.n344 dvss.n217 27.8593
R527 dvss.n304 dvss.n234 27.8593
R528 dvss.n264 dvss.n251 27.8593
R529 dvss.n512 dvss.n131 27.8593
R530 dvss.n474 dvss.n473 27.8593
R531 dvss.n435 dvss.n434 27.8593
R532 dvss.n552 dvss.n3 25.977
R533 dvss.n219 dvss.t166 25.4291
R534 dvss.n236 dvss.t77 25.4291
R535 dvss.n253 dvss.t130 25.4291
R536 dvss.n129 dvss.t147 25.4291
R537 dvss.n146 dvss.t82 25.4291
R538 dvss.n163 dvss.t194 25.4291
R539 dvss.n2 dvss.t141 24.9236
R540 dvss.n6 dvss.t60 24.9236
R541 dvss.n25 dvss.n17 24.3755
R542 dvss.n45 dvss.n17 24.3755
R543 dvss.n49 dvss.n18 24.3755
R544 dvss.n45 dvss.n18 24.3755
R545 dvss.n384 dvss.n204 23.7737
R546 dvss.n398 dvss.n397 23.7737
R547 dvss.n81 dvss.n80 23.7181
R548 dvss.n541 dvss.n7 23.7181
R549 dvss.n389 dvss.n388 23.7181
R550 dvss.n377 dvss.n205 23.7181
R551 dvss.n377 dvss.n376 23.7181
R552 dvss.n338 dvss.n337 23.7181
R553 dvss.n337 dvss.n336 23.7181
R554 dvss.n298 dvss.n297 23.7181
R555 dvss.n297 dvss.n296 23.7181
R556 dvss.n258 dvss.n257 23.7181
R557 dvss.n522 dvss.n521 23.7181
R558 dvss.n486 dvss.n144 23.7181
R559 dvss.n482 dvss.n144 23.7181
R560 dvss.n447 dvss.n161 23.7181
R561 dvss.n443 dvss.n161 23.7181
R562 dvss.n404 dvss.n403 23.7181
R563 dvss.n403 dvss.n402 23.7181
R564 dvss.n396 dvss.n393 23.7181
R565 dvss.n105 dvss.n104 23.7181
R566 dvss.n542 dvss.n5 22.9652
R567 dvss.n372 dvss.n208 22.9652
R568 dvss.n332 dvss.n225 22.9652
R569 dvss.n292 dvss.n242 22.9652
R570 dvss.n488 dvss.n487 22.9652
R571 dvss.n449 dvss.n448 22.9652
R572 dvss.n408 dvss.n179 22.9652
R573 dvss.n542 dvss.n541 21.4593
R574 dvss.n376 dvss.n208 21.4593
R575 dvss.n336 dvss.n225 21.4593
R576 dvss.n296 dvss.n242 21.4593
R577 dvss.n487 dvss.n486 21.4593
R578 dvss.n448 dvss.n447 21.4593
R579 dvss.n404 dvss.n179 21.4593
R580 dvss.n556 dvss.n555 21.4265
R581 dvss.n48 dvss.t210 21.1687
R582 dvss.n50 dvss.t36 21.1687
R583 dvss.n199 dvss.t8 21.1543
R584 dvss.n383 dvss.n381 20.9718
R585 dvss.n185 dvss.n182 20.9718
R586 dvss.n33 dvss.n9 19.9405
R587 dvss.n23 dvss.n19 18.4515
R588 dvss.n22 dvss.n20 18.4515
R589 dvss.n28 dvss.n27 18.4515
R590 dvss.n29 dvss.n26 18.4515
R591 dvss.n548 dvss.n3 18.4476
R592 dvss.n351 dvss.n350 17.6946
R593 dvss.n311 dvss.n310 17.6946
R594 dvss.n271 dvss.n270 17.6946
R595 dvss.n510 dvss.n134 17.6946
R596 dvss.n152 dvss.n149 17.6946
R597 dvss.n169 dvss.n166 17.6946
R598 dvss.n112 dvss.t72 16.6567
R599 dvss.n77 dvss 15.0593
R600 dvss.n102 dvss 15.0593
R601 dvss.n371 dvss.n370 14.6829
R602 dvss.n331 dvss.n330 14.6829
R603 dvss.n291 dvss.n290 14.6829
R604 dvss.n492 dvss.n141 14.6829
R605 dvss.n453 dvss.n158 14.6829
R606 dvss.n410 dvss.n409 14.6829
R607 dvss.t136 dvss.n59 13.7828
R608 dvss.n40 dvss.n9 13.3461
R609 dvss.n39 dvss.n38 13.0158
R610 dvss.n34 dvss.n33 11.7338
R611 dvss.n41 dvss.n40 10.1755
R612 dvss.n120 dvss 9.488
R613 dvss.n80 dvss.n79 9.3005
R614 dvss.n81 dvss.n60 9.3005
R615 dvss.n394 dvss.n393 9.3005
R616 dvss.n412 dvss.n175 9.3005
R617 dvss.n411 dvss.n410 9.3005
R618 dvss.n409 dvss.n177 9.3005
R619 dvss.n408 dvss.n407 9.3005
R620 dvss.n406 dvss.n179 9.3005
R621 dvss.n405 dvss.n404 9.3005
R622 dvss.n403 dvss.n181 9.3005
R623 dvss.n402 dvss.n401 9.3005
R624 dvss.n400 dvss.n182 9.3005
R625 dvss.n399 dvss.n398 9.3005
R626 dvss.n397 dvss.n183 9.3005
R627 dvss.n396 dvss.n395 9.3005
R628 dvss.n522 dvss.n126 9.3005
R629 dvss.n521 dvss.n520 9.3005
R630 dvss.n519 dvss.n127 9.3005
R631 dvss.n518 dvss.n517 9.3005
R632 dvss.n516 dvss.n128 9.3005
R633 dvss.n515 dvss.n514 9.3005
R634 dvss.n513 dvss.n512 9.3005
R635 dvss.n511 dvss.n132 9.3005
R636 dvss.n510 dvss.n509 9.3005
R637 dvss.n508 dvss.n507 9.3005
R638 dvss.n506 dvss.n135 9.3005
R639 dvss.n505 dvss.n504 9.3005
R640 dvss.n503 dvss.n136 9.3005
R641 dvss.n502 dvss.n501 9.3005
R642 dvss.n499 dvss.n137 9.3005
R643 dvss.n498 dvss.n497 9.3005
R644 dvss.n496 dvss.n139 9.3005
R645 dvss.n495 dvss.n494 9.3005
R646 dvss.n493 dvss.n140 9.3005
R647 dvss.n492 dvss.n491 9.3005
R648 dvss.n490 dvss.n141 9.3005
R649 dvss.n489 dvss.n488 9.3005
R650 dvss.n487 dvss.n142 9.3005
R651 dvss.n486 dvss.n485 9.3005
R652 dvss.n484 dvss.n144 9.3005
R653 dvss.n483 dvss.n482 9.3005
R654 dvss.n481 dvss.n145 9.3005
R655 dvss.n479 dvss.n478 9.3005
R656 dvss.n477 dvss.n147 9.3005
R657 dvss.n476 dvss.n475 9.3005
R658 dvss.n473 dvss.n148 9.3005
R659 dvss.n472 dvss.n471 9.3005
R660 dvss.n470 dvss.n149 9.3005
R661 dvss.n469 dvss.n468 9.3005
R662 dvss.n467 dvss.n150 9.3005
R663 dvss.n466 dvss.n465 9.3005
R664 dvss.n464 dvss.n153 9.3005
R665 dvss.n463 dvss.n462 9.3005
R666 dvss.n460 dvss.n154 9.3005
R667 dvss.n459 dvss.n458 9.3005
R668 dvss.n457 dvss.n156 9.3005
R669 dvss.n456 dvss.n455 9.3005
R670 dvss.n454 dvss.n157 9.3005
R671 dvss.n453 dvss.n452 9.3005
R672 dvss.n451 dvss.n158 9.3005
R673 dvss.n450 dvss.n449 9.3005
R674 dvss.n448 dvss.n159 9.3005
R675 dvss.n447 dvss.n446 9.3005
R676 dvss.n445 dvss.n161 9.3005
R677 dvss.n444 dvss.n443 9.3005
R678 dvss.n442 dvss.n162 9.3005
R679 dvss.n440 dvss.n439 9.3005
R680 dvss.n438 dvss.n164 9.3005
R681 dvss.n437 dvss.n436 9.3005
R682 dvss.n434 dvss.n165 9.3005
R683 dvss.n433 dvss.n432 9.3005
R684 dvss.n431 dvss.n166 9.3005
R685 dvss.n430 dvss.n429 9.3005
R686 dvss.n428 dvss.n427 9.3005
R687 dvss.n426 dvss.n170 9.3005
R688 dvss.n425 dvss.n424 9.3005
R689 dvss.n423 dvss.n171 9.3005
R690 dvss.n421 dvss.n420 9.3005
R691 dvss.n419 dvss.n173 9.3005
R692 dvss.n418 dvss.n417 9.3005
R693 dvss.n416 dvss.n415 9.3005
R694 dvss.n257 dvss.n256 9.3005
R695 dvss.n258 dvss.n255 9.3005
R696 dvss.n260 dvss.n259 9.3005
R697 dvss.n262 dvss.n261 9.3005
R698 dvss.n263 dvss.n252 9.3005
R699 dvss.n266 dvss.n265 9.3005
R700 dvss.n267 dvss.n251 9.3005
R701 dvss.n269 dvss.n268 9.3005
R702 dvss.n270 dvss.n249 9.3005
R703 dvss.n273 dvss.n272 9.3005
R704 dvss.n274 dvss.n248 9.3005
R705 dvss.n276 dvss.n275 9.3005
R706 dvss.n277 dvss.n247 9.3005
R707 dvss.n281 dvss.n280 9.3005
R708 dvss.n282 dvss.n246 9.3005
R709 dvss.n284 dvss.n283 9.3005
R710 dvss.n285 dvss.n245 9.3005
R711 dvss.n287 dvss.n286 9.3005
R712 dvss.n288 dvss.n244 9.3005
R713 dvss.n290 dvss.n289 9.3005
R714 dvss.n291 dvss.n243 9.3005
R715 dvss.n293 dvss.n292 9.3005
R716 dvss.n294 dvss.n242 9.3005
R717 dvss.n296 dvss.n295 9.3005
R718 dvss.n297 dvss.n239 9.3005
R719 dvss.n298 dvss.n238 9.3005
R720 dvss.n300 dvss.n299 9.3005
R721 dvss.n302 dvss.n301 9.3005
R722 dvss.n303 dvss.n235 9.3005
R723 dvss.n306 dvss.n305 9.3005
R724 dvss.n307 dvss.n234 9.3005
R725 dvss.n309 dvss.n308 9.3005
R726 dvss.n310 dvss.n232 9.3005
R727 dvss.n313 dvss.n312 9.3005
R728 dvss.n314 dvss.n231 9.3005
R729 dvss.n316 dvss.n315 9.3005
R730 dvss.n317 dvss.n230 9.3005
R731 dvss.n321 dvss.n320 9.3005
R732 dvss.n322 dvss.n229 9.3005
R733 dvss.n324 dvss.n323 9.3005
R734 dvss.n325 dvss.n228 9.3005
R735 dvss.n327 dvss.n326 9.3005
R736 dvss.n328 dvss.n227 9.3005
R737 dvss.n330 dvss.n329 9.3005
R738 dvss.n331 dvss.n226 9.3005
R739 dvss.n333 dvss.n332 9.3005
R740 dvss.n334 dvss.n225 9.3005
R741 dvss.n336 dvss.n335 9.3005
R742 dvss.n337 dvss.n222 9.3005
R743 dvss.n338 dvss.n221 9.3005
R744 dvss.n340 dvss.n339 9.3005
R745 dvss.n342 dvss.n341 9.3005
R746 dvss.n343 dvss.n218 9.3005
R747 dvss.n346 dvss.n345 9.3005
R748 dvss.n347 dvss.n217 9.3005
R749 dvss.n349 dvss.n348 9.3005
R750 dvss.n350 dvss.n215 9.3005
R751 dvss.n353 dvss.n352 9.3005
R752 dvss.n354 dvss.n214 9.3005
R753 dvss.n356 dvss.n355 9.3005
R754 dvss.n357 dvss.n213 9.3005
R755 dvss.n361 dvss.n360 9.3005
R756 dvss.n362 dvss.n212 9.3005
R757 dvss.n364 dvss.n363 9.3005
R758 dvss.n365 dvss.n211 9.3005
R759 dvss.n367 dvss.n366 9.3005
R760 dvss.n368 dvss.n210 9.3005
R761 dvss.n370 dvss.n369 9.3005
R762 dvss.n371 dvss.n209 9.3005
R763 dvss.n373 dvss.n372 9.3005
R764 dvss.n374 dvss.n208 9.3005
R765 dvss.n376 dvss.n375 9.3005
R766 dvss.n378 dvss.n377 9.3005
R767 dvss.n379 dvss.n205 9.3005
R768 dvss.n381 dvss.n380 9.3005
R769 dvss.n385 dvss.n384 9.3005
R770 dvss.n386 dvss.n204 9.3005
R771 dvss.n388 dvss.n387 9.3005
R772 dvss.n389 dvss.n203 9.3005
R773 dvss.n538 dvss.n7 9.3005
R774 dvss.n543 dvss.n542 9.3005
R775 dvss.n549 dvss.n548 9.3005
R776 dvss.n547 dvss.n4 9.3005
R777 dvss.n546 dvss.n545 9.3005
R778 dvss.n544 dvss.n5 9.3005
R779 dvss.n541 dvss.n540 9.3005
R780 dvss.n550 dvss.n3 9.3005
R781 dvss.n552 dvss.n551 9.3005
R782 dvss.n106 dvss.n105 9.3005
R783 dvss.n104 dvss.n103 9.3005
R784 dvss.n98 dvss.n13 9.3005
R785 dvss.n531 dvss.n530 9.3005
R786 dvss.n73 dvss.n56 9.3005
R787 dvss.n109 dvss.n108 8.88939
R788 dvss.n69 dvss.n68 8.77764
R789 dvss.n359 dvss.n212 7.90638
R790 dvss.n319 dvss.n229 7.90638
R791 dvss.n279 dvss.n246 7.90638
R792 dvss.n500 dvss.n499 7.90638
R793 dvss.n461 dvss.n460 7.90638
R794 dvss.n422 dvss.n421 7.90638
R795 dvss.n103 dvss.n102 7.18226
R796 dvss.n78 dvss.n77 7.17078
R797 dvss.n80 dvss 7.15344
R798 dvss.n104 dvss 7.15344
R799 dvss.n345 dvss.n344 6.77697
R800 dvss.n305 dvss.n304 6.77697
R801 dvss.n265 dvss.n264 6.77697
R802 dvss.n515 dvss.n131 6.77697
R803 dvss.n475 dvss.n474 6.77697
R804 dvss.n436 dvss.n435 6.77697
R805 dvss.n195 dvss.n176 6.7005
R806 dvss.n555 dvss.n553 6.56103
R807 dvss.n41 dvss.n35 5.66204
R808 dvss.n39 dvss.n35 5.19708
R809 dvss.n19 dvss.t208 4.3505
R810 dvss.n19 dvss.t106 4.3505
R811 dvss.n20 dvss.t134 4.3505
R812 dvss.n20 dvss.t200 4.3505
R813 dvss.n27 dvss.t57 4.3505
R814 dvss.n27 dvss.t102 4.3505
R815 dvss.n26 dvss.t108 4.3505
R816 dvss.n26 dvss.t38 4.3505
R817 dvss.n339 dvss.n220 3.38874
R818 dvss.n299 dvss.n237 3.38874
R819 dvss.n259 dvss.n254 3.38874
R820 dvss.n130 dvss.n127 3.38874
R821 dvss.n481 dvss.n480 3.38874
R822 dvss.n442 dvss.n441 3.38874
R823 dvss.n542 dvss 3.29747
R824 dvss.n556 dvss.n1 3.21038
R825 dvss.n75 dvss.n70 3.17391
R826 dvss.n352 dvss.n351 2.63579
R827 dvss.n312 dvss.n311 2.63579
R828 dvss.n272 dvss.n271 2.63579
R829 dvss.n507 dvss.n134 2.63579
R830 dvss.n468 dvss.n152 2.63579
R831 dvss.n429 dvss.n169 2.63579
R832 dvss.n40 dvss.n39 2.50662
R833 dvss.n107 dvss.n95 2.44193
R834 dvss.n69 dvss.n60 2.41042
R835 dvss.n108 dvss.n107 2.3255
R836 dvss.n553 dvss.n1 1.93239
R837 dvss.n360 dvss.n359 1.88285
R838 dvss.n320 dvss.n319 1.88285
R839 dvss.n280 dvss.n279 1.88285
R840 dvss.n501 dvss.n500 1.88285
R841 dvss.n462 dvss.n461 1.88285
R842 dvss.n423 dvss.n422 1.88285
R843 dvss.n38 dvss.n37 1.85983
R844 dvss.n24 dvss.n23 1.57196
R845 dvss.n30 dvss.n29 1.57139
R846 dvss.n188 dvss.n174 1.5505
R847 dvss.n70 dvss.n61 1.46336
R848 dvss.n529 dvss.n14 1.32907
R849 dvss.n121 dvss.n57 1.32907
R850 dvss.n414 dvss.n176 1.11858
R851 dvss.n193 dvss.n188 0.649775
R852 dvss dvss.n119 0.637219
R853 dvss.n384 dvss.n383 0.630008
R854 dvss.n398 dvss.n185 0.630008
R855 dvss.t61 dvss.n533 0.474702
R856 dvss.n533 dvss 0.36436
R857 dvss.n533 dvss.n532 0.357983
R858 dvss.n38 dvss 0.326572
R859 dvss.n538 dvss.n537 0.274194
R860 dvss.n100 dvss.n99 0.260009
R861 dvss.n256 dvss.n126 0.240996
R862 dvss.n167 dvss.t88 0.189075
R863 dvss.n74 dvss 0.178871
R864 dvss.n95 dvss.n91 0.178278
R865 dvss dvss.n536 0.150986
R866 dvss.n532 dvss.n531 0.148545
R867 dvss.n72 dvss 0.145311
R868 dvss.n413 dvss 0.142307
R869 dvss.n201 dvss 0.140841
R870 dvss.n99 dvss 0.140381
R871 dvss.n531 dvss.n11 0.136163
R872 dvss.n536 dvss.n535 0.13579
R873 dvss.n202 dvss 0.127978
R874 dvss.n202 dvss.n201 0.123227
R875 dvss.n412 dvss.n411 0.120292
R876 dvss.n411 dvss.n177 0.120292
R877 dvss.n407 dvss.n177 0.120292
R878 dvss.n407 dvss.n406 0.120292
R879 dvss.n406 dvss.n405 0.120292
R880 dvss.n401 dvss.n400 0.120292
R881 dvss.n399 dvss.n183 0.120292
R882 dvss.n395 dvss.n183 0.120292
R883 dvss.n544 dvss.n543 0.120292
R884 dvss.n545 dvss.n544 0.120292
R885 dvss.n545 dvss.n4 0.120292
R886 dvss.n549 dvss.n4 0.120292
R887 dvss.n550 dvss.n549 0.120292
R888 dvss.n551 dvss.n550 0.120292
R889 dvss.n97 dvss 0.115052
R890 dvss.n119 dvss.n118 0.109875
R891 dvss.n75 dvss.n74 0.109468
R892 dvss.n400 dvss 0.104667
R893 dvss.n414 dvss 0.0999624
R894 dvss.n543 dvss 0.0968542
R895 dvss.n100 dvss 0.0959969
R896 dvss.n78 dvss 0.080434
R897 dvss.n200 dvss 0.0781256
R898 dvss.n79 dvss.n78 0.0777204
R899 dvss.t87 dvss.t62 0.070611
R900 dvss.n50 dvss.n24 0.0678684
R901 dvss.n534 dvss.t61 0.0675999
R902 dvss.n48 dvss.n30 0.0671667
R903 dvss.n536 dvss.n9 0.0664942
R904 dvss.n201 dvss.n200 0.0638562
R905 dvss.n21 dvss 0.0633141
R906 dvss.n118 dvss.n57 0.0606266
R907 dvss.n532 dvss 0.060557
R908 dvss.n535 dvss.t88 0.060491
R909 dvss.n181 dvss 0.0603958
R910 dvss.n401 dvss 0.0603958
R911 dvss dvss.n394 0.0603958
R912 dvss.n540 dvss 0.0603958
R913 dvss.n72 dvss.n71 0.0603629
R914 dvss.n200 dvss.n8 0.0586797
R915 dvss.n1 dvss 0.0525833
R916 dvss.n14 dvss.n11 0.0495635
R917 dvss.n107 dvss.n106 0.0482484
R918 dvss.n97 dvss.n96 0.0467134
R919 dvss.n29 dvss.n28 0.0457733
R920 dvss.n413 dvss.n412 0.0447708
R921 dvss.n118 dvss 0.0421667
R922 dvss.n534 dvss.n10 0.0405094
R923 dvss.n23 dvss 0.0346686
R924 dvss dvss.n100 0.0335285
R925 dvss dvss.n181 0.0330521
R926 dvss.n394 dvss 0.0330521
R927 dvss.n11 dvss 0.0300195
R928 dvss.n74 dvss.n73 0.028566
R929 dvss dvss.n538 0.0271393
R930 dvss.n103 dvss 0.0248902
R931 dvss.n540 dvss 0.0239375
R932 dvss.n28 dvss.n10 0.0228519
R933 dvss.n405 dvss 0.0226354
R934 dvss.n395 dvss 0.0226354
R935 dvss.n75 dvss 0.0215598
R936 dvss.n99 dvss.n98 0.0208358
R937 dvss.n8 dvss 0.0206613
R938 dvss.n539 dvss 0.0199672
R939 dvss.n119 dvss 0.0193397
R940 dvss.n22 dvss.n21 0.0184385
R941 dvss dvss.n60 0.0174837
R942 dvss dvss.n399 0.016125
R943 dvss.n520 dvss.n519 0.015957
R944 dvss.n519 dvss.n518 0.015957
R945 dvss.n518 dvss.n128 0.015957
R946 dvss.n514 dvss.n128 0.015957
R947 dvss.n514 dvss.n513 0.015957
R948 dvss.n513 dvss.n132 0.015957
R949 dvss.n509 dvss.n132 0.015957
R950 dvss.n509 dvss.n508 0.015957
R951 dvss.n508 dvss.n135 0.015957
R952 dvss.n504 dvss.n135 0.015957
R953 dvss.n504 dvss.n503 0.015957
R954 dvss.n503 dvss.n502 0.015957
R955 dvss.n502 dvss.n137 0.015957
R956 dvss.n497 dvss.n137 0.015957
R957 dvss.n497 dvss.n496 0.015957
R958 dvss.n496 dvss.n495 0.015957
R959 dvss.n495 dvss.n140 0.015957
R960 dvss.n491 dvss.n140 0.015957
R961 dvss.n491 dvss.n490 0.015957
R962 dvss.n490 dvss.n489 0.015957
R963 dvss.n489 dvss.n142 0.015957
R964 dvss.n485 dvss.n142 0.015957
R965 dvss.n483 dvss.n145 0.015957
R966 dvss.n478 dvss.n145 0.015957
R967 dvss.n478 dvss.n477 0.015957
R968 dvss.n477 dvss.n476 0.015957
R969 dvss.n476 dvss.n148 0.015957
R970 dvss.n471 dvss.n148 0.015957
R971 dvss.n471 dvss.n470 0.015957
R972 dvss.n470 dvss.n469 0.015957
R973 dvss.n469 dvss.n150 0.015957
R974 dvss.n465 dvss.n150 0.015957
R975 dvss.n465 dvss.n464 0.015957
R976 dvss.n464 dvss.n463 0.015957
R977 dvss.n463 dvss.n154 0.015957
R978 dvss.n458 dvss.n154 0.015957
R979 dvss.n458 dvss.n457 0.015957
R980 dvss.n457 dvss.n456 0.015957
R981 dvss.n456 dvss.n157 0.015957
R982 dvss.n452 dvss.n157 0.015957
R983 dvss.n452 dvss.n451 0.015957
R984 dvss.n451 dvss.n450 0.015957
R985 dvss.n450 dvss.n159 0.015957
R986 dvss.n446 dvss.n159 0.015957
R987 dvss.n444 dvss.n162 0.015957
R988 dvss.n439 dvss.n162 0.015957
R989 dvss.n439 dvss.n438 0.015957
R990 dvss.n438 dvss.n437 0.015957
R991 dvss.n437 dvss.n165 0.015957
R992 dvss.n432 dvss.n165 0.015957
R993 dvss.n432 dvss.n431 0.015957
R994 dvss.n431 dvss.n430 0.015957
R995 dvss.n427 dvss.n426 0.015957
R996 dvss.n426 dvss.n425 0.015957
R997 dvss.n425 dvss.n171 0.015957
R998 dvss.n420 dvss.n171 0.015957
R999 dvss.n420 dvss.n419 0.015957
R1000 dvss.n419 dvss.n418 0.015957
R1001 dvss.n414 dvss.n413 0.0141555
R1002 dvss.n260 dvss.n255 0.0125293
R1003 dvss.n261 dvss.n260 0.0125293
R1004 dvss.n261 dvss.n252 0.0125293
R1005 dvss.n266 dvss.n252 0.0125293
R1006 dvss.n267 dvss.n266 0.0125293
R1007 dvss.n268 dvss.n267 0.0125293
R1008 dvss.n268 dvss.n249 0.0125293
R1009 dvss.n273 dvss.n249 0.0125293
R1010 dvss.n274 dvss.n273 0.0125293
R1011 dvss.n275 dvss.n274 0.0125293
R1012 dvss.n275 dvss.n247 0.0125293
R1013 dvss.n281 dvss.n247 0.0125293
R1014 dvss.n282 dvss.n281 0.0125293
R1015 dvss.n283 dvss.n282 0.0125293
R1016 dvss.n283 dvss.n245 0.0125293
R1017 dvss.n287 dvss.n245 0.0125293
R1018 dvss.n288 dvss.n287 0.0125293
R1019 dvss.n289 dvss.n288 0.0125293
R1020 dvss.n289 dvss.n243 0.0125293
R1021 dvss.n293 dvss.n243 0.0125293
R1022 dvss.n294 dvss.n293 0.0125293
R1023 dvss.n295 dvss.n294 0.0125293
R1024 dvss.n300 dvss.n238 0.0125293
R1025 dvss.n301 dvss.n300 0.0125293
R1026 dvss.n301 dvss.n235 0.0125293
R1027 dvss.n306 dvss.n235 0.0125293
R1028 dvss.n307 dvss.n306 0.0125293
R1029 dvss.n308 dvss.n307 0.0125293
R1030 dvss.n308 dvss.n232 0.0125293
R1031 dvss.n313 dvss.n232 0.0125293
R1032 dvss.n314 dvss.n313 0.0125293
R1033 dvss.n315 dvss.n314 0.0125293
R1034 dvss.n315 dvss.n230 0.0125293
R1035 dvss.n321 dvss.n230 0.0125293
R1036 dvss.n322 dvss.n321 0.0125293
R1037 dvss.n323 dvss.n322 0.0125293
R1038 dvss.n323 dvss.n228 0.0125293
R1039 dvss.n327 dvss.n228 0.0125293
R1040 dvss.n328 dvss.n327 0.0125293
R1041 dvss.n329 dvss.n328 0.0125293
R1042 dvss.n329 dvss.n226 0.0125293
R1043 dvss.n333 dvss.n226 0.0125293
R1044 dvss.n334 dvss.n333 0.0125293
R1045 dvss.n335 dvss.n334 0.0125293
R1046 dvss.n340 dvss.n221 0.0125293
R1047 dvss.n341 dvss.n340 0.0125293
R1048 dvss.n341 dvss.n218 0.0125293
R1049 dvss.n346 dvss.n218 0.0125293
R1050 dvss.n347 dvss.n346 0.0125293
R1051 dvss.n348 dvss.n347 0.0125293
R1052 dvss.n348 dvss.n215 0.0125293
R1053 dvss.n353 dvss.n215 0.0125293
R1054 dvss.n354 dvss.n353 0.0125293
R1055 dvss.n355 dvss.n354 0.0125293
R1056 dvss.n355 dvss.n213 0.0125293
R1057 dvss.n361 dvss.n213 0.0125293
R1058 dvss.n362 dvss.n361 0.0125293
R1059 dvss.n363 dvss.n362 0.0125293
R1060 dvss.n363 dvss.n211 0.0125293
R1061 dvss.n367 dvss.n211 0.0125293
R1062 dvss.n368 dvss.n367 0.0125293
R1063 dvss.n369 dvss.n368 0.0125293
R1064 dvss.n369 dvss.n209 0.0125293
R1065 dvss.n373 dvss.n209 0.0125293
R1066 dvss.n374 dvss.n373 0.0125293
R1067 dvss.n375 dvss.n374 0.0125293
R1068 dvss.n380 dvss.n379 0.0125293
R1069 dvss.n386 dvss.n385 0.0125293
R1070 dvss.n387 dvss.n386 0.0125293
R1071 dvss.n427 dvss.n167 0.0122608
R1072 dvss.n100 dvss 0.012146
R1073 dvss dvss.n22 0.0110353
R1074 dvss.n380 dvss 0.0109603
R1075 dvss.n79 dvss.n75 0.0106902
R1076 dvss.n535 dvss.t87 0.0106199
R1077 dvss.n106 dvss 0.0105932
R1078 dvss.n415 dvss.n174 0.0099086
R1079 dvss.n537 dvss.n8 0.00990439
R1080 dvss.n551 dvss.n1 0.0083125
R1081 dvss.n520 dvss 0.00822849
R1082 dvss dvss.n484 0.00822849
R1083 dvss dvss.n483 0.00822849
R1084 dvss dvss.n445 0.00822849
R1085 dvss dvss.n444 0.00822849
R1086 dvss.n73 dvss.n72 0.00733962
R1087 dvss.n418 dvss.n174 0.00654839
R1088 dvss dvss.n255 0.00651464
R1089 dvss dvss.n239 0.00651464
R1090 dvss dvss.n238 0.00651464
R1091 dvss dvss.n222 0.00651464
R1092 dvss dvss.n221 0.00651464
R1093 dvss.n378 dvss 0.00651464
R1094 dvss.n379 dvss 0.00651464
R1095 dvss dvss.n203 0.00651464
R1096 dvss.n98 dvss.n97 0.00591045
R1097 dvss dvss.n1 0.00570833
R1098 dvss.n21 dvss.n10 0.00519818
R1099 dvss.n537 dvss 0.00481034
R1100 dvss dvss.n126 0.00470027
R1101 dvss.n484 dvss 0.00470027
R1102 dvss.n445 dvss 0.00470027
R1103 dvss.n430 dvss.n167 0.00419624
R1104 dvss.n256 dvss 0.00376883
R1105 dvss.n239 dvss 0.00376883
R1106 dvss.n222 dvss 0.00376883
R1107 dvss dvss.n378 0.00376883
R1108 dvss.n203 dvss 0.00376883
R1109 dvss.t62 dvss.n534 0.00351108
R1110 dvss.n485 dvss 0.00335618
R1111 dvss.n446 dvss 0.00335618
R1112 dvss.n295 dvss 0.0027228
R1113 dvss.n335 dvss 0.0027228
R1114 dvss.n375 dvss 0.0027228
R1115 dvss.n387 dvss 0.0027228
R1116 dvss.n385 dvss 0.00206904
R1117 dvss dvss.n539 0.00180208
R1118 dvss.n539 dvss 0.00152459
R1119 dvss.n415 dvss.n414 0.00150806
R1120 dvss dvss.n202 0.00077533
R1121 dvss.n71 dvss.n57 0.000763713
R1122 dvss.n96 dvss.n14 0.000703583
R1123 x7.stby_done_b.n8 x7.stby_done_b.t1 373.866
R1124 x7.stby_done_b.n6 x7.stby_done_b.t6 333.651
R1125 x7.stby_done_b.n6 x7.stby_done_b.t2 297.233
R1126 x7.stby_done_b.n1 x7.stby_done_b.t5 241.536
R1127 x7.stby_done_b x7.stby_done_b.t0 237.101
R1128 x7.stby_done_b.n4 x7.stby_done_b.t3 207.423
R1129 x7.stby_done_b.n3 x7.stby_done_b.t4 202.133
R1130 x7.stby_done_b x7.stby_done_b.n6 195.701
R1131 x7.stby_done_b.n1 x7.stby_done_b.t7 169.237
R1132 x7.stby_done_b.n5 x7.stby_done_b.n4 159.758
R1133 x7.stby_done_b.n3 x7.stby_done_b 154.91
R1134 x7.stby_done_b.n2 x7.stby_done_b.n1 152
R1135 x7.stby_done_b.n4 x7.stby_done_b.n3 36.8275
R1136 x7.stby_done_b x7.stby_done_b.n8 26.7478
R1137 x7.stby_done_b.n7 x7.stby_done_b 15.8995
R1138 x7.stby_done_b.n7 x7.stby_done_b.n0 15.8481
R1139 x7.stby_done_b.n0 x7.stby_done_b.n5 13.8109
R1140 x7.stby_done_b x7.stby_done_b.n2 13.3943
R1141 x7.stby_done_b.n8 x7.stby_done_b.n7 3.1005
R1142 x7.stby_done_b.n5 x7.stby_done_b 2.52171
R1143 x7.stby_done_b.n2 x7.stby_done_b 1.9205
R1144 x7.stby_done_b.n0 x7.stby_done_b 1.418
R1145 dvdd.n294 dvdd.n285 5128.23
R1146 dvdd.n294 dvdd.n286 5128.23
R1147 dvdd.n292 dvdd.n286 5128.23
R1148 dvdd.n292 dvdd.n285 5128.23
R1149 dvdd.n42 dvdd.n5 1736.47
R1150 dvdd.n45 dvdd.n4 1736.47
R1151 dvdd.n30 dvdd.n27 1736.47
R1152 dvdd.n33 dvdd.n29 1736.47
R1153 dvdd.n254 dvdd.t15 838.817
R1154 dvdd.n69 dvdd.t51 806.511
R1155 dvdd.n69 dvdd.t9 806.511
R1156 dvdd.n90 dvdd.t116 806.511
R1157 dvdd.n90 dvdd.t1 806.511
R1158 dvdd.n111 dvdd.t99 806.511
R1159 dvdd.n111 dvdd.t29 806.511
R1160 dvdd.n291 dvdd.n283 787.447
R1161 dvdd.n291 dvdd.n284 786.827
R1162 dvdd.n56 dvdd.t144 668.683
R1163 dvdd.n56 dvdd.t75 668.683
R1164 dvdd.n227 dvdd.t19 667.778
R1165 dvdd.n227 dvdd.t95 667.778
R1166 dvdd.n189 dvdd.t113 667.778
R1167 dvdd.n189 dvdd.t23 667.778
R1168 dvdd.n151 dvdd.t25 667.778
R1169 dvdd.n151 dvdd.t140 667.778
R1170 dvdd.n295 dvdd.n283 604.574
R1171 dvdd.n73 dvdd.n71 604.457
R1172 dvdd.n73 dvdd.n72 604.457
R1173 dvdd.n94 dvdd.n92 604.457
R1174 dvdd.n94 dvdd.n93 604.457
R1175 dvdd.n115 dvdd.n113 604.457
R1176 dvdd.n115 dvdd.n114 604.457
R1177 dvdd.n232 dvdd.n61 604.394
R1178 dvdd.n232 dvdd.n62 604.394
R1179 dvdd.n194 dvdd.n82 604.394
R1180 dvdd.n194 dvdd.n83 604.394
R1181 dvdd.n156 dvdd.n103 604.394
R1182 dvdd.n156 dvdd.n104 604.394
R1183 dvdd.n220 dvdd.n67 601.679
R1184 dvdd.n220 dvdd.n68 601.679
R1185 dvdd.n182 dvdd.n88 601.679
R1186 dvdd.n182 dvdd.n89 601.679
R1187 dvdd.n144 dvdd.n109 601.679
R1188 dvdd.n144 dvdd.n110 601.679
R1189 dvdd.n259 dvdd.n258 585
R1190 dvdd.t92 dvdd.t14 556.386
R1191 dvdd.n246 dvdd 538.664
R1192 dvdd.n18 dvdd 535.705
R1193 dvdd.n11 dvdd 535.705
R1194 dvdd.t10 dvdd 473.521
R1195 dvdd.t24 dvdd.t81 448.146
R1196 dvdd.t22 dvdd.t4 448.146
R1197 dvdd.t18 dvdd.t12 448.146
R1198 dvdd.n295 dvdd.n284 423.062
R1199 dvdd.t100 dvdd.t58 367.579
R1200 dvdd.t135 dvdd.t145 367.579
R1201 dvdd.t64 dvdd.t66 367.579
R1202 dvdd.n273 dvdd.t52 360.005
R1203 dvdd.t28 dvdd.t61 330.654
R1204 dvdd.t0 dvdd.t16 330.654
R1205 dvdd.t8 dvdd.t106 330.654
R1206 dvdd.n43 dvdd.n4 314.781
R1207 dvdd.n44 dvdd.n5 314.781
R1208 dvdd.n31 dvdd.n29 314.781
R1209 dvdd.n32 dvdd.n27 314.781
R1210 dvdd.n23 dvdd.n17 312.053
R1211 dvdd.n9 dvdd.n8 312.051
R1212 dvdd.n265 dvdd.n255 312.051
R1213 dvdd.t47 dvdd.t45 304.829
R1214 dvdd.t14 dvdd.t137 284.113
R1215 dvdd.t58 dvdd.t86 275.265
R1216 dvdd.t145 dvdd.t111 275.265
R1217 dvdd.t66 dvdd.t125 275.265
R1218 dvdd.t137 dvdd.t10 275.235
R1219 dvdd.n270 dvdd.t33 261.837
R1220 dvdd.t114 dvdd.t127 260.437
R1221 dvdd.t148 dvdd.t108 260.437
R1222 dvdd.n207 dvdd.n76 259.707
R1223 dvdd.n207 dvdd.n75 259.707
R1224 dvdd.n169 dvdd.n97 259.707
R1225 dvdd.n169 dvdd.n96 259.707
R1226 dvdd.n131 dvdd.n118 259.707
R1227 dvdd.n131 dvdd.n117 259.707
R1228 dvdd.t33 dvdd.t26 258.481
R1229 dvdd.n272 dvdd.t129 253.446
R1230 dvdd.n271 dvdd.t133 253.446
R1231 dvdd.t44 dvdd.t124 248.599
R1232 dvdd.t124 dvdd.t92 248.599
R1233 dvdd.n201 dvdd.n80 242.607
R1234 dvdd.n163 dvdd.n101 242.607
R1235 dvdd.n125 dvdd.n123 242.607
R1236 dvdd.n201 dvdd.n79 242.607
R1237 dvdd.n163 dvdd.n100 242.607
R1238 dvdd.n125 dvdd.n122 242.607
R1239 dvdd.t49 dvdd.t142 234.982
R1240 dvdd.t152 dvdd.t7 234.982
R1241 dvdd.t31 dvdd.t63 234.982
R1242 dvdd dvdd.n269 232.445
R1243 dvdd.n0 dvdd.t39 228.215
R1244 dvdd.n0 dvdd.t37 228.215
R1245 dvdd.n239 dvdd.n59 215.123
R1246 dvdd.n239 dvdd.n238 215.123
R1247 dvdd.t45 dvdd.t76 213.084
R1248 dvdd.n41 dvdd.n3 185.225
R1249 dvdd.n46 dvdd.n3 185.225
R1250 dvdd.n34 dvdd.n28 185.225
R1251 dvdd.n28 dvdd.n26 185.225
R1252 dvdd.t102 dvdd.t84 181.273
R1253 dvdd.t72 dvdd.t120 181.273
R1254 dvdd.t90 dvdd.t117 181.273
R1255 dvdd.t57 dvdd.t28 166.167
R1256 dvdd.t142 dvdd.t158 166.167
R1257 dvdd.t6 dvdd.t0 166.167
R1258 dvdd.t7 dvdd.t159 166.167
R1259 dvdd.t110 dvdd.t8 166.167
R1260 dvdd.t63 dvdd.t98 166.167
R1261 dvdd.t52 dvdd.t100 162.81
R1262 dvdd.t61 dvdd.t49 162.81
R1263 dvdd.t129 dvdd.t135 162.81
R1264 dvdd.t16 dvdd.t152 162.81
R1265 dvdd.t133 dvdd.t64 162.81
R1266 dvdd.t106 dvdd.t31 162.81
R1267 dvdd.t68 dvdd.n292 161.316
R1268 dvdd.n294 dvdd.t169 161.316
R1269 dvdd.t158 dvdd.t24 154.417
R1270 dvdd.t159 dvdd.t22 154.417
R1271 dvdd.t98 dvdd.t18 154.417
R1272 dvdd.t26 dvdd.t74 147.703
R1273 dvdd.n75 dvdd.t141 147.111
R1274 dvdd.n76 dvdd.t126 147.111
R1275 dvdd.n96 dvdd.t112 147.111
R1276 dvdd.n97 dvdd.t147 147.111
R1277 dvdd.n117 dvdd.t87 147.111
R1278 dvdd.n118 dvdd.t166 147.111
R1279 dvdd.t83 dvdd.t57 144.346
R1280 dvdd.t96 dvdd.t6 144.346
R1281 dvdd.t97 dvdd.t110 144.346
R1282 dvdd.t86 dvdd.t102 140.989
R1283 dvdd.t84 dvdd.t83 140.989
R1284 dvdd.t81 dvdd.t93 140.989
R1285 dvdd.t111 dvdd.t72 140.989
R1286 dvdd.t120 dvdd.t96 140.989
R1287 dvdd.t4 dvdd.t20 140.989
R1288 dvdd.t125 dvdd.t90 140.989
R1289 dvdd.t117 dvdd.t97 140.989
R1290 dvdd.t12 dvdd.t2 140.989
R1291 dvdd.t74 dvdd 132.597
R1292 dvdd dvdd.n272 125.883
R1293 dvdd dvdd.n271 125.883
R1294 dvdd dvdd.n270 125.883
R1295 dvdd.t79 dvdd.t68 121.245
R1296 dvdd.t77 dvdd.t79 121.245
R1297 dvdd.t167 dvdd.t77 121.245
R1298 dvdd.t42 dvdd.t167 121.245
R1299 dvdd.t55 dvdd.t171 121.245
R1300 dvdd.t40 dvdd.t55 121.245
R1301 dvdd.t70 dvdd.t40 121.245
R1302 dvdd.t169 dvdd.t70 121.245
R1303 dvdd.n71 dvdd.t155 119.608
R1304 dvdd.n72 dvdd.t118 119.608
R1305 dvdd.n92 dvdd.t121 119.608
R1306 dvdd.n93 dvdd.t154 119.608
R1307 dvdd.n113 dvdd.t85 119.608
R1308 dvdd.n114 dvdd.t143 119.608
R1309 dvdd.t93 dvdd 109.1
R1310 dvdd.t20 dvdd 109.1
R1311 dvdd.t2 dvdd 109.1
R1312 dvdd.n75 dvdd.t67 108.413
R1313 dvdd.n76 dvdd.t151 108.413
R1314 dvdd.n96 dvdd.t146 108.413
R1315 dvdd.n97 dvdd.t150 108.413
R1316 dvdd.n117 dvdd.t89 108.413
R1317 dvdd.n118 dvdd.t59 108.413
R1318 dvdd.n270 dvdd.n55 106.559
R1319 dvdd.n271 dvdd.n54 106.559
R1320 dvdd.n272 dvdd.n53 106.559
R1321 dvdd.n47 dvdd.n2 105.412
R1322 dvdd.n40 dvdd.n2 105.412
R1323 dvdd.n37 dvdd.n36 105.412
R1324 dvdd.n36 dvdd.n35 105.412
R1325 dvdd dvdd.t47 100.624
R1326 dvdd.n67 dvdd.t119 93.81
R1327 dvdd.n68 dvdd.t32 93.81
R1328 dvdd.n88 dvdd.t174 93.81
R1329 dvdd.n89 dvdd.t153 93.81
R1330 dvdd.n109 dvdd.t50 93.81
R1331 dvdd.n110 dvdd.t54 93.81
R1332 dvdd dvdd.t114 91.745
R1333 dvdd dvdd.t148 91.745
R1334 dvdd dvdd.t44 88.7855
R1335 dvdd.n258 dvdd.t48 86.7743
R1336 dvdd.n47 dvdd.n46 79.8123
R1337 dvdd.n41 dvdd.n40 79.8123
R1338 dvdd.n35 dvdd.n34 79.8123
R1339 dvdd.n37 dvdd.n26 79.8123
R1340 dvdd.n59 dvdd.t27 74.7554
R1341 dvdd.n238 dvdd.t139 74.7554
R1342 dvdd.n67 dvdd.t107 63.3219
R1343 dvdd.n68 dvdd.t122 63.3219
R1344 dvdd.n71 dvdd.t105 63.3219
R1345 dvdd.n72 dvdd.t91 63.3219
R1346 dvdd.n88 dvdd.t88 63.3219
R1347 dvdd.n89 dvdd.t17 63.3219
R1348 dvdd.n92 dvdd.t73 63.3219
R1349 dvdd.n93 dvdd.t123 63.3219
R1350 dvdd.n109 dvdd.t62 63.3219
R1351 dvdd.n110 dvdd.t104 63.3219
R1352 dvdd.n113 dvdd.t157 63.3219
R1353 dvdd.n114 dvdd.t103 63.3219
R1354 dvdd.n79 dvdd.t65 61.9829
R1355 dvdd.n100 dvdd.t163 61.9829
R1356 dvdd.n122 dvdd.t131 61.9829
R1357 dvdd.n80 dvdd.t156 61.9826
R1358 dvdd.n101 dvdd.t136 61.9826
R1359 dvdd.n123 dvdd.t101 61.9826
R1360 dvdd.n258 dvdd.t46 61.05
R1361 dvdd.n293 dvdd.t42 60.6225
R1362 dvdd.t171 dvdd.n293 60.6225
R1363 dvdd.n291 dvdd.t69 60.3236
R1364 dvdd.n295 dvdd.t170 60.3236
R1365 dvdd.n296 dvdd.n282 54.7085
R1366 dvdd.n297 dvdd.n281 54.7085
R1367 dvdd.n289 dvdd.n288 54.7085
R1368 dvdd.n290 dvdd.n287 54.7085
R1369 dvdd.n61 dvdd.t13 41.5552
R1370 dvdd.n61 dvdd.t3 41.5552
R1371 dvdd.n62 dvdd.t132 41.5552
R1372 dvdd.n62 dvdd.t30 41.5552
R1373 dvdd.n82 dvdd.t35 41.5552
R1374 dvdd.n82 dvdd.t21 41.5552
R1375 dvdd.n83 dvdd.t5 41.5552
R1376 dvdd.n83 dvdd.t60 41.5552
R1377 dvdd.n103 dvdd.t162 41.5552
R1378 dvdd.n103 dvdd.t94 41.5552
R1379 dvdd.n104 dvdd.t82 41.5552
R1380 dvdd.n104 dvdd.t173 41.5552
R1381 dvdd.n46 dvdd.n45 37.0005
R1382 dvdd.n42 dvdd.n41 37.0005
R1383 dvdd.n34 dvdd.n33 37.0005
R1384 dvdd.n30 dvdd.n26 37.0005
R1385 dvdd.n17 dvdd.t115 36.1587
R1386 dvdd.n17 dvdd.t128 36.1587
R1387 dvdd.n8 dvdd.t149 36.1587
R1388 dvdd.n8 dvdd.t109 36.1587
R1389 dvdd.n255 dvdd.t138 35.4605
R1390 dvdd.n249 dvdd.n248 34.6358
R1391 dvdd.n253 dvdd.n245 34.6358
R1392 dvdd.n264 dvdd.n256 34.6358
R1393 dvdd.n231 dvdd.n63 34.6358
R1394 dvdd.n221 dvdd.n65 34.6358
R1395 dvdd.n225 dvdd.n65 34.6358
R1396 dvdd.n226 dvdd.n225 34.6358
R1397 dvdd.n219 dvdd.n218 34.6358
R1398 dvdd.n213 dvdd.n212 34.6358
R1399 dvdd.n214 dvdd.n213 34.6358
R1400 dvdd.n200 dvdd.n199 34.6358
R1401 dvdd.n202 dvdd.n77 34.6358
R1402 dvdd.n206 dvdd.n77 34.6358
R1403 dvdd.n193 dvdd.n84 34.6358
R1404 dvdd.n183 dvdd.n86 34.6358
R1405 dvdd.n187 dvdd.n86 34.6358
R1406 dvdd.n188 dvdd.n187 34.6358
R1407 dvdd.n181 dvdd.n180 34.6358
R1408 dvdd.n175 dvdd.n174 34.6358
R1409 dvdd.n176 dvdd.n175 34.6358
R1410 dvdd.n162 dvdd.n161 34.6358
R1411 dvdd.n164 dvdd.n98 34.6358
R1412 dvdd.n168 dvdd.n98 34.6358
R1413 dvdd.n155 dvdd.n105 34.6358
R1414 dvdd.n145 dvdd.n107 34.6358
R1415 dvdd.n149 dvdd.n107 34.6358
R1416 dvdd.n150 dvdd.n149 34.6358
R1417 dvdd.n143 dvdd.n142 34.6358
R1418 dvdd.n137 dvdd.n136 34.6358
R1419 dvdd.n138 dvdd.n137 34.6358
R1420 dvdd.n124 dvdd.n52 34.6358
R1421 dvdd.n126 dvdd.n119 34.6358
R1422 dvdd.n130 dvdd.n119 34.6358
R1423 dvdd.n239 dvdd.n58 33.8829
R1424 dvdd.n227 dvdd.n226 32.377
R1425 dvdd.n189 dvdd.n188 32.377
R1426 dvdd.n151 dvdd.n150 32.377
R1427 dvdd.n214 dvdd.n69 32.0005
R1428 dvdd.n176 dvdd.n90 32.0005
R1429 dvdd.n138 dvdd.n111 32.0005
R1430 dvdd.n240 dvdd.n239 31.624
R1431 dvdd.n202 dvdd.n201 31.2476
R1432 dvdd.n164 dvdd.n163 31.2476
R1433 dvdd.n126 dvdd.n125 31.2476
R1434 dvdd.n5 dvdd.n3 30.8338
R1435 dvdd.n4 dvdd.n2 30.8338
R1436 dvdd.n36 dvdd.n27 30.8338
R1437 dvdd.n29 dvdd.n28 30.8338
R1438 dvdd.n79 dvdd.t134 30.1745
R1439 dvdd.n100 dvdd.t164 30.1745
R1440 dvdd.n122 dvdd.t53 30.1745
R1441 dvdd.n80 dvdd.t165 30.1738
R1442 dvdd.n101 dvdd.t130 30.1738
R1443 dvdd.n123 dvdd.t161 30.1738
R1444 dvdd.n208 dvdd.n73 30.1181
R1445 dvdd.n170 dvdd.n94 30.1181
R1446 dvdd.n132 dvdd.n115 30.1181
R1447 dvdd.n43 dvdd.n42 29.6618
R1448 dvdd.n45 dvdd.n44 29.6618
R1449 dvdd.n31 dvdd.n30 29.6618
R1450 dvdd.n33 dvdd.n32 29.6618
R1451 dvdd.n59 dvdd.t34 28.5349
R1452 dvdd.n238 dvdd.t160 28.5349
R1453 dvdd.n260 dvdd.n256 28.2952
R1454 dvdd dvdd.n245 27.8593
R1455 dvdd.n255 dvdd.t11 26.5955
R1456 dvdd.n259 dvdd.n257 25.2079
R1457 dvdd.n22 dvdd.n18 23.7181
R1458 dvdd.n11 dvdd.n10 23.7181
R1459 dvdd.n248 dvdd.n246 23.7181
R1460 dvdd.n233 dvdd.n55 23.7181
R1461 dvdd.n199 dvdd.n54 23.7181
R1462 dvdd.n195 dvdd.n54 23.7181
R1463 dvdd.n161 dvdd.n53 23.7181
R1464 dvdd.n157 dvdd.n53 23.7181
R1465 dvdd.n273 dvdd.n52 23.7181
R1466 dvdd.n58 dvdd.n55 23.7181
R1467 dvdd.n232 dvdd.n231 22.9652
R1468 dvdd.n194 dvdd.n193 22.9652
R1469 dvdd.n156 dvdd.n155 22.9652
R1470 dvdd.n266 dvdd.n254 22.5887
R1471 dvdd.n265 dvdd.n264 22.5887
R1472 dvdd.n266 dvdd.n265 21.8358
R1473 dvdd.n233 dvdd.n232 21.4593
R1474 dvdd.n195 dvdd.n194 21.4593
R1475 dvdd.n157 dvdd.n156 21.4593
R1476 dvdd.n212 dvdd.n73 20.3299
R1477 dvdd.n174 dvdd.n94 20.3299
R1478 dvdd.n136 dvdd.n115 20.3299
R1479 dvdd.n254 dvdd.n253 19.9534
R1480 dvdd.n240 dvdd.n56 19.577
R1481 dvdd.n269 dvdd.n56 18.4476
R1482 dvdd.n227 dvdd.n63 18.0711
R1483 dvdd.n189 dvdd.n84 18.0711
R1484 dvdd.n151 dvdd.n105 18.0711
R1485 dvdd.n23 dvdd 15.8123
R1486 dvdd dvdd.n9 15.8123
R1487 dvdd.n295 dvdd.n294 13.2148
R1488 dvdd.n292 dvdd.n291 13.2148
R1489 dvdd.n38 dvdd.n37 10.0436
R1490 dvdd.n35 dvdd.n1 9.59217
R1491 dvdd.n218 dvdd.n69 9.41227
R1492 dvdd.n180 dvdd.n90 9.41227
R1493 dvdd.n142 dvdd.n111 9.41227
R1494 dvdd.n19 dvdd.n18 9.3005
R1495 dvdd.n22 dvdd.n21 9.3005
R1496 dvdd.n10 dvdd.n6 9.3005
R1497 dvdd.n12 dvdd.n11 9.3005
R1498 dvdd.n40 dvdd.n39 9.3005
R1499 dvdd.n48 dvdd.n47 9.3005
R1500 dvdd.n261 dvdd.n260 9.3005
R1501 dvdd.n262 dvdd.n256 9.3005
R1502 dvdd.n264 dvdd.n263 9.3005
R1503 dvdd.n265 dvdd.n243 9.3005
R1504 dvdd.n254 dvdd.n244 9.3005
R1505 dvdd.n253 dvdd.n252 9.3005
R1506 dvdd.n251 dvdd.n245 9.3005
R1507 dvdd.n250 dvdd.n249 9.3005
R1508 dvdd.n248 dvdd.n247 9.3005
R1509 dvdd.n246 dvdd.n51 9.3005
R1510 dvdd.n269 dvdd.n268 9.3005
R1511 dvdd.n274 dvdd.n273 9.3005
R1512 dvdd.n120 dvdd.n52 9.3005
R1513 dvdd.n124 dvdd.n121 9.3005
R1514 dvdd.n127 dvdd.n126 9.3005
R1515 dvdd.n128 dvdd.n119 9.3005
R1516 dvdd.n130 dvdd.n129 9.3005
R1517 dvdd.n131 dvdd.n116 9.3005
R1518 dvdd.n133 dvdd.n132 9.3005
R1519 dvdd.n134 dvdd.n115 9.3005
R1520 dvdd.n136 dvdd.n135 9.3005
R1521 dvdd.n137 dvdd.n112 9.3005
R1522 dvdd.n139 dvdd.n138 9.3005
R1523 dvdd.n140 dvdd.n111 9.3005
R1524 dvdd.n142 dvdd.n141 9.3005
R1525 dvdd.n143 dvdd.n108 9.3005
R1526 dvdd.n146 dvdd.n145 9.3005
R1527 dvdd.n147 dvdd.n107 9.3005
R1528 dvdd.n149 dvdd.n148 9.3005
R1529 dvdd.n150 dvdd.n106 9.3005
R1530 dvdd.n152 dvdd.n151 9.3005
R1531 dvdd.n153 dvdd.n105 9.3005
R1532 dvdd.n155 dvdd.n154 9.3005
R1533 dvdd.n156 dvdd.n102 9.3005
R1534 dvdd.n158 dvdd.n157 9.3005
R1535 dvdd.n159 dvdd.n53 9.3005
R1536 dvdd.n161 dvdd.n160 9.3005
R1537 dvdd.n162 dvdd.n99 9.3005
R1538 dvdd.n165 dvdd.n164 9.3005
R1539 dvdd.n166 dvdd.n98 9.3005
R1540 dvdd.n168 dvdd.n167 9.3005
R1541 dvdd.n169 dvdd.n95 9.3005
R1542 dvdd.n171 dvdd.n170 9.3005
R1543 dvdd.n172 dvdd.n94 9.3005
R1544 dvdd.n174 dvdd.n173 9.3005
R1545 dvdd.n175 dvdd.n91 9.3005
R1546 dvdd.n177 dvdd.n176 9.3005
R1547 dvdd.n178 dvdd.n90 9.3005
R1548 dvdd.n180 dvdd.n179 9.3005
R1549 dvdd.n181 dvdd.n87 9.3005
R1550 dvdd.n184 dvdd.n183 9.3005
R1551 dvdd.n185 dvdd.n86 9.3005
R1552 dvdd.n187 dvdd.n186 9.3005
R1553 dvdd.n188 dvdd.n85 9.3005
R1554 dvdd.n190 dvdd.n189 9.3005
R1555 dvdd.n191 dvdd.n84 9.3005
R1556 dvdd.n193 dvdd.n192 9.3005
R1557 dvdd.n194 dvdd.n81 9.3005
R1558 dvdd.n196 dvdd.n195 9.3005
R1559 dvdd.n197 dvdd.n54 9.3005
R1560 dvdd.n199 dvdd.n198 9.3005
R1561 dvdd.n200 dvdd.n78 9.3005
R1562 dvdd.n203 dvdd.n202 9.3005
R1563 dvdd.n204 dvdd.n77 9.3005
R1564 dvdd.n206 dvdd.n205 9.3005
R1565 dvdd.n207 dvdd.n74 9.3005
R1566 dvdd.n209 dvdd.n208 9.3005
R1567 dvdd.n210 dvdd.n73 9.3005
R1568 dvdd.n212 dvdd.n211 9.3005
R1569 dvdd.n213 dvdd.n70 9.3005
R1570 dvdd.n215 dvdd.n214 9.3005
R1571 dvdd.n216 dvdd.n69 9.3005
R1572 dvdd.n218 dvdd.n217 9.3005
R1573 dvdd.n219 dvdd.n66 9.3005
R1574 dvdd.n222 dvdd.n221 9.3005
R1575 dvdd.n223 dvdd.n65 9.3005
R1576 dvdd.n225 dvdd.n224 9.3005
R1577 dvdd.n226 dvdd.n64 9.3005
R1578 dvdd.n228 dvdd.n227 9.3005
R1579 dvdd.n229 dvdd.n63 9.3005
R1580 dvdd.n231 dvdd.n230 9.3005
R1581 dvdd.n232 dvdd.n60 9.3005
R1582 dvdd.n234 dvdd.n233 9.3005
R1583 dvdd.n235 dvdd.n55 9.3005
R1584 dvdd.n236 dvdd.n58 9.3005
R1585 dvdd.n239 dvdd.n237 9.3005
R1586 dvdd.n239 dvdd.n57 9.3005
R1587 dvdd.n241 dvdd.n240 9.3005
R1588 dvdd.n242 dvdd.n56 9.3005
R1589 dvdd.n267 dvdd.n266 9.3005
R1590 dvdd.n208 dvdd.n207 9.03579
R1591 dvdd.n170 dvdd.n169 9.03579
R1592 dvdd.n132 dvdd.n131 9.03579
R1593 dvdd.n285 dvdd.n283 7.70883
R1594 dvdd.n293 dvdd.n285 7.70883
R1595 dvdd.n286 dvdd.n284 7.70883
R1596 dvdd.n293 dvdd.n286 7.70883
R1597 dvdd.n24 dvdd.n23 7.17001
R1598 dvdd.n9 dvdd.n7 7.15376
R1599 dvdd.n282 dvdd.t41 7.14175
R1600 dvdd.n282 dvdd.t71 7.14175
R1601 dvdd.n281 dvdd.t172 7.14175
R1602 dvdd.n281 dvdd.t56 7.14175
R1603 dvdd.n288 dvdd.t168 7.14175
R1604 dvdd.n288 dvdd.t43 7.14175
R1605 dvdd.n287 dvdd.t80 7.14175
R1606 dvdd.n287 dvdd.t78 7.14175
R1607 dvdd.n249 dvdd 6.77697
R1608 dvdd.n44 dvdd.t36 6.70818
R1609 dvdd.t36 dvdd.n43 6.70818
R1610 dvdd.n32 dvdd.t38 6.70818
R1611 dvdd.t38 dvdd.n31 6.70818
R1612 dvdd dvdd.n22 6.4005
R1613 dvdd.n10 dvdd 6.4005
R1614 dvdd.n221 dvdd.n220 6.02403
R1615 dvdd.n207 dvdd.n206 6.02403
R1616 dvdd.n183 dvdd.n182 6.02403
R1617 dvdd.n169 dvdd.n168 6.02403
R1618 dvdd.n145 dvdd.n144 6.02403
R1619 dvdd.n131 dvdd.n130 6.02403
R1620 dvdd.n220 dvdd.n219 3.76521
R1621 dvdd.n182 dvdd.n181 3.76521
R1622 dvdd.n144 dvdd.n143 3.76521
R1623 dvdd.n201 dvdd.n200 3.38874
R1624 dvdd.n163 dvdd.n162 3.38874
R1625 dvdd.n125 dvdd.n124 3.38874
R1626 dvdd.n296 dvdd.n295 1.66909
R1627 dvdd.n291 dvdd.n290 1.57188
R1628 dvdd.n36 dvdd.n0 1.32907
R1629 dvdd.n2 dvdd.n0 1.32907
R1630 dvdd.n260 dvdd.n259 1.23559
R1631 dvdd.n275 dvdd.n51 0.776793
R1632 dvdd.n275 dvdd.n274 0.637387
R1633 dvdd dvdd.n267 0.438
R1634 dvdd.n50 dvdd.n49 0.432317
R1635 dvdd.n16 dvdd 0.42713
R1636 dvdd dvdd.n16 0.32387
R1637 dvdd.n267 dvdd 0.313
R1638 dvdd.n7 dvdd 0.203706
R1639 dvdd.n13 dvdd 0.167167
R1640 dvdd.n19 dvdd 0.164848
R1641 dvdd.n257 dvdd 0.159538
R1642 dvdd.n38 dvdd.n15 0.141704
R1643 dvdd.n261 dvdd.n257 0.141672
R1644 dvdd.n38 dvdd.n25 0.139389
R1645 dvdd.n14 dvdd.n6 0.127236
R1646 dvdd.n263 dvdd.n243 0.120292
R1647 dvdd.n251 dvdd.n250 0.120292
R1648 dvdd.n252 dvdd.n251 0.120292
R1649 dvdd.n252 dvdd.n244 0.120292
R1650 dvdd.n121 dvdd.n120 0.120292
R1651 dvdd.n127 dvdd.n121 0.120292
R1652 dvdd.n128 dvdd.n127 0.120292
R1653 dvdd.n129 dvdd.n128 0.120292
R1654 dvdd.n129 dvdd.n116 0.120292
R1655 dvdd.n133 dvdd.n116 0.120292
R1656 dvdd.n134 dvdd.n133 0.120292
R1657 dvdd.n135 dvdd.n134 0.120292
R1658 dvdd.n135 dvdd.n112 0.120292
R1659 dvdd.n139 dvdd.n112 0.120292
R1660 dvdd.n140 dvdd.n139 0.120292
R1661 dvdd.n141 dvdd.n140 0.120292
R1662 dvdd.n141 dvdd.n108 0.120292
R1663 dvdd.n146 dvdd.n108 0.120292
R1664 dvdd.n147 dvdd.n146 0.120292
R1665 dvdd.n148 dvdd.n147 0.120292
R1666 dvdd.n148 dvdd.n106 0.120292
R1667 dvdd.n152 dvdd.n106 0.120292
R1668 dvdd.n153 dvdd.n152 0.120292
R1669 dvdd.n154 dvdd.n153 0.120292
R1670 dvdd.n154 dvdd.n102 0.120292
R1671 dvdd.n158 dvdd.n102 0.120292
R1672 dvdd.n160 dvdd.n99 0.120292
R1673 dvdd.n165 dvdd.n99 0.120292
R1674 dvdd.n166 dvdd.n165 0.120292
R1675 dvdd.n167 dvdd.n166 0.120292
R1676 dvdd.n167 dvdd.n95 0.120292
R1677 dvdd.n171 dvdd.n95 0.120292
R1678 dvdd.n172 dvdd.n171 0.120292
R1679 dvdd.n173 dvdd.n172 0.120292
R1680 dvdd.n173 dvdd.n91 0.120292
R1681 dvdd.n177 dvdd.n91 0.120292
R1682 dvdd.n178 dvdd.n177 0.120292
R1683 dvdd.n179 dvdd.n178 0.120292
R1684 dvdd.n179 dvdd.n87 0.120292
R1685 dvdd.n184 dvdd.n87 0.120292
R1686 dvdd.n185 dvdd.n184 0.120292
R1687 dvdd.n186 dvdd.n185 0.120292
R1688 dvdd.n186 dvdd.n85 0.120292
R1689 dvdd.n190 dvdd.n85 0.120292
R1690 dvdd.n191 dvdd.n190 0.120292
R1691 dvdd.n192 dvdd.n191 0.120292
R1692 dvdd.n192 dvdd.n81 0.120292
R1693 dvdd.n196 dvdd.n81 0.120292
R1694 dvdd.n198 dvdd.n78 0.120292
R1695 dvdd.n203 dvdd.n78 0.120292
R1696 dvdd.n204 dvdd.n203 0.120292
R1697 dvdd.n205 dvdd.n204 0.120292
R1698 dvdd.n205 dvdd.n74 0.120292
R1699 dvdd.n209 dvdd.n74 0.120292
R1700 dvdd.n210 dvdd.n209 0.120292
R1701 dvdd.n211 dvdd.n210 0.120292
R1702 dvdd.n211 dvdd.n70 0.120292
R1703 dvdd.n215 dvdd.n70 0.120292
R1704 dvdd.n216 dvdd.n215 0.120292
R1705 dvdd.n217 dvdd.n216 0.120292
R1706 dvdd.n217 dvdd.n66 0.120292
R1707 dvdd.n222 dvdd.n66 0.120292
R1708 dvdd.n223 dvdd.n222 0.120292
R1709 dvdd.n224 dvdd.n223 0.120292
R1710 dvdd.n224 dvdd.n64 0.120292
R1711 dvdd.n228 dvdd.n64 0.120292
R1712 dvdd.n229 dvdd.n228 0.120292
R1713 dvdd.n230 dvdd.n229 0.120292
R1714 dvdd.n230 dvdd.n60 0.120292
R1715 dvdd.n234 dvdd.n60 0.120292
R1716 dvdd.n237 dvdd.n236 0.120292
R1717 dvdd.n241 dvdd.n57 0.120292
R1718 dvdd.n242 dvdd.n241 0.120292
R1719 dvdd.n276 dvdd.n275 0.109494
R1720 dvdd.n15 dvdd.n14 0.109053
R1721 dvdd.n267 dvdd.n244 0.107271
R1722 dvdd.n14 dvdd 0.0983618
R1723 dvdd dvdd.n261 0.0981562
R1724 dvdd.n250 dvdd 0.0968542
R1725 dvdd.n280 dvdd.n279 0.0944312
R1726 dvdd.n277 dvdd.n276 0.0856755
R1727 dvdd.n278 dvdd.n277 0.0856755
R1728 dvdd.n237 dvdd 0.0812292
R1729 dvdd dvdd.n6 0.0803611
R1730 dvdd.n279 dvdd.n278 0.0777774
R1731 dvdd.n14 dvdd.n7 0.070241
R1732 dvdd.n25 dvdd.n24 0.0685285
R1733 dvdd.n267 dvdd 0.063
R1734 dvdd.n263 dvdd 0.0603958
R1735 dvdd dvdd.n262 0.0603958
R1736 dvdd.n247 dvdd 0.0603958
R1737 dvdd.n120 dvdd 0.0603958
R1738 dvdd.n159 dvdd 0.0603958
R1739 dvdd.n160 dvdd 0.0603958
R1740 dvdd.n197 dvdd 0.0603958
R1741 dvdd.n198 dvdd 0.0603958
R1742 dvdd.n235 dvdd 0.0603958
R1743 dvdd.n236 dvdd 0.0603958
R1744 dvdd.n268 dvdd 0.0603958
R1745 dvdd dvdd.n13 0.0595278
R1746 dvdd.n21 dvdd.n16 0.0535523
R1747 dvdd.n12 dvdd 0.0508472
R1748 dvdd.n290 dvdd.n289 0.0456945
R1749 dvdd.n39 dvdd.n38 0.0456858
R1750 dvdd.n20 dvdd 0.0405
R1751 dvdd dvdd.n57 0.0395625
R1752 dvdd dvdd.n296 0.0385435
R1753 dvdd dvdd.n51 0.0382604
R1754 dvdd.n39 dvdd.n0 0.0379437
R1755 dvdd.n21 dvdd 0.0339302
R1756 dvdd.n13 dvdd.n12 0.0334861
R1757 dvdd.n274 dvdd 0.03175
R1758 dvdd dvdd.n159 0.03175
R1759 dvdd dvdd.n197 0.03175
R1760 dvdd dvdd.n235 0.03175
R1761 dvdd.n268 dvdd 0.03175
R1762 dvdd.n24 dvdd.n16 0.0300191
R1763 dvdd.n247 dvdd 0.0239375
R1764 dvdd.n49 dvdd.n0 0.0233041
R1765 dvdd.n262 dvdd 0.0226354
R1766 dvdd dvdd.n158 0.0226354
R1767 dvdd dvdd.n196 0.0226354
R1768 dvdd dvdd.n234 0.0226354
R1769 dvdd dvdd.n242 0.0226354
R1770 dvdd.n298 dvdd.n297 0.0219531
R1771 dvdd.n15 dvdd 0.0210592
R1772 dvdd.n20 dvdd.n19 0.0205
R1773 dvdd.n48 dvdd.n1 0.0182365
R1774 dvdd.n25 dvdd 0.0179419
R1775 dvdd.n49 dvdd.n48 0.0151396
R1776 dvdd.n289 dvdd.n280 0.0150881
R1777 dvdd dvdd.n20 0.0121279
R1778 dvdd.n298 dvdd.n280 0.00936728
R1779 dvdd.n267 dvdd.n243 0.0083125
R1780 dvdd.n276 dvdd.t178 0.0083125
R1781 dvdd.n277 dvdd.t177 0.0083125
R1782 dvdd.n278 dvdd.t176 0.0083125
R1783 dvdd.n50 dvdd.t175 0.0083125
R1784 dvdd.n297 dvdd 0.00765103
R1785 dvdd.n279 dvdd.n50 0.00754239
R1786 dvdd.n1 dvdd 0.00176689
R1787 dvdd.n298 dvdd 0.001125
R1788 a_20376_n2791.n1 a_20376_n2791.n0 926.024
R1789 a_20376_n2791.n1 a_20376_n2791.t3 82.0838
R1790 a_20376_n2791.n0 a_20376_n2791.t0 63.3338
R1791 a_20376_n2791.t1 a_20376_n2791.n1 63.3219
R1792 a_20376_n2791.n0 a_20376_n2791.t2 29.7268
R1793 a_19955_n2241.n1 a_19955_n2241.t7 530.01
R1794 a_19955_n2241.t0 a_19955_n2241.n5 421.021
R1795 a_19955_n2241.n0 a_19955_n2241.t2 337.142
R1796 a_19955_n2241.n3 a_19955_n2241.t1 280.223
R1797 a_19955_n2241.n4 a_19955_n2241.t3 263.173
R1798 a_19955_n2241.n4 a_19955_n2241.t5 227.826
R1799 a_19955_n2241.n0 a_19955_n2241.t4 199.762
R1800 a_19955_n2241.n2 a_19955_n2241.n1 170.81
R1801 a_19955_n2241.n2 a_19955_n2241.n0 167.321
R1802 a_19955_n2241.n5 a_19955_n2241.n4 152
R1803 a_19955_n2241.n1 a_19955_n2241.t6 141.923
R1804 a_19955_n2241.n3 a_19955_n2241.n2 10.8376
R1805 a_19955_n2241.n5 a_19955_n2241.n3 2.50485
R1806 a_20689_n2273.n3 a_20689_n2273.n2 647.119
R1807 a_20689_n2273.n1 a_20689_n2273.t4 350.253
R1808 a_20689_n2273.n2 a_20689_n2273.n0 260.339
R1809 a_20689_n2273.n2 a_20689_n2273.n1 246.119
R1810 a_20689_n2273.n1 a_20689_n2273.t5 189.588
R1811 a_20689_n2273.n3 a_20689_n2273.t2 89.1195
R1812 a_20689_n2273.n0 a_20689_n2273.t1 63.3338
R1813 a_20689_n2273.t0 a_20689_n2273.n3 41.0422
R1814 a_20689_n2273.n0 a_20689_n2273.t3 31.9797
R1815 a_21036_n1869.n3 a_21036_n1869.n2 636.953
R1816 a_21036_n1869.n1 a_21036_n1869.t5 366.856
R1817 a_21036_n1869.n2 a_21036_n1869.n0 300.2
R1818 a_21036_n1869.n2 a_21036_n1869.n1 225.036
R1819 a_21036_n1869.n1 a_21036_n1869.t4 174.056
R1820 a_21036_n1869.n0 a_21036_n1869.t0 70.0005
R1821 a_21036_n1869.n3 a_21036_n1869.t3 68.0124
R1822 a_21036_n1869.t1 a_21036_n1869.n3 63.3219
R1823 a_21036_n1869.n0 a_21036_n1869.t2 61.6672
R1824 a_10620_n8338.t0 a_10620_n8338.t1 83.9243
R1825 a_24220_n8172.t0 a_24220_n8172.t1 83.56
R1826 a_16620_n2791.n3 a_16620_n2791.n2 636.953
R1827 a_16620_n2791.n1 a_16620_n2791.t4 366.856
R1828 a_16620_n2791.n2 a_16620_n2791.n0 300.2
R1829 a_16620_n2791.n2 a_16620_n2791.n1 225.036
R1830 a_16620_n2791.n1 a_16620_n2791.t5 174.056
R1831 a_16620_n2791.n0 a_16620_n2791.t0 70.0005
R1832 a_16620_n2791.t1 a_16620_n2791.n3 68.0124
R1833 a_16620_n2791.n3 a_16620_n2791.t3 63.3219
R1834 a_16620_n2791.n0 a_16620_n2791.t2 61.6672
R1835 a_16974_n2791.t0 a_16974_n2791.t1 87.1434
R1836 a_16795_n2817.n6 a_16795_n2817.n5 746.659
R1837 a_16795_n2817.n0 a_16795_n2817.t3 389.183
R1838 a_16795_n2817.n2 a_16795_n2817.t7 256.988
R1839 a_16795_n2817.n1 a_16795_n2817.n0 251.167
R1840 a_16795_n2817.n1 a_16795_n2817.t1 223.571
R1841 a_16795_n2817.n4 a_16795_n2817.t5 212.081
R1842 a_16795_n2817.n5 a_16795_n2817.n4 181.942
R1843 a_16795_n2817.n0 a_16795_n2817.t8 174.891
R1844 a_16795_n2817.n2 a_16795_n2817.t4 163.803
R1845 a_16795_n2817.n3 a_16795_n2817.t6 139.78
R1846 a_16795_n2817.n3 a_16795_n2817.n2 129.264
R1847 a_16795_n2817.n6 a_16795_n2817.t2 63.3219
R1848 a_16795_n2817.t0 a_16795_n2817.n6 63.3219
R1849 a_16795_n2817.n5 a_16795_n2817.n1 24.6993
R1850 a_16795_n2817.n4 a_16795_n2817.n3 22.6399
R1851 ena_ip.t0 ena_ip.n0 744.115
R1852 ena_ip ena_ip.t0 732.75
R1853 ena_ip.n15 ena_ip.t7 408.63
R1854 ena_ip.n11 ena_ip.t13 408.63
R1855 ena_ip.n7 ena_ip.t4 408.63
R1856 ena_ip.n12 ena_ip.t6 347.577
R1857 ena_ip.n8 ena_ip.t8 347.577
R1858 ena_ip.n4 ena_ip.t16 347.577
R1859 ena_ip.n2 ena_ip.t14 332.752
R1860 ena_ip.t14 ena_ip.n1 332.752
R1861 ena_ip.n2 ena_ip.t17 332.411
R1862 ena_ip.t17 ena_ip.n1 332.411
R1863 ena_ip.n16 ena_ip.t19 239.505
R1864 ena_ip ena_ip.t1 216.155
R1865 ena_ip.n12 ena_ip.t9 193.337
R1866 ena_ip.n8 ena_ip.t10 193.337
R1867 ena_ip.n4 ena_ip.t18 193.337
R1868 ena_ip.n16 ena_ip.t11 167.204
R1869 ena_ip ena_ip.n15 165.089
R1870 ena_ip ena_ip.n11 165.089
R1871 ena_ip ena_ip.n7 165.089
R1872 ena_ip ena_ip.n16 157.12
R1873 ena_ip.n13 ena_ip.n12 152
R1874 ena_ip.n9 ena_ip.n8 152
R1875 ena_ip.n5 ena_ip.n4 152
R1876 ena_ip.n15 ena_ip.t3 132.282
R1877 ena_ip.n11 ena_ip.t5 132.282
R1878 ena_ip.n7 ena_ip.t15 132.282
R1879 ena_ip ena_ip.t2 59.9857
R1880 ena_ip ena_ip.t12 59.0936
R1881 ena_ip.n0 ena_ip 57.4755
R1882 ena_ip ena_ip.n17 13.8078
R1883 ena_ip.n17 ena_ip 9.82907
R1884 ena_ip ena_ip.n6 9.3005
R1885 ena_ip ena_ip.n10 9.3005
R1886 ena_ip ena_ip.n14 9.3005
R1887 ena_ip ena_ip.n18 8.84514
R1888 ena_ip.n17 ena_ip 5.71479
R1889 ena_ip.n3 ena_ip.n1 5.53161
R1890 ena_ip.n13 ena_ip 4.67077
R1891 ena_ip.n9 ena_ip 4.67077
R1892 ena_ip.n5 ena_ip 4.67077
R1893 ena_ip.n3 ena_ip.n2 4.67076
R1894 ena_ip.n18 ena_ip 4.17561
R1895 ena_ip.n0 ena_ip 3.62625
R1896 ena_ip ena_ip.n3 3.51723
R1897 ena_ip.n14 ena_ip 2.94104
R1898 ena_ip.n10 ena_ip 2.94104
R1899 ena_ip.n6 ena_ip 2.94104
R1900 ena_ip.n18 ena_ip 2.93705
R1901 ena_ip.n14 ena_ip.n13 2.76807
R1902 ena_ip.n10 ena_ip.n9 2.76807
R1903 ena_ip.n6 ena_ip.n5 2.76807
R1904 x3.in_b.n1 x3.in_b.n0 3.2348
R1905 x3.in_b.n1 x3.in_b.t3 166.376
R1906 x3.in_b.n1 x3.in_b.t2 166.207
R1907 x3.in_b.n0 x3.in_b.t0 228.429
R1908 x3.in_b.n0 x3.in_b.t1 83.9309
R1909 a_21211_n1943.n6 a_21211_n1943.n5 746.659
R1910 a_21211_n1943.n0 a_21211_n1943.t6 389.183
R1911 a_21211_n1943.n2 a_21211_n1943.t4 256.988
R1912 a_21211_n1943.n1 a_21211_n1943.n0 251.167
R1913 a_21211_n1943.n1 a_21211_n1943.t1 223.571
R1914 a_21211_n1943.n4 a_21211_n1943.t7 212.081
R1915 a_21211_n1943.n5 a_21211_n1943.n4 181.942
R1916 a_21211_n1943.n0 a_21211_n1943.t8 174.891
R1917 a_21211_n1943.n2 a_21211_n1943.t5 163.803
R1918 a_21211_n1943.n3 a_21211_n1943.t3 139.78
R1919 a_21211_n1943.n3 a_21211_n1943.n2 129.264
R1920 a_21211_n1943.n6 a_21211_n1943.t2 63.3219
R1921 a_21211_n1943.t0 a_21211_n1943.n6 63.3219
R1922 a_21211_n1943.n5 a_21211_n1943.n1 24.6993
R1923 a_21211_n1943.n4 a_21211_n1943.n3 22.6399
R1924 a_17913_n2791.t0 a_17913_n2791.n3 370.026
R1925 a_17913_n2791.n0 a_17913_n2791.t2 351.356
R1926 a_17913_n2791.n1 a_17913_n2791.t5 334.717
R1927 a_17913_n2791.n3 a_17913_n2791.t1 325.971
R1928 a_17913_n2791.n1 a_17913_n2791.t4 309.935
R1929 a_17913_n2791.n0 a_17913_n2791.t3 305.683
R1930 a_17913_n2791.n2 a_17913_n2791.n0 16.879
R1931 a_17913_n2791.n3 a_17913_n2791.n2 10.8867
R1932 a_17913_n2791.n2 a_17913_n2791.n1 9.3005
R1933 a_18481_n2549.n3 a_18481_n2549.n2 647.119
R1934 a_18481_n2549.n1 a_18481_n2549.t4 350.253
R1935 a_18481_n2549.n2 a_18481_n2549.n0 260.339
R1936 a_18481_n2549.n2 a_18481_n2549.n1 246.119
R1937 a_18481_n2549.n1 a_18481_n2549.t5 189.588
R1938 a_18481_n2549.n3 a_18481_n2549.t2 89.1195
R1939 a_18481_n2549.n0 a_18481_n2549.t3 63.3338
R1940 a_18481_n2549.t0 a_18481_n2549.n3 41.0422
R1941 a_18481_n2549.n0 a_18481_n2549.t1 31.9797
R1942 a_18828_n2791.n3 a_18828_n2791.n2 636.953
R1943 a_18828_n2791.n1 a_18828_n2791.t4 366.856
R1944 a_18828_n2791.n2 a_18828_n2791.n0 300.2
R1945 a_18828_n2791.n2 a_18828_n2791.n1 225.036
R1946 a_18828_n2791.n1 a_18828_n2791.t5 174.056
R1947 a_18828_n2791.n0 a_18828_n2791.t2 70.0005
R1948 a_18828_n2791.t1 a_18828_n2791.n3 68.0124
R1949 a_18828_n2791.n3 a_18828_n2791.t3 63.3219
R1950 a_18828_n2791.n0 a_18828_n2791.t0 61.6672
R1951 a_2130_n19848.t0 a_2130_n19848.t1 82.0028
R1952 a_24530_n20014.t0 a_24530_n20014.t1 81.9478
R1953 icnode.t1 icnode.t0 84.1171
R1954 a_11526_n12394.t0 a_11526_n12394.t1 78.7148
R1955 vbreg.n21 vbreg.t2 244.944
R1956 vbreg.n49 vbreg.n2 202.542
R1957 vbreg.n40 vbreg.n10 201.036
R1958 vbreg.n33 vbreg.n7 200.282
R1959 vbreg.n20 vbreg.n21 0.962138
R1960 vbreg.n35 vbreg.n10 179.201
R1961 vbreg.n2 vbreg.n24 178.447
R1962 vbreg.n35 vbreg.n7 176.941
R1963 vbreg.n42 vbreg.n24 160.376
R1964 vbreg.n35 vbreg.n19 116.609
R1965 vbreg.n35 vbreg.n15 116.609
R1966 vbreg.n30 vbreg.n10 116.609
R1967 vbreg.n17 vbreg.n10 116.609
R1968 vbreg.n44 vbreg.n24 116.609
R1969 vbreg.n56 vbreg.n24 116.609
R1970 vbreg.n53 vbreg.n2 116.609
R1971 vbreg.n2 vbreg.n25 116.609
R1972 vbreg.n18 vbreg.n7 116.609
R1973 vbreg.n16 vbreg.n7 116.609
R1974 vbreg.n42 vbreg.n26 115.005
R1975 vbreg.n42 vbreg.n40 110.683
R1976 vbreg.t13 vbreg.n31 86.3125
R1977 vbreg.n14 vbreg.t10 88.4838
R1978 vbreg.n18 vbreg.t14 86.3125
R1979 vbreg.t12 vbreg.n16 86.3125
R1980 vbreg.t23 vbreg.n12 88.4979
R1981 vbreg.n51 vbreg.t25 86.3125
R1982 vbreg.t17 vbreg.n38 86.3125
R1983 vbreg.n28 vbreg.t18 86.3125
R1984 vbreg.n15 vbreg.t9 86.3125
R1985 vbreg.n19 vbreg.t11 86.3125
R1986 vbreg.n37 vbreg.t15 86.3125
R1987 vbreg.n29 vbreg.t16 86.3125
R1988 vbreg.n57 vbreg.t7 86.3125
R1989 vbreg.n43 vbreg.t20 86.3125
R1990 vbreg.n55 vbreg.t19 86.3125
R1991 vbreg.n54 vbreg.t22 86.3125
R1992 vbreg.n47 vbreg.t21 86.3125
R1993 vbreg.n52 vbreg.t24 86.3125
R1994 vbreg.n16 vbreg.n14 2.64048
R1995 vbreg.n38 vbreg.n37 72.5338
R1996 vbreg.n12 vbreg.n47 2.18593
R1997 vbreg.n18 vbreg.n31 72.5338
R1998 vbreg.n29 vbreg.n28 72.5338
R1999 vbreg.n52 vbreg.n51 72.5338
R2000 vbreg.n15 vbreg.n17 71.7809
R2001 vbreg.n57 vbreg.n56 71.7809
R2002 vbreg.n19 vbreg.n30 71.7809
R2003 vbreg.n28 vbreg.n26 71.7809
R2004 vbreg.n44 vbreg.n43 71.7809
R2005 vbreg.n16 vbreg.n15 71.5299
R2006 vbreg.n13 vbreg.n18 2.62088
R2007 vbreg.n55 vbreg.n25 71.2789
R2008 vbreg.n54 vbreg.n53 71.2789
R2009 vbreg.n38 vbreg.n23 60.7378
R2010 vbreg.n11 vbreg.t8 60.1061
R2011 vbreg.n32 vbreg.t13 55.9125
R2012 vbreg.n32 vbreg.t10 55.9125
R2013 vbreg.t14 vbreg.n34 55.9125
R2014 vbreg.n34 vbreg.t12 55.9125
R2015 vbreg.n48 vbreg.t23 55.9125
R2016 vbreg.n48 vbreg.t25 55.9125
R2017 vbreg.n39 vbreg.t17 55.9125
R2018 vbreg.n39 vbreg.t18 55.9125
R2019 vbreg.t9 vbreg.n36 55.9125
R2020 vbreg.n36 vbreg.t11 55.9125
R2021 vbreg.n27 vbreg.t15 55.9125
R2022 vbreg.t16 vbreg.n27 55.9125
R2023 vbreg.n41 vbreg.t7 55.9125
R2024 vbreg.n41 vbreg.t20 55.9125
R2025 vbreg.n45 vbreg.t19 55.9125
R2026 vbreg.t22 vbreg.n45 55.9125
R2027 vbreg.t21 vbreg.n46 55.9125
R2028 vbreg.n46 vbreg.t24 55.9125
R2029 vbreg.n33 vbreg.n32 30.4005
R2030 vbreg.n49 vbreg.n48 30.4005
R2031 vbreg.n36 vbreg.n35 30.4005
R2032 vbreg.n27 vbreg.n10 30.4005
R2033 vbreg.n40 vbreg.n39 30.4005
R2034 vbreg.n42 vbreg.n41 30.4005
R2035 vbreg.n45 vbreg.n24 30.4005
R2036 vbreg.n46 vbreg.n2 30.4005
R2037 vbreg.n34 vbreg.n7 30.4005
R2038 vbreg.n21 vbreg.t1 22.4019
R2039 vbreg.n22 vbreg.t3 21.1527
R2040 vbreg.n21 vbreg.t0 21.0621
R2041 vbreg.n42 vbreg.n11 2.00645
R2042 vbreg.n11 vbreg.n23 15.0573
R2043 vbreg.n57 vbreg.n23 11.7966
R2044 vbreg.n21 vbreg.n22 0.632464
R2045 vbreg.n40 vbreg.n3 3.01598
R2046 vbreg.n51 vbreg.n50 2.92951
R2047 vbreg.n4 vbreg.n31 2.92951
R2048 vbreg.n50 vbreg.n49 2.3255
R2049 vbreg.n0 vbreg.n2 2.3255
R2050 vbreg.n38 vbreg.n3 2.3255
R2051 vbreg.n55 vbreg.n3 2.3255
R2052 vbreg.n0 vbreg.n54 2.3255
R2053 vbreg.n52 vbreg.n0 2.3255
R2054 vbreg.n4 vbreg.n33 2.3255
R2055 vbreg.n5 vbreg.n7 2.3255
R2056 vbreg.n37 vbreg.n9 2.3255
R2057 vbreg.n9 vbreg.n10 2.3255
R2058 vbreg.n29 vbreg.n9 2.3255
R2059 vbreg.n28 vbreg.n8 2.3255
R2060 vbreg.n43 vbreg.n8 2.3255
R2061 vbreg.n3 vbreg.n57 2.3255
R2062 vbreg.n8 vbreg.n11 1.77359
R2063 vbreg.n3 vbreg.n20 1.69825
R2064 vbreg.n47 vbreg.n25 1.2554
R2065 vbreg.n53 vbreg.n52 1.2554
R2066 vbreg.n20 vbreg.t4 21.8362
R2067 vbreg.n21 vbreg.t6 21.6418
R2068 vbreg.n22 vbreg.t5 21.6076
R2069 vbreg.n19 vbreg.n13 2.62088
R2070 vbreg.n9 vbreg.n15 2.82746
R2071 vbreg.n6 vbreg.n5 0.489702
R2072 vbreg.n9 vbreg.n6 0.553315
R2073 vbreg.n1 vbreg.n0 0.420519
R2074 vbreg.n9 vbreg.n8 1.22324
R2075 vbreg.n6 vbreg.n35 2.715
R2076 vbreg.n12 vbreg.n0 1.45199
R2077 vbreg.n50 vbreg.n0 1.13148
R2078 vbreg.n5 vbreg.n4 1.12454
R2079 vbreg.n1 vbreg.n3 0.237615
R2080 vbreg.n5 vbreg.n13 0.795018
R2081 vbreg.n14 vbreg.n5 0.776083
R2082 vbreg.n3 vbreg.n11 0.753999
R2083 vbreg.n37 vbreg.n17 0.753441
R2084 vbreg.n56 vbreg.n55 0.753441
R2085 vbreg.n30 vbreg.n29 0.753441
R2086 vbreg.n43 vbreg.n26 0.753441
R2087 vbreg.n54 vbreg.n44 0.753441
R2088 vbreg.n1 vbreg.n24 2.61619
R2089 a_15000_n2791.n2 a_15000_n2791.n1 682.193
R2090 a_15000_n2791.n0 a_15000_n2791.t4 279.142
R2091 a_15000_n2791.n1 a_15000_n2791.t2 250.526
R2092 a_15000_n2791.n0 a_15000_n2791.t3 145.958
R2093 a_15000_n2791.n1 a_15000_n2791.n0 118.642
R2094 a_15000_n2791.t0 a_15000_n2791.n2 70.3576
R2095 a_15000_n2791.n2 a_15000_n2791.t1 65.6672
R2096 x7.x2.x2.CLK x7.x2.x2.CLK.t0 721.571
R2097 x7.x2.x2.CLK.n2 x7.x2.x2.CLK.t0 707.66
R2098 x7.x2.x2.CLK.n0 x7.x2.x2.CLK.t2 294.557
R2099 x7.x2.x2.CLK.n1 x7.x2.x2.CLK.t1 271.777
R2100 x7.x2.x2.CLK.n0 x7.x2.x2.CLK.t3 211.01
R2101 x7.x2.x2.CLK x7.x2.x2.CLK.n0 152
R2102 x7.x2.x2.CLK.n2 x7.x2.x2.CLK.n1 38.2982
R2103 x7.x2.x2.CLK.n1 x7.x2.x2.CLK 32.5125
R2104 x7.x2.x2.CLK x7.x2.x2.CLK.n2 3.76521
R2105 x7.x1.Qb2.n4 x7.x1.Qb2.t1 372.361
R2106 x7.x1.Qb2.n2 x7.x1.Qb2.t2 333.651
R2107 x7.x1.Qb2.n2 x7.x1.Qb2.t5 297.233
R2108 x7.x1.Qb2.n0 x7.x1.Qb2.t3 294.557
R2109 x7.x1.Qb2.n5 x7.x1.Qb2.t0 231.921
R2110 x7.x1.Qb2.n0 x7.x1.Qb2.t4 211.01
R2111 x7.x1.Qb2 x7.x1.Qb2.n2 195.701
R2112 x7.x1.Qb2.n1 x7.x1.Qb2.n0 152
R2113 x7.x1.Qb2.n5 x7.x1.Qb2.n1 41.5091
R2114 x7.x1.Qb2.n5 x7.x1.Qb2.n4 18.1966
R2115 x7.x1.Qb2.n4 x7.x1.Qb2.n3 9.36092
R2116 x7.x1.Qb2.n3 x7.x1.Qb2 6.49269
R2117 x7.x1.Qb2.n1 x7.x1.Qb2 4.20621
R2118 x7.x1.Qb2.n3 x7.x1.Qb2 3.52967
R2119 x7.x1.Qb2 x7.x1.Qb2.n5 2.5605
R2120 a_18168_n1881.n1 a_18168_n1881.n0 926.024
R2121 a_18168_n1881.n1 a_18168_n1881.t2 82.0838
R2122 a_18168_n1881.n0 a_18168_n1881.t3 63.3338
R2123 a_18168_n1881.t0 a_18168_n1881.n1 63.3219
R2124 a_18168_n1881.n0 a_18168_n1881.t1 29.7268
R2125 vbp.n3 vbp.n4 26.3414
R2126 vbp.n0 vbp 26.2397
R2127 vbp vbp.t2 112.21
R2128 vbp.n5 vbp.t12 21.3971
R2129 vbp.t10 vbp.n7 21.2714
R2130 vbp.n1 vbp.t13 21.3971
R2131 vbp.n3 vbp.n6 8.08368
R2132 vbp.n3 vbp.n5 8.21681
R2133 vbp.t17 vbp.n4 16.1817
R2134 vbp vbp.n2 8.77241
R2135 vbp vbp.t0 40.0025
R2136 vbp.t6 vbp 21.3013
R2137 vbp vbp.t16 21.3065
R2138 vbp.t3 vbp.n7 21.3313
R2139 vbp.n6 vbp.t14 21.0504
R2140 vbp.t4 vbp.n6 21.0498
R2141 vbp.n5 vbp.t7 20.9537
R2142 vbp.t11 vbp.n4 33.1891
R2143 vbp.t1 vbp.n2 21.7234
R2144 vbp.t9 vbp.n2 21.1857
R2145 vbp.t8 vbp.n1 20.9537
R2146 vbp.n0 vbp.t15 33.1158
R2147 vbp.n7 vbp 17.5035
R2148 vbp.n3 vbp 12.5283
R2149 vbp.n0 vbp.t5 16.2176
R2150 vbp vbp.n1 13.871
R2151 dvdd_ip.n100 dvdd_ip.n43 36575
R2152 dvdd_ip.n101 dvdd_ip.n100 36575
R2153 dvdd_ip.n102 dvdd_ip.n43 36575
R2154 dvdd_ip.n102 dvdd_ip.n101 36575
R2155 dvdd_ip.n99 dvdd_ip.n41 18251.4
R2156 dvdd_ip.n99 dvdd_ip.n42 18251.4
R2157 dvdd_ip.n103 dvdd_ip.n41 18251.4
R2158 dvdd_ip.n103 dvdd_ip.n42 18251.4
R2159 dvdd_ip.n79 dvdd_ip.n57 10440
R2160 dvdd_ip.n81 dvdd_ip.n57 10440
R2161 dvdd_ip.n81 dvdd_ip.n58 10440
R2162 dvdd_ip.n79 dvdd_ip.n58 10440
R2163 dvdd_ip.n105 dvdd_ip.n104 4516.33
R2164 dvdd_ip.n104 dvdd_ip.n40 4243.24
R2165 dvdd_ip.n38 dvdd_ip.n32 4030.59
R2166 dvdd_ip.n36 dvdd_ip.n35 4030.59
R2167 dvdd_ip.n65 dvdd_ip.n64 4030.59
R2168 dvdd_ip.n62 dvdd_ip.n61 4030.59
R2169 dvdd_ip.n98 dvdd_ip.n5 3741.35
R2170 dvdd_ip.n98 dvdd_ip.n97 3618.82
R2171 dvdd_ip.n74 dvdd_ip.n70 3190.03
R2172 dvdd_ip.n74 dvdd_ip.n71 3190.03
R2173 dvdd_ip.n72 dvdd_ip.n71 3190.03
R2174 dvdd_ip.n72 dvdd_ip.n70 3190.03
R2175 dvdd_ip.n96 dvdd_ip.n95 2795.29
R2176 dvdd_ip.n93 dvdd_ip.n45 2795.29
R2177 dvdd_ip.n90 dvdd_ip.n46 2417.65
R2178 dvdd_ip.n90 dvdd_ip.n47 2417.65
R2179 dvdd_ip.n92 dvdd_ip.n47 2417.65
R2180 dvdd_ip.n92 dvdd_ip.n46 2417.65
R2181 dvdd_ip.n65 dvdd_ip.n60 1199.77
R2182 dvdd_ip.n63 dvdd_ip.n62 1199.77
R2183 dvdd_ip.n96 dvdd_ip.n44 703.912
R2184 dvdd_ip.n94 dvdd_ip.n93 703.912
R2185 dvdd_ip.n105 dvdd_ip.n39 654.165
R2186 dvdd_ip.n56 dvdd_ip.t17 642.13
R2187 dvdd_ip.n88 dvdd_ip.t14 642.13
R2188 dvdd_ip.n29 dvdd_ip.t1 642.13
R2189 dvdd_ip.n11 dvdd_ip.n83 594.953
R2190 dvdd_ip.n11 dvdd_ip.n84 594.301
R2191 dvdd_ip.n39 dvdd_ip.n31 429.93
R2192 dvdd_ip.n33 dvdd_ip.n31 429.93
R2193 dvdd_ip.t40 dvdd_ip.t24 397.805
R2194 dvdd_ip.t32 dvdd_ip.t40 397.805
R2195 dvdd_ip.t34 dvdd_ip.t32 397.805
R2196 dvdd_ip.t27 dvdd_ip.t42 397.805
R2197 dvdd_ip.t38 dvdd_ip.t27 397.805
R2198 dvdd_ip.t29 dvdd_ip.t38 397.805
R2199 dvdd_ip.n33 dvdd_ip.n30 340.42
R2200 dvdd_ip.n92 dvdd_ip.t9 327.8
R2201 dvdd_ip.t7 dvdd_ip.n90 327.8
R2202 dvdd_ip.t19 dvdd_ip.t23 312.123
R2203 dvdd_ip.t22 dvdd_ip.t18 312.123
R2204 dvdd_ip.t23 dvdd_ip.n70 259.716
R2205 dvdd_ip.t18 dvdd_ip.n71 259.716
R2206 dvdd_ip.t24 dvdd_ip.n79 250.107
R2207 dvdd_ip.n81 dvdd_ip.t29 250.107
R2208 dvdd_ip.n2 dvdd_ip.n26 221.308
R2209 dvdd_ip.n80 dvdd_ip.t34 198.903
R2210 dvdd_ip.t42 dvdd_ip.n80 198.903
R2211 dvdd_ip.t9 dvdd_ip.n91 159.988
R2212 dvdd_ip.n91 dvdd_ip.t7 159.988
R2213 dvdd_ip.n73 dvdd_ip.t19 156.062
R2214 dvdd_ip.n73 dvdd_ip.t22 156.062
R2215 dvdd_ip.n24 dvdd_ip.n23 146.071
R2216 dvdd_ip.n82 dvdd_ip.n0 138.667
R2217 dvdd_ip.n51 dvdd_ip.t43 126.082
R2218 dvdd_ip.n54 dvdd_ip.t39 115.43
R2219 dvdd_ip.n52 dvdd_ip.t46 115.43
R2220 dvdd_ip.n77 dvdd_ip.t47 115.43
R2221 dvdd_ip.n75 dvdd_ip.t41 115.43
R2222 dvdd_ip.n1 dvdd_ip.t33 113.624
R2223 dvdd_ip.n4 dvdd_ip.t51 113.624
R2224 dvdd_ip.n21 dvdd_ip.t48 113.624
R2225 dvdd_ip.n1 dvdd_ip.t45 113.501
R2226 dvdd_ip.n4 dvdd_ip.t35 113.501
R2227 dvdd_ip.n55 dvdd_ip.t50 111.784
R2228 dvdd_ip.n54 dvdd_ip.t49 111.784
R2229 dvdd_ip.n53 dvdd_ip.t31 111.784
R2230 dvdd_ip.n52 dvdd_ip.t30 111.784
R2231 dvdd_ip.n77 dvdd_ip.t37 111.784
R2232 dvdd_ip.n78 dvdd_ip.t36 111.784
R2233 dvdd_ip.n75 dvdd_ip.t26 111.784
R2234 dvdd_ip.n76 dvdd_ip.t25 111.784
R2235 dvdd_ip.n22 dvdd_ip.t28 111.784
R2236 dvdd_ip.n22 dvdd_ip.t52 111.784
R2237 dvdd_ip.n51 dvdd_ip.t44 111.784
R2238 dvdd_ip.n35 dvdd_ip.n34 106.282
R2239 dvdd_ip.n38 dvdd_ip.n37 106.282
R2240 dvdd_ip.n27 dvdd_ip 1.37849
R2241 dvdd_ip.n68 dvdd_ip.n50 89.4643
R2242 dvdd_ip.n17 dvdd_ip.n82 64.1367
R2243 dvdd_ip.n28 dvdd_ip.t21 60.3236
R2244 dvdd_ip.n84 dvdd_ip.t15 57.1305
R2245 dvdd_ip.n84 dvdd_ip.t13 57.1305
R2246 dvdd_ip.n83 dvdd_ip.t10 57.1305
R2247 dvdd_ip.n83 dvdd_ip.t8 57.1305
R2248 dvdd_ip.n85 dvdd_ip.n19 55.1223
R2249 dvdd_ip.n111 dvdd_ip.n108 54.7105
R2250 dvdd_ip.n111 dvdd_ip.n106 54.7105
R2251 dvdd_ip.n111 dvdd_ip.n109 54.7085
R2252 dvdd_ip.n111 dvdd_ip.n107 54.7085
R2253 dvdd_ip.n111 dvdd_ip.n110 54.7085
R2254 dvdd_ip.n88 dvdd_ip.n48 53.6981
R2255 dvdd_ip.n14 dvdd_ip.n30 46.6446
R2256 dvdd_ip.n62 dvdd_ip.n49 46.2505
R2257 dvdd_ip.n66 dvdd_ip.n65 46.2505
R2258 dvdd_ip.n36 dvdd_ip.n31 46.2505
R2259 dvdd_ip.n32 dvdd_ip.n30 46.2505
R2260 dvdd_ip.n34 dvdd_ip.n32 44.5206
R2261 dvdd_ip.n37 dvdd_ip.n36 44.5206
R2262 dvdd_ip.n18 dvdd_ip.n16 0.871339
R2263 dvdd_ip.n67 dvdd_ip.n66 37.2058
R2264 dvdd_ip.n93 dvdd_ip.n15 37.0005
R2265 dvdd_ip.n5 dvdd_ip.n96 37.0005
R2266 dvdd_ip.n89 dvdd_ip.n19 33.5615
R2267 dvdd_ip.n10 dvdd_ip.n9 1.04644
R2268 dvdd_ip.n68 dvdd_ip.n67 31.3351
R2269 dvdd_ip.n15 dvdd_ip.n92 26.4291
R2270 dvdd_ip.n90 dvdd_ip.n89 26.4291
R2271 dvdd_ip.n61 dvdd_ip.n6 12.8793
R2272 dvdd_ip.n14 dvdd_ip.n105 23.3225
R2273 dvdd_ip.n67 dvdd_ip.n7 22.576
R2274 dvdd_ip.n85 dvdd_ip.n46 20.5561
R2275 dvdd_ip.n91 dvdd_ip.n46 20.5561
R2276 dvdd_ip.n87 dvdd_ip.n47 20.5561
R2277 dvdd_ip.n91 dvdd_ip.n47 20.5561
R2278 dvdd_ip.n87 dvdd_ip.n48 19.0763
R2279 dvdd_ip.n2 dvdd_ip.n0 18.9635
R2280 dvdd_ip.n89 dvdd_ip.n88 17.7956
R2281 dvdd_ip.n86 dvdd_ip.n5 17.833
R2282 dvdd_ip.n20 dvdd_ip.n86 17.8749
R2283 dvdd_ip.n78 dvdd_ip.n77 14.6565
R2284 dvdd_ip.n76 dvdd_ip.n75 14.6565
R2285 dvdd_ip.n53 dvdd_ip.n52 14.6565
R2286 dvdd_ip.n55 dvdd_ip.n54 14.6565
R2287 dvdd_ip.n59 dvdd_ip.n16 10.2385
R2288 dvdd_ip.n12 dvdd_ip.n28 0.591844
R2289 dvdd_ip.n20 dvdd_ip.n85 13.513
R2290 dvdd_ip.n86 dvdd_ip.n45 13.2148
R2291 dvdd_ip.n95 dvdd_ip.n28 13.2148
R2292 dvdd_ip.n70 dvdd_ip.n69 12.3338
R2293 dvdd_ip.n71 dvdd_ip.n0 12.3338
R2294 dvdd_ip.n24 dvdd_ip.n81 11.563
R2295 dvdd_ip.n66 dvdd_ip.n59 11.1792
R2296 dvdd_ip.n8 dvdd_ip.n13 1.8903
R2297 dvdd_ip.n18 dvdd_ip.n68 11.0012
R2298 dvdd_ip.n25 dvdd_ip.n23 139.684
R2299 dvdd_ip.n45 dvdd_ip.n44 9.84115
R2300 dvdd_ip.n95 dvdd_ip.n94 9.84115
R2301 dvdd_ip.n88 dvdd_ip.n9 9.4314
R2302 dvdd_ip dvdd_ip.n56 9.39134
R2303 dvdd_ip.n18 dvdd_ip.n29 9.30175
R2304 dvdd_ip.n25 dvdd_ip.n2 1.1019
R2305 dvdd_ip.n17 dvdd_ip.n50 8.03454
R2306 dvdd_ip.n57 dvdd_ip.n27 15.3109
R2307 dvdd_ip.n64 dvdd_ip.n7 7.4005
R2308 dvdd_ip.n39 dvdd_ip.n38 7.4005
R2309 dvdd_ip.n35 dvdd_ip.n33 7.4005
R2310 dvdd_ip.n6 dvdd_ip.n18 0.167749
R2311 dvdd_ip.n109 dvdd_ip.t5 7.14175
R2312 dvdd_ip.n109 dvdd_ip.t12 7.14175
R2313 dvdd_ip.n108 dvdd_ip.t3 7.14175
R2314 dvdd_ip.n108 dvdd_ip.t55 7.14175
R2315 dvdd_ip.n107 dvdd_ip.t6 7.14175
R2316 dvdd_ip.n107 dvdd_ip.t54 7.14175
R2317 dvdd_ip.n106 dvdd_ip.t11 7.14175
R2318 dvdd_ip.n106 dvdd_ip.t53 7.14175
R2319 dvdd_ip.n110 dvdd_ip.t4 7.14175
R2320 dvdd_ip.n110 dvdd_ip.t2 7.14175
R2321 dvdd_ip.n26 dvdd_ip.n74 6.37981
R2322 dvdd_ip.n74 dvdd_ip.n73 6.37981
R2323 dvdd_ip.n72 dvdd_ip.n50 6.37981
R2324 dvdd_ip.n73 dvdd_ip.n72 6.37981
R2325 dvdd_ip.n49 dvdd_ip.n19 5.51614
R2326 dvdd_ip.n61 dvdd_ip.n60 5.18874
R2327 dvdd_ip.n64 dvdd_ip.n63 5.18874
R2328 dvdd_ip.n13 dvdd_ip.n40 5.53168
R2329 dvdd_ip.n97 dvdd_ip.n14 4.95261
R2330 dvdd_ip.n25 dvdd_ip.n82 3.23758
R2331 dvdd_ip.n20 dvdd_ip.n8 0.738278
R2332 dvdd_ip.n8 dvdd_ip.n87 3.8204
R2333 dvdd_ip.n24 dvdd_ip 3.55088
R2334 dvdd_ip.t20 dvdd_ip.n44 3.32862
R2335 dvdd_ip.n94 dvdd_ip.t20 3.32862
R2336 dvdd_ip.n9 dvdd_ip.n19 3.14232
R2337 dvdd_ip.n2 dvdd_ip.n78 3.1045
R2338 dvdd_ip.n2 dvdd_ip.n76 3.1045
R2339 dvdd_ip.n24 dvdd_ip.n55 3.1045
R2340 dvdd_ip.n12 dvdd_ip.n8 0.0238734
R2341 dvdd_ip.n80 dvdd_ip.n57 2.76169
R2342 dvdd_ip.n58 dvdd_ip.n23 2.76169
R2343 dvdd_ip.n80 dvdd_ip.n58 2.76169
R2344 dvdd_ip.n10 dvdd_ip.n49 2.74244
R2345 dvdd_ip.n69 dvdd_ip.n18 2.32363
R2346 dvdd_ip.n63 dvdd_ip.t0 2.20373
R2347 dvdd_ip.t0 dvdd_ip.n60 2.20373
R2348 dvdd_ip.n97 dvdd_ip.n42 2.07915
R2349 dvdd_ip.n101 dvdd_ip.n42 2.07915
R2350 dvdd_ip.n41 dvdd_ip.n40 2.07915
R2351 dvdd_ip.n43 dvdd_ip.n41 2.07915
R2352 dvdd_ip.n10 dvdd_ip.n48 9.20625
R2353 dvdd_ip.n21 dvdd_ip.n51 1.71757
R2354 dvdd_ip.n27 dvdd_ip.n2 1.42317
R2355 dvdd_ip.n56 dvdd_ip.n30 1.51323
R2356 dvdd_ip.n16 dvdd_ip.n26 82.9703
R2357 dvdd_ip.n24 dvdd_ip.n53 3.23543
R2358 dvdd_ip.n37 dvdd_ip.t16 1.22055
R2359 dvdd_ip.n34 dvdd_ip.t16 1.22055
R2360 dvdd_ip.n9 dvdd_ip.n7 1.02666
R2361 dvdd_ip.n9 dvdd_ip.n8 0.868735
R2362 dvdd_ip.n66 dvdd_ip.n29 0.83013
R2363 dvdd_ip.n18 dvdd_ip.n17 0.810159
R2364 dvdd_ip.n99 dvdd_ip.n98 0.768135
R2365 dvdd_ip.n100 dvdd_ip.n99 0.768135
R2366 dvdd_ip.n104 dvdd_ip.n103 0.768135
R2367 dvdd_ip.n103 dvdd_ip.n102 0.768135
R2368 dvdd_ip.n3 dvdd_ip 0.748986
R2369 dvdd_ip.n1 dvdd_ip.n4 0.726273
R2370 dvdd_ip.n69 dvdd_ip.n59 0.70655
R2371 dvdd_ip.n3 dvdd_ip.n21 0.67791
R2372 dvdd_ip.n8 dvdd_ip.n11 0.621489
R2373 dvdd_ip.n111 dvdd_ip 0.569502
R2374 dvdd_ip.n79 dvdd_ip.n2 11.6172
R2375 dvdd_ip.n17 dvdd_ip.n2 1.64329
R2376 dvdd_ip dvdd_ip.n14 0.563996
R2377 dvdd_ip.n9 dvdd_ip.n6 0.547509
R2378 dvdd_ip.n3 dvdd_ip.n22 0.721964
R2379 dvdd_ip.n8 dvdd_ip.t56 0.442304
R2380 dvdd_ip.n2 dvdd_ip.n1 0.719176
R2381 dvdd_ip.n15 dvdd_ip.n12 1.41519
R2382 dvdd_ip.n5 dvdd_ip.n13 1.39615
R2383 dvdd_ip.n1 dvdd_ip.n3 1.26452
R2384 tail tail.t6 113.688
R2385 tail.n3 tail.t5 113.688
R2386 tail tail.t8 113.624
R2387 tail.n0 tail.t4 113.562
R2388 tail.n0 tail.t9 113.562
R2389 tail.n1 tail.t7 113.562
R2390 tail.n1 tail.t2 113.562
R2391 tail tail.t3 113.501
R2392 tail tail.t11 113.438
R2393 tail.n3 tail.t10 113.438
R2394 tail tail.n2 53.5531
R2395 tail.n2 tail.t0 6.92425
R2396 tail.n2 tail.t1 6.92425
R2397 tail tail.n1 1.9055
R2398 tail.n1 tail.n0 1.13844
R2399 tail.n3 tail 1.13636
R2400 a_16273_n2549.n3 a_16273_n2549.n2 647.119
R2401 a_16273_n2549.n1 a_16273_n2549.t4 350.253
R2402 a_16273_n2549.n2 a_16273_n2549.n0 260.339
R2403 a_16273_n2549.n2 a_16273_n2549.n1 246.119
R2404 a_16273_n2549.n1 a_16273_n2549.t5 189.588
R2405 a_16273_n2549.n3 a_16273_n2549.t3 89.1195
R2406 a_16273_n2549.n0 a_16273_n2549.t1 63.3338
R2407 a_16273_n2549.t0 a_16273_n2549.n3 41.0422
R2408 a_16273_n2549.n0 a_16273_n2549.t2 31.9797
R2409 a_16151_n2791.t0 a_16151_n2791.t1 198.571
R2410 a_16317_n2791.t0 a_16317_n2791.t1 60.0005
R2411 standby_b.n18 standby_b.t16 408.63
R2412 standby_b.n20 standby_b.t27 408.63
R2413 standby_b.n22 standby_b.t13 408.63
R2414 standby_b.n12 standby_b.t8 401.051
R2415 standby_b.t8 standby_b.n11 401.051
R2416 standby_b.t21 standby_b.n3 401.051
R2417 standby_b.n4 standby_b.t21 401.051
R2418 standby_b.n12 standby_b.t18 371.31
R2419 standby_b.t18 standby_b.n11 371.31
R2420 standby_b.t20 standby_b.n13 371.31
R2421 standby_b.n14 standby_b.t20 371.31
R2422 standby_b.t2 standby_b.n10 371.31
R2423 standby_b.n15 standby_b.t2 371.31
R2424 standby_b.n17 standby_b.t5 371.31
R2425 standby_b.t5 standby_b.n16 371.31
R2426 standby_b.n9 standby_b.t23 371.31
R2427 standby_b.t23 standby_b.n8 371.31
R2428 standby_b.t25 standby_b.n2 371.31
R2429 standby_b.n7 standby_b.t25 371.31
R2430 standby_b.t9 standby_b.n5 371.31
R2431 standby_b.n6 standby_b.t9 371.31
R2432 standby_b.n4 standby_b.t19 371.31
R2433 standby_b.t19 standby_b.n3 371.31
R2434 standby_b.n26 standby_b.t15 347.577
R2435 standby_b.n25 standby_b.t17 347.577
R2436 standby_b.n24 standby_b.t4 347.577
R2437 standby_b.t14 standby_b.n0 166.376
R2438 standby_b.n0 standby_b.t6 166.207
R2439 standby_b.n0 standby_b.t1 3.2348
R2440 standby_b.n27 standby_b.t26 236.552
R2441 standby_b.t1 standby_b.t0 228.429
R2442 standby_b.n26 standby_b.t10 193.337
R2443 standby_b.n25 standby_b.t11 193.337
R2444 standby_b.n24 standby_b.t24 193.337
R2445 x7.x2.x4.RESET_B standby_b.n18 165.089
R2446 x7.x2.x4.RESET_B standby_b.n20 165.089
R2447 x7.x2.x4.RESET_B standby_b.n22 165.089
R2448 standby_b.n27 standby_b.t12 164.251
R2449 x7.x3.A1 standby_b.n27 154.47
R2450 x7.x2.x2.RESET_B standby_b.n26 152
R2451 x7.x2.x3.RESET_B standby_b.n25 152
R2452 x7.x2.x4.RESET_B standby_b.n24 152
R2453 standby_b.n18 standby_b.t3 132.282
R2454 standby_b.n20 standby_b.t7 132.282
R2455 standby_b.n22 standby_b.t22 132.282
R2456 standby_b.n6 standby_b.n3 29.7417
R2457 standby_b.n7 standby_b.n6 29.7417
R2458 standby_b.n8 standby_b.n7 29.7417
R2459 standby_b.n16 standby_b.n15 29.7417
R2460 standby_b.n15 standby_b.n14 29.7417
R2461 standby_b.n14 standby_b.n11 29.7417
R2462 standby_b.n5 standby_b.n4 29.7417
R2463 standby_b.n5 standby_b.n2 29.7417
R2464 standby_b.n9 standby_b.n2 29.7417
R2465 standby_b.n17 standby_b.n10 29.7417
R2466 standby_b.n13 standby_b.n10 29.7417
R2467 standby_b.n13 standby_b.n12 29.7417
R2468 standby_b.n8 standby_b.n1 17.6946
R2469 standby_b.n1 standby_b.n9 17.5064
R2470 standby_b.n19 x7.x2.x4.RESET_B 16.7098
R2471 standby_b.n1 x7.stby_b 15.0825
R2472 x7.x2.x2.RESET_B standby_b.n19 14.0185
R2473 x7.x2.x3.RESET_B standby_b.n21 14.0185
R2474 x7.x2.x4.RESET_B standby_b.n23 14.0185
R2475 x7.stby_b x7.x3.A1 13.8064
R2476 standby_b.n1 standby_b.n17 12.2358
R2477 standby_b.n16 standby_b.n1 12.0476
R2478 standby_b.n19 x7.x2.x2.RESET_B 11.4672
R2479 standby_b.n21 x7.x2.x3.RESET_B 11.4672
R2480 standby_b.n23 x7.x2.x4.RESET_B 11.4672
R2481 x7.stby_b x7.x2.x4.RESET_B 10.5569
R2482 standby_b.t1 standby_b.n1 10.4718
R2483 standby_b.n23 x7.x2.x4.RESET_B 9.3005
R2484 x7.x2.x4.RESET_B x7.x2.x3.RESET_B 9.3005
R2485 standby_b.n21 x7.x2.x4.RESET_B 9.3005
R2486 x7.x2.x4.RESET_B x7.x2.x2.RESET_B 9.3005
R2487 a_9120_n9346.n1 a_9120_n9346.t2 649.659
R2488 a_9120_n9346.n0 a_9120_n9346.t4 227.685
R2489 a_9120_n9346.t0 a_9120_n9346.n2 44.6806
R2490 a_9120_n9346.n1 a_9120_n9346.t1 5.45407
R2491 a_9120_n9346.n0 a_9120_n9346.t3 5.07473
R2492 a_9120_n9346.n2 a_9120_n9346.n0 0.639781
R2493 a_9120_n9346.n2 a_9120_n9346.n1 0.0621233
R2494 a_24220_n9832.t0 a_24220_n9832.t1 83.56
R2495 a_16974_n1881.t0 a_16974_n1881.t1 87.1434
R2496 a_16795_n1943.n6 a_16795_n1943.n5 746.659
R2497 a_16795_n1943.n0 a_16795_n1943.t8 389.183
R2498 a_16795_n1943.n2 a_16795_n1943.t4 256.988
R2499 a_16795_n1943.n1 a_16795_n1943.n0 251.167
R2500 a_16795_n1943.n1 a_16795_n1943.t1 223.571
R2501 a_16795_n1943.n4 a_16795_n1943.t5 212.081
R2502 a_16795_n1943.n5 a_16795_n1943.n4 181.942
R2503 a_16795_n1943.n0 a_16795_n1943.t7 174.891
R2504 a_16795_n1943.n2 a_16795_n1943.t6 163.803
R2505 a_16795_n1943.n3 a_16795_n1943.t3 139.78
R2506 a_16795_n1943.n3 a_16795_n1943.n2 129.264
R2507 a_16795_n1943.n6 a_16795_n1943.t2 63.3219
R2508 a_16795_n1943.t0 a_16795_n1943.n6 63.3219
R2509 a_16795_n1943.n5 a_16795_n1943.n1 24.6993
R2510 a_16795_n1943.n4 a_16795_n1943.n3 22.6399
R2511 a_21775_n2247.t0 a_21775_n2247.n1 386.31
R2512 a_21775_n2247.n1 a_21775_n2247.t1 249.956
R2513 a_21775_n2247.n0 a_21775_n2247.t2 239.04
R2514 a_21775_n2247.n1 a_21775_n2247.n0 175.661
R2515 a_21775_n2247.n0 a_21775_n2247.t3 166.739
R2516 x7.ena_done_b.n8 x7.ena_done_b.t0 373.866
R2517 x7.ena_done_b.n6 x7.ena_done_b.t5 333.651
R2518 x7.ena_done_b.n6 x7.ena_done_b.t6 297.233
R2519 x7.ena_done_b x7.ena_done_b.t1 247.159
R2520 x7.ena_done_b.n0 x7.ena_done_b.t3 241.536
R2521 x7.ena_done_b.n2 x7.ena_done_b.t4 207.423
R2522 x7.ena_done_b.n3 x7.ena_done_b.t7 202.133
R2523 x7.ena_done_b x7.ena_done_b.n6 195.701
R2524 x7.ena_done_b.n0 x7.ena_done_b.t2 169.237
R2525 x7.ena_done_b.n5 x7.ena_done_b.n2 159.758
R2526 x7.ena_done_b.n1 x7.ena_done_b.n0 155.84
R2527 x7.ena_done_b.n4 x7.ena_done_b.n3 152
R2528 x7.ena_done_b.n3 x7.ena_done_b.n2 36.8275
R2529 x7.ena_done_b x7.ena_done_b.n8 16.6907
R2530 x7.ena_done_b.n7 x7.ena_done_b 15.8995
R2531 x7.ena_done_b.n7 x7.ena_done_b 15.6656
R2532 x7.ena_done_b x7.ena_done_b.n5 13.8109
R2533 x7.ena_done_b x7.ena_done_b.n1 11.2245
R2534 x7.ena_done_b.n5 x7.ena_done_b.n4 5.4308
R2535 x7.ena_done_b.n4 x7.ena_done_b 3.68535
R2536 x7.ena_done_b.n1 x7.ena_done_b 3.2005
R2537 x7.ena_done_b.n8 x7.ena_done_b.n7 3.1005
R2538 a_20121_n2241.t0 a_20121_n2241.n3 370.026
R2539 a_20121_n2241.n0 a_20121_n2241.t2 351.356
R2540 a_20121_n2241.n1 a_20121_n2241.t4 334.717
R2541 a_20121_n2241.n3 a_20121_n2241.t1 325.971
R2542 a_20121_n2241.n1 a_20121_n2241.t5 309.935
R2543 a_20121_n2241.n0 a_20121_n2241.t3 305.683
R2544 a_20121_n2241.n2 a_20121_n2241.n0 16.879
R2545 a_20121_n2241.n3 a_20121_n2241.n2 10.8867
R2546 a_20121_n2241.n2 a_20121_n2241.n1 9.3005
R2547 a_2130_n21176.t0 a_2130_n21176.t1 82.0028
R2548 a_24530_n21342.t0 a_24530_n21342.t1 81.9492
R2549 standby_33.n0 standby_33.t0 227.886
R2550 standby_33 standby_33.t3 216.05
R2551 standby_33.n0 standby_33.n1 25.0903
R2552 standby_33.n0 standby_33.t4 12.7763
R2553 standby_33.n1 standby_33.t1 5.5105
R2554 standby_33.n1 standby_33.t2 5.5105
R2555 standby_33.n0 standby_33 1.67737
R2556 ibias.n7 ibias.n1 1544.9
R2557 ibias.n4 ibias.n3 1544.9
R2558 ibias.n2 ibias.n0 300.425
R2559 ibias.n8 ibias.n2 300.425
R2560 ibias.n9 ibias.n0 177.746
R2561 ibias.n9 ibias.n8 177.746
R2562 ibias.n5 ibias.n1 139.143
R2563 ibias.n6 ibias.n3 139.143
R2564 ibias.n9 ibias.t1 60.1061
R2565 ibias.n4 ibias.n0 46.2505
R2566 ibias.n8 ibias.n7 46.2505
R2567 ibias.n5 ibias.n4 40.8622
R2568 ibias.n7 ibias.n6 40.8622
R2569 ibias.n3 ibias.n2 12.3338
R2570 ibias.n9 ibias.n1 12.3338
R2571 ibias.n6 ibias.t0 4.16651
R2572 ibias.t0 ibias.n5 4.16651
R2573 ibias ibias.n9 1.58676
R2574 ibias_ip ibias_ip.t13 31.8332
R2575 ibias_ip.t12 ibias_ip 31.4808
R2576 ibias_ip ibias_ip.t0 61.7027
R2577 ibias_ip.t1 ibias_ip 31.3394
R2578 ibias_ip ibias_ip.t2 39.498
R2579 ibias_ip.n0 ibias_ip.t11 31.8633
R2580 ibias_ip ibias_ip.t7 31.1832
R2581 ibias_ip.n1 ibias_ip.t3 31.1727
R2582 ibias_ip.n0 ibias_ip.t9 31.193
R2583 ibias_ip.n0 ibias_ip.t5 31.1967
R2584 ibias_ip.t4 ibias_ip.n1 39.8957
R2585 ibias_ip ibias_ip.t8 39.8329
R2586 ibias_ip.t6 ibias_ip.n0 39.8506
R2587 ibias_ip.n0 ibias_ip.t10 39.8715
R2588 ibias_ip ibias_ip.n1 1.87886
R2589 ibias_ip ibias_ip.n0 1.34188
R2590 avdd_ip.n53 avdd_ip.n49 58547.9
R2591 avdd_ip.n55 avdd_ip.n49 58547.9
R2592 avdd_ip.n54 avdd_ip.n53 58547.9
R2593 avdd_ip.n55 avdd_ip.n54 58547.9
R2594 avdd_ip.n77 avdd_ip.n76 50679.6
R2595 avdd_ip.n52 avdd_ip.n47 28978.4
R2596 avdd_ip.n56 avdd_ip.n47 28978.4
R2597 avdd_ip.n52 avdd_ip.n48 28978.4
R2598 avdd_ip.n56 avdd_ip.n48 28978.4
R2599 avdd_ip.n95 avdd_ip.n15 7296
R2600 avdd_ip.n93 avdd_ip.n15 7296
R2601 avdd_ip.n95 avdd_ip.n16 7296
R2602 avdd_ip.n93 avdd_ip.n16 7296
R2603 avdd_ip.n57 avdd_ip.n25 6735.06
R2604 avdd_ip.n51 avdd_ip.n25 6735.06
R2605 avdd_ip.n51 avdd_ip.n50 3209.98
R2606 avdd_ip.n86 avdd_ip.n57 2921.68
R2607 avdd_ip.n79 avdd_ip.n78 857.648
R2608 avdd_ip.n81 avdd_ip.n73 857.648
R2609 avdd_ip.n78 avdd_ip.n73 857.648
R2610 avdd_ip.n67 avdd_ip.n60 857.648
R2611 avdd_ip.n64 avdd_ip.n61 857.648
R2612 avdd_ip.n77 avdd_ip.t2 337.433
R2613 avdd_ip.n65 avdd_ip.n64 267.182
R2614 avdd_ip.n67 avdd_ip.n66 267.182
R2615 avdd_ip.n81 avdd_ip.n80 267.182
R2616 avdd_ip.n24 avdd_ip.n23 212.139
R2617 avdd_ip.n92 avdd_ip.n91 202.696
R2618 avdd_ip.n87 avdd_ip.n24 201.294
R2619 avdd_ip.n90 avdd_ip.n18 134.065
R2620 avdd_ip.n50 avdd_ip.n18 110.358
R2621 avdd_ip.t7 avdd_ip.n15 105.665
R2622 avdd_ip.t11 avdd_ip.n16 105.665
R2623 avdd_ip.n64 avdd_ip.n63 92.5005
R2624 avdd_ip.n60 avdd_ip.n59 92.5005
R2625 avdd_ip.n68 avdd_ip.n67 92.5005
R2626 avdd_ip.n62 avdd_ip.n61 92.5005
R2627 avdd_ip.n78 avdd_ip.n75 92.5005
R2628 avdd_ip.n78 avdd_ip.n77 92.5005
R2629 avdd_ip.n74 avdd_ip.n73 92.5005
R2630 avdd_ip.t2 avdd_ip.n73 92.5005
R2631 avdd_ip.n82 avdd_ip.n81 92.5005
R2632 avdd_ip.n79 avdd_ip.n72 92.5005
R2633 avdd_ip.n63 avdd_ip.n59 91.4872
R2634 avdd_ip.n75 avdd_ip.n72 91.4829
R2635 avdd_ip.n94 avdd_ip.t7 79.5673
R2636 avdd_ip.n94 avdd_ip.t11 79.5673
R2637 avdd_ip.n87 avdd_ip.n86 75.3225
R2638 avdd_ip.n63 avdd_ip.n62 66.8331
R2639 avdd_ip.n75 avdd_ip.n74 66.3131
R2640 avdd_ip.n69 avdd_ip.n59 63.936
R2641 avdd_ip.n83 avdd_ip.n72 63.936
R2642 avdd_ip.n2 avdd_ip.t1 62.0945
R2643 avdd_ip.n39 avdd_ip.t23 61.1041
R2644 avdd_ip.n37 avdd_ip.t24 60.1061
R2645 avdd_ip.n33 avdd_ip.t21 60.1061
R2646 avdd_ip.n34 avdd_ip.t26 60.1061
R2647 avdd_ip.n31 avdd_ip.t20 60.1061
R2648 avdd_ip.n91 avdd_ip.t15 60.1061
R2649 avdd_ip.n91 avdd_ip.t12 60.1061
R2650 avdd_ip.n91 avdd_ip.t13 60.1061
R2651 avdd_ip.n23 avdd_ip.t10 60.1061
R2652 avdd_ip.n23 avdd_ip.t8 60.1061
R2653 avdd_ip.n23 avdd_ip.t9 60.1061
R2654 avdd_ip.n20 avdd_ip.t16 60.1061
R2655 avdd_ip.n20 avdd_ip.t14 60.1061
R2656 avdd_ip.n19 avdd_ip.t18 60.1061
R2657 avdd_ip.n19 avdd_ip.t17 60.1061
R2658 avdd_ip.n28 avdd_ip.t27 60.1061
R2659 avdd_ip.n28 avdd_ip.t19 60.1061
R2660 avdd_ip.n27 avdd_ip.t28 60.1061
R2661 avdd_ip.n27 avdd_ip.t22 60.1061
R2662 avdd_ip.n38 avdd_ip.t25 60.1061
R2663 avdd_ip.n80 avdd_ip.n79 57.4849
R2664 avdd_ip.n65 avdd_ip.n60 57.4849
R2665 avdd_ip.n66 avdd_ip.n61 57.4849
R2666 avdd_ip.n2 avdd_ip.n1 55.1707
R2667 avdd_ip.n2 avdd_ip.n0 54.9038
R2668 avdd_ip.n44 avdd_ip.n26 44.6614
R2669 avdd_ip.n68 avdd_ip.n58 43.3376
R2670 avdd_ip.n82 avdd_ip.n71 43.3376
R2671 avdd_ip.n46 avdd_ip.n45 30.1747
R2672 avdd_ip.n66 avdd_ip.t5 28.8172
R2673 avdd_ip.t5 avdd_ip.n65 28.8172
R2674 avdd_ip.n80 avdd_ip.t2 28.8172
R2675 avdd_ip.n92 avdd_ip.n17 10.6324
R2676 avdd_ip.n98 avdd_ip.n97 9.3005
R2677 avdd_ip.n50 avdd_ip.n14 8.37369
R2678 avdd_ip.n38 avdd_ip.n37 7.25561
R2679 avdd_ip.n0 avdd_ip.t4 6.92425
R2680 avdd_ip.n0 avdd_ip.t3 6.92425
R2681 avdd_ip.n1 avdd_ip.t6 6.92425
R2682 avdd_ip.n1 avdd_ip.t0 6.92425
R2683 avdd_ip.n93 avdd_ip.n92 6.37981
R2684 avdd_ip.n94 avdd_ip.n93 6.37981
R2685 avdd_ip.n96 avdd_ip.n95 6.37981
R2686 avdd_ip.n95 avdd_ip.n94 6.37981
R2687 avdd_ip.n32 avdd_ip.n31 6.17839
R2688 avdd_ip.n96 avdd_ip.n14 5.31953
R2689 avdd_ip.n62 avdd_ip.n58 4.38907
R2690 avdd_ip.n74 avdd_ip.n71 4.38907
R2691 avdd_ip.n97 avdd_ip.n96 3.70667
R2692 avdd_ip.n46 avdd_ip.n24 3.6009
R2693 avdd_ip.n84 avdd_ip.n71 2.4925
R2694 avdd_ip.n70 avdd_ip.n58 2.44611
R2695 avdd_ip.n18 avdd_ip.n16 2.43471
R2696 avdd_ip.n45 avdd_ip.n15 2.43471
R2697 avdd_ip.n69 avdd_ip.n68 2.37764
R2698 avdd_ip.n83 avdd_ip.n82 2.37764
R2699 avdd_ip.n70 avdd_ip.n69 2.3255
R2700 avdd_ip.n84 avdd_ip.n83 2.3255
R2701 avdd_ip.n88 avdd_ip.n87 2.09243
R2702 avdd_ip.n34 avdd_ip.n30 1.87566
R2703 avdd_ip.n26 avdd_ip.n13 1.57905
R2704 avdd_ip.n4 avdd_ip.n3 1.18871
R2705 avdd_ip.n33 avdd_ip.n32 1.07773
R2706 avdd_ip.n48 avdd_ip.n25 1.05764
R2707 avdd_ip.n54 avdd_ip.n48 1.05764
R2708 avdd_ip.n47 avdd_ip.n46 1.05764
R2709 avdd_ip.n49 avdd_ip.n47 1.05764
R2710 avdd_ip.n35 avdd_ip.n34 0.982678
R2711 avdd_ip.n35 avdd_ip.n33 0.919312
R2712 avdd_ip.n39 avdd_ip.n38 0.90347
R2713 avdd_ip.n32 avdd_ip.n30 0.845955
R2714 avdd_ip.n11 avdd_ip.n4 0.827286
R2715 avdd_ip avdd_ip.n11 0.808179
R2716 avdd_ip.n29 avdd_ip.n27 0.65712
R2717 avdd_ip.n21 avdd_ip.n19 0.652725
R2718 avdd_ip.n90 avdd_ip.n89 0.613954
R2719 avdd_ip.n57 avdd_ip.n56 0.530586
R2720 avdd_ip.n56 avdd_ip.n55 0.530586
R2721 avdd_ip.n52 avdd_ip.n51 0.530586
R2722 avdd_ip.n53 avdd_ip.n52 0.530586
R2723 avdd_ip.n3 avdd_ip.n2 0.507794
R2724 avdd_ip.n45 avdd_ip.n44 0.448948
R2725 avdd_ip.n40 avdd_ip.n36 0.402976
R2726 avdd_ip.n22 avdd_ip.n21 0.319749
R2727 avdd_ip.n89 avdd_ip.n88 0.319015
R2728 avdd_ip.n42 avdd_ip.n29 0.319015
R2729 avdd_ip.n41 avdd_ip.n40 0.319015
R2730 avdd_ip.n36 avdd_ip.n35 0.282318
R2731 avdd_ip.n11 avdd_ip.n10 0.255087
R2732 avdd_ip.n21 avdd_ip.n20 0.25137
R2733 avdd_ip.n29 avdd_ip.n28 0.25137
R2734 avdd_ip.n41 avdd_ip.n12 0.245735
R2735 avdd_ip avdd_ip.n99 0.213307
R2736 avdd_ip.n89 avdd_ip.n17 0.211864
R2737 avdd_ip.n40 avdd_ip.n39 0.211864
R2738 avdd_ip.n99 avdd_ip 0.18211
R2739 avdd_ip.n31 avdd_ip.n14 0.174542
R2740 avdd_ip.n37 avdd_ip.n26 0.174542
R2741 avdd_ip.n86 avdd_ip.n85 0.166571
R2742 avdd_ip.n42 avdd_ip.n41 0.150396
R2743 avdd_ip.n88 avdd_ip.n22 0.150396
R2744 avdd_ip.n3 avdd_ip.t33 0.125045
R2745 avdd_ip.n7 avdd_ip.n4 0.123905
R2746 avdd_ip.n43 avdd_ip.n22 0.117461
R2747 avdd_ip.n10 avdd_ip.n9 0.111971
R2748 avdd_ip.n8 avdd_ip.n7 0.110265
R2749 avdd_ip.n43 avdd_ip.n42 0.108384
R2750 avdd_ip.n6 avdd_ip.n5 0.106696
R2751 avdd_ip.n9 avdd_ip.n8 0.106696
R2752 avdd_ip.n85 avdd_ip.n70 0.0839309
R2753 avdd_ip.n85 avdd_ip.n84 0.0812962
R2754 avdd_ip.n5 avdd_ip.t30 0.0180781
R2755 avdd_ip.n9 avdd_ip.t32 0.0180781
R2756 avdd_ip.n8 avdd_ip.t29 0.0180781
R2757 avdd_ip.n6 avdd_ip.t31 0.0180781
R2758 avdd_ip.n10 avdd_ip.n5 0.0174228
R2759 avdd_ip.n13 avdd_ip.n12 0.0173478
R2760 avdd_ip.n23 avdd_ip.n17 0.0154184
R2761 avdd_ip.n91 avdd_ip.n90 0.0154184
R2762 avdd_ip.n7 avdd_ip.n6 0.0150053
R2763 avdd_ip.n97 avdd_ip.n13 0.0119388
R2764 avdd_ip.n44 avdd_ip.n43 0.0117727
R2765 avdd_ip.n99 avdd_ip.n98 0.00101125
R2766 avdd_ip.n36 avdd_ip.n30 0.000885802
R2767 avdd_ip.n98 avdd_ip.n12 0.000627812
R2768 xout.n29 xout.t26 594.784
R2769 xout.n29 xout.t24 194.649
R2770 xout.n25 xout.t23 124.457
R2771 xout.n25 xout.t25 106.793
R2772 xout.t23 xout.n24 86.3125
R2773 xout.t25 xout.n23 86.3125
R2774 xout.n3 xout.t14 62.0071
R2775 xout.n4 xout.t12 62.0071
R2776 xout.n3 xout.t19 60.1061
R2777 xout.n4 xout.t20 60.1061
R2778 xout.n8 xout.t10 60.1061
R2779 xout.n8 xout.t9 60.1061
R2780 xout.n10 xout.t13 60.1061
R2781 xout.n10 xout.t11 60.1061
R2782 xout.n0 xout.t16 60.1061
R2783 xout.n0 xout.t18 60.1061
R2784 xout.n1 xout.t15 60.1061
R2785 xout.n1 xout.t17 60.1061
R2786 xout.n24 xout.n23 58.6245
R2787 xout.n22 xout.t0 43.5339
R2788 xout.n28 xout.n27 21.3269
R2789 xout.n16 xout.n15 18.5533
R2790 xout.n20 xout.n13 18.553
R2791 xout.n19 xout.n18 18.4723
R2792 xout.n19 xout.n17 18.4564
R2793 xout.n16 xout.n14 18.4564
R2794 xout.n27 xout.n23 12.2455
R2795 xout.n18 xout.t1 4.133
R2796 xout.n18 xout.t8 4.133
R2797 xout.n17 xout.t21 4.133
R2798 xout.n17 xout.t22 4.133
R2799 xout.n15 xout.t2 4.133
R2800 xout.n15 xout.t4 4.133
R2801 xout.n14 xout.t3 4.133
R2802 xout.n14 xout.t6 4.133
R2803 xout.n13 xout.t5 4.133
R2804 xout.n13 xout.t7 4.133
R2805 xout.n5 xout.n4 3.64406
R2806 xout.n5 xout.n3 3.61238
R2807 xout.n26 xout.n24 3.56553
R2808 xout.n22 xout.n21 2.24362
R2809 xout.n29 xout.n28 2.18092
R2810 xout.n28 xout.n22 1.03102
R2811 xout.n27 xout.n26 0.742745
R2812 xout.n26 xout.n25 0.715885
R2813 xout.n21 xout.n12 0.464586
R2814 xout.n2 xout.n0 0.424187
R2815 xout.n11 xout.n9 0.402558
R2816 xout xout.n29 0.377063
R2817 xout.n6 xout.n2 0.316998
R2818 xout.n2 xout.n1 0.310571
R2819 xout.n12 xout.n7 0.273717
R2820 xout.n7 xout.n6 0.261913
R2821 xout.n9 xout.n8 0.254998
R2822 xout.n11 xout.n10 0.25137
R2823 xout.n6 xout.n5 0.143668
R2824 xout.n9 xout.n7 0.126918
R2825 xout.n12 xout.n11 0.125886
R2826 xout.n21 xout.n20 0.0947164
R2827 xout.n20 xout.n16 0.0657574
R2828 xout.n20 xout.n19 0.0480746
R2829 inv_in.n19 inv_in.t0 47.4896
R2830 inv_in.n18 inv_in.t3 6.48745
R2831 inv_in.n19 inv_in.t1 6.24255
R2832 inv_in inv_in.n17 2.2182
R2833 inv_in.n18 inv_in 0.342687
R2834 inv_in inv_in.n18 0.217687
R2835 inv_in.n5 inv_in.n4 0.110198
R2836 inv_in.n7 inv_in.n6 0.110101
R2837 inv_in.n10 inv_in.n9 0.110101
R2838 inv_in.n8 inv_in.n2 0.110101
R2839 inv_in.n16 inv_in.n15 0.109734
R2840 inv_in.n14 inv_in.n0 0.109734
R2841 inv_in.n13 inv_in.n12 0.109709
R2842 inv_in.n11 inv_in.n1 0.109709
R2843 inv_in.n9 inv_in.n7 0.109325
R2844 inv_in.n9 inv_in.n8 0.109325
R2845 inv_in.n12 inv_in.n11 0.109325
R2846 inv_in.n11 inv_in.n3 0.109325
R2847 inv_in.n15 inv_in.n14 0.1086
R2848 inv_in.n16 inv_in.n0 0.1086
R2849 inv_in.n4 inv_in.n3 0.10222
R2850 inv_in.n7 inv_in.n5 0.101755
R2851 inv_in inv_in.n19 0.09425
R2852 inv_in.n18 inv_in 0.063
R2853 inv_in.n0 inv_in.t11 0.00880157
R2854 inv_in.n7 inv_in.t9 0.00848368
R2855 inv_in.n9 inv_in.t10 0.00848368
R2856 inv_in.n8 inv_in.t2 0.00848368
R2857 inv_in.n5 inv_in.t12 0.00838586
R2858 inv_in.n4 inv_in.t14 0.0083125
R2859 inv_in.n6 inv_in.t13 0.0083125
R2860 inv_in.n2 inv_in.t6 0.0083125
R2861 inv_in.n10 inv_in.t4 0.0083125
R2862 inv_in.n1 inv_in.t5 0.0083125
R2863 inv_in.n13 inv_in.t8 0.0083125
R2864 inv_in.n17 inv_in.t7 0.0083125
R2865 inv_in.n6 inv_in.n3 0.00106244
R2866 inv_in.n12 inv_in.n2 0.00106244
R2867 inv_in.n11 inv_in.n10 0.00106244
R2868 inv_in.n17 inv_in.n16 0.000989074
R2869 inv_in.n15 inv_in.n1 0.000548907
R2870 inv_in.n14 inv_in.n13 0.000548907
R2871 inv_m1.t0 inv_m1.n0 652.083
R2872 inv_m1.n0 inv_m1.t1 229.685
R2873 inv_m1 inv_m1.n0 4.5555
R2874 inv_m1 inv_m1.n3 1.058
R2875 inv_m1.n3 inv_m1.n2 24.8426
R2876 inv_m1.n2 inv_m1.t4 20.438
R2877 inv_m1.n2 inv_m1.t3 20.4375
R2878 inv_m1.n3 inv_m1.n1 24.7082
R2879 inv_m1.n1 inv_m1.t5 21.9207
R2880 inv_m1.n1 inv_m1.t2 21.9202
R2881 a_2132_n15590.t0 a_2132_n15590.t1 82.3309
R2882 a_18932_n15756.t0 a_18932_n15756.t1 83.5579
R2883 inv_m2 inv_m2.t0 651.861
R2884 inv_m2 inv_m2.t1 229.522
R2885 inv_m2 inv_m2.t2 108.124
R2886 inv_m2.t5 inv_m2 108.124
R2887 inv_m2.n0 inv_m2 80.6505
R2888 inv_m2.t2 inv_m2.n0 27.4745
R2889 inv_m2.n0 inv_m2.t5 27.4745
R2890 inv_m2 inv_m2.n1 24.0208
R2891 inv_m2.n1 inv_m2.t3 20.4885
R2892 inv_m2.n1 inv_m2.t4 20.387
R2893 dout_ip.n0 dout_ip.t0 651.692
R2894 dout_ip.n0 dout_ip.t1 651.431
R2895 dout_ip.n1 dout_ip.t9 288.204
R2896 dout_ip.n5 dout_ip.t5 264.103
R2897 dout_ip.n2 dout_ip.t6 264.103
R2898 dout_ip.n0 dout_ip.t3 229.352
R2899 dout_ip.n0 dout_ip.t2 229.101
R2900 dout_ip.n1 dout_ip.t7 195.017
R2901 x7.x2.clkin dout_ip.n5 159.236
R2902 x7.x1.clkin dout_ip.n2 159.236
R2903 x7.x5.A dout_ip.n1 153.153
R2904 dout_ip.n4 x7.x2.x1.A 152
R2905 x7.x1.x1.A dout_ip.n3 152
R2906 dout_ip.n4 dout_ip.t8 145.209
R2907 dout_ip.n3 dout_ip.t4 145.209
R2908 dout_ip.n7 dout_ip.n6 117.519
R2909 dout_ip.n6 x7.x1.clkin 68.1959
R2910 dout_ip.n5 dout_ip.n4 37.6741
R2911 dout_ip.n3 dout_ip.n2 37.6741
R2912 x7.clkin dout_ip.n7 31.6505
R2913 dout_ip.n7 x7.x5.A 24.4485
R2914 x7.clkin dout_ip.n0 11.4719
R2915 x7.x2.clkin x7.x2.x1.A 10.3444
R2916 x7.x1.clkin x7.x1.x1.A 10.3444
R2917 dout_ip.n6 x7.x2.clkin 9.3005
R2918 a_20689_n2549.n3 a_20689_n2549.n2 647.119
R2919 a_20689_n2549.n1 a_20689_n2549.t4 350.253
R2920 a_20689_n2549.n2 a_20689_n2549.n0 260.339
R2921 a_20689_n2549.n2 a_20689_n2549.n1 246.119
R2922 a_20689_n2549.n1 a_20689_n2549.t5 189.588
R2923 a_20689_n2549.n3 a_20689_n2549.t2 89.1195
R2924 a_20689_n2549.n0 a_20689_n2549.t3 63.3338
R2925 a_20689_n2549.t0 a_20689_n2549.n3 41.0422
R2926 a_20689_n2549.n0 a_20689_n2549.t1 31.9797
R2927 a_20567_n2791.t1 a_20567_n2791.t0 198.571
R2928 a_20733_n2791.t0 a_20733_n2791.t1 60.0005
R2929 xin_buf.n0 xin_buf.t2 9.98044
R2930 xin_buf.n1 xin_buf.t3 6.0819
R2931 xin_buf.n0 xin_buf.t1 3.49292
R2932 xin_buf.n1 xin_buf.t4 2.23853
R2933 xin_buf.n1 xin_buf.t0 10.3359
R2934 xin_buf.n0 xin_buf.t0 28.8094
R2935 a_15000_n1881.n2 a_15000_n1881.n1 682.193
R2936 a_15000_n1881.n0 a_15000_n1881.t4 279.142
R2937 a_15000_n1881.n1 a_15000_n1881.t1 250.737
R2938 a_15000_n1881.n0 a_15000_n1881.t3 145.958
R2939 a_15000_n1881.n1 a_15000_n1881.n0 118.45
R2940 a_15000_n1881.n2 a_15000_n1881.t2 70.3576
R2941 a_15000_n1881.t0 a_15000_n1881.n2 65.6672
R2942 x7.x1.x2.CLK x7.x1.x2.CLK.t0 716.451
R2943 x7.x1.x2.CLK.t0 x7.x1.x2.CLK.n3 707.66
R2944 x7.x1.x2.CLK.n0 x7.x1.x2.CLK.t2 294.557
R2945 x7.x1.x2.CLK.n2 x7.x1.x2.CLK.t1 271.777
R2946 x7.x1.x2.CLK.n0 x7.x1.x2.CLK.t3 211.01
R2947 x7.x1.x2.CLK.n1 x7.x1.x2.CLK.n0 152
R2948 x7.x1.x2.CLK.n3 x7.x1.x2.CLK.n2 38.2982
R2949 x7.x1.x2.CLK.n2 x7.x1.x2.CLK.n1 33.0611
R2950 x7.x1.x2.CLK x7.x1.x2.CLK.n3 8.88521
R2951 x7.x1.x2.CLK.n1 x7.x1.x2.CLK 4.20621
R2952 a_16151_n1869.t1 a_16151_n1869.t0 198.571
R2953 a_16317_n1881.t0 a_16317_n1881.t1 60.0005
R2954 a_21775_n2791.t1 a_21775_n2791.n1 386.31
R2955 a_21775_n2791.n1 a_21775_n2791.t0 249.956
R2956 a_21775_n2791.n0 a_21775_n2791.t3 239.04
R2957 a_21775_n2791.n1 a_21775_n2791.n0 175.661
R2958 a_21775_n2791.n0 a_21775_n2791.t2 166.739
R2959 x7.clk_disable.n3 x7.clk_disable.t1 319.219
R2960 x7.clk_disable.n1 x7.clk_disable.t4 268.313
R2961 x7.clk_disable x7.clk_disable.t0 249.867
R2962 x7.clk_disable.n2 x7.clk_disable.t2 206.19
R2963 x7.clk_disable.n1 x7.clk_disable.t5 186.374
R2964 x7.clk_disable x7.clk_disable.n2 152
R2965 x7.clk_disable.n2 x7.clk_disable.n1 148.35
R2966 x7.clk_disable x7.clk_disable.n0 32.2121
R2967 x7.clk_disable x7.clk_disable.t3 21.881
R2968 x7.clk_disable.n3 x7.clk_disable 21.8175
R2969 x7.clk_disable.n0 x7.clk_disable 11.0708
R2970 x7.clk_disable.n0 x7.clk_disable 8.03187
R2971 x7.clk_disable x7.clk_disable.n3 4.14393
R2972 a_14009_n2701.t0 a_14009_n2701.n0 753.673
R2973 a_14009_n2701.n0 a_14009_n2701.t2 354.81
R2974 a_14009_n2701.n0 a_14009_n2701.t1 303.562
R2975 standby_ip.t0 standby_ip.n3 368.26
R2976 standby_ip.n2 standby_ip.n3 1.85916
R2977 standby_ip.n17 standby_ip.t4 405.389
R2978 standby_ip.t4 standby_ip.n16 405.389
R2979 standby_ip.t15 standby_ip.n8 405.389
R2980 standby_ip.n9 standby_ip.t15 405.389
R2981 standby_ip.n17 standby_ip.t6 375.649
R2982 standby_ip.t6 standby_ip.n16 375.649
R2983 standby_ip.t17 standby_ip.n18 375.649
R2984 standby_ip.n19 standby_ip.t17 375.649
R2985 standby_ip.t18 standby_ip.n15 375.649
R2986 standby_ip.n20 standby_ip.t18 375.649
R2987 standby_ip.n22 standby_ip.t5 375.649
R2988 standby_ip.t5 standby_ip.n21 375.649
R2989 standby_ip.n14 standby_ip.t11 375.649
R2990 standby_ip.t11 standby_ip.n13 375.649
R2991 standby_ip.t12 standby_ip.n7 375.649
R2992 standby_ip.n12 standby_ip.t12 375.649
R2993 standby_ip.t8 standby_ip.n10 375.649
R2994 standby_ip.n11 standby_ip.t8 375.649
R2995 standby_ip.n9 standby_ip.t9 375.649
R2996 standby_ip.t9 standby_ip.n8 375.649
R2997 standby_ip.t13 standby_ip.n23 332.752
R2998 standby_ip.n24 standby_ip.t13 332.75
R2999 standby_ip.t7 standby_ip.n23 332.411
R3000 standby_ip.n24 standby_ip.t7 332.411
R3001 standby_ip.n4 standby_ip.t3 231.718
R3002 standby_ip standby_ip.t1 216.155
R3003 standby_ip standby_ip.n5 161.314
R3004 standby_ip.n4 standby_ip.t14 159.417
R3005 standby_ip.n5 standby_ip.n4 152
R3006 standby_ip standby_ip.t16 59.9857
R3007 standby_ip standby_ip.t2 59.3654
R3008 standby_ip standby_ip.n2 46.2227
R3009 standby_ip.n11 standby_ip.n8 29.7417
R3010 standby_ip.n12 standby_ip.n11 29.7417
R3011 standby_ip.n13 standby_ip.n12 29.7417
R3012 standby_ip.n21 standby_ip.n20 29.7417
R3013 standby_ip.n20 standby_ip.n19 29.7417
R3014 standby_ip.n19 standby_ip.n16 29.7417
R3015 standby_ip.n10 standby_ip.n9 29.7417
R3016 standby_ip.n10 standby_ip.n7 29.7417
R3017 standby_ip.n14 standby_ip.n7 29.7417
R3018 standby_ip.n22 standby_ip.n15 29.7417
R3019 standby_ip.n18 standby_ip.n15 29.7417
R3020 standby_ip.n18 standby_ip.n17 29.7417
R3021 standby_ip.n13 standby_ip.n6 16.7534
R3022 standby_ip.n0 standby_ip.n14 16.7534
R3023 standby_ip.n1 standby_ip 13.0593
R3024 standby_ip.n21 standby_ip.n6 12.9887
R3025 standby_ip.n0 standby_ip.n22 12.9887
R3026 standby_ip standby_ip.t10 12.6603
R3027 standby_ip standby_ip.n26 9.27339
R3028 standby_ip.n25 standby_ip.n23 5.53161
R3029 standby_ip.n26 standby_ip.n2 5.46183
R3030 standby_ip standby_ip.n1 5.4255
R3031 standby_ip.n25 standby_ip.n24 4.67076
R3032 standby_ip.n3 standby_ip 1.88798
R3033 standby_ip standby_ip.n25 3.51723
R3034 standby_ip.n2 standby_ip 2.98717
R3035 standby_ip.n1 standby_ip.n6 2.80971
R3036 standby_ip.n26 standby_ip 2.78266
R3037 standby_ip.n5 standby_ip 2.74336
R3038 standby_ip.n1 standby_ip.n0 2.49791
R3039 a_2971_n1521.t1 a_2971_n1521.n1 405.735
R3040 a_2971_n1521.n1 a_2971_n1521.t0 294.611
R3041 a_2971_n1521.n0 a_2971_n1521.t3 254.389
R3042 a_2971_n1521.n0 a_2971_n1521.t2 211.01
R3043 a_2971_n1521.n1 a_2971_n1521.n0 152
R3044 a_14035_n1997.t0 a_14035_n1997.t1 38.7697
R3045 a_2132_n17582.t0 a_2132_n17582.t1 83.9053
R3046 a_18932_n17416.t0 a_18932_n17416.t1 83.5579
R3047 avss.n20 avss.n19 18580.7
R3048 avss.n38 avss.n37 15308.7
R3049 avss.n76 avss.n20 12246.6
R3050 avss.n40 avss.n35 3599.36
R3051 avss.n41 avss.n35 3599.36
R3052 avss.n41 avss.n34 3599.36
R3053 avss.n40 avss.n34 3599.36
R3054 avss.n67 avss.n25 2489.59
R3055 avss.n67 avss.n26 2489.59
R3056 avss.n69 avss.n26 2489.59
R3057 avss.n69 avss.n25 2489.59
R3058 avss.n28 avss.n21 2489.59
R3059 avss.n28 avss.n22 2489.59
R3060 avss.n74 avss.n22 2489.59
R3061 avss.n74 avss.n21 2489.59
R3062 avss.n78 avss.n13 2489.59
R3063 avss.n78 avss.n14 2489.59
R3064 avss.n16 avss.n14 2489.59
R3065 avss.n16 avss.n13 2489.59
R3066 avss.n88 avss.n6 2489.59
R3067 avss.n90 avss.n6 2489.59
R3068 avss.n90 avss.n5 2489.59
R3069 avss.n88 avss.n5 2489.59
R3070 avss.n36 avss.n20 2342.14
R3071 avss.n77 avss.n76 930.542
R3072 avss.n76 avss.n75 930.542
R3073 avss.n43 avss.n42 881.42
R3074 avss.n19 avss.t18 633.244
R3075 avss.n15 avss.t16 633.244
R3076 avss.t12 avss.n17 633.244
R3077 avss.n77 avss.t14 633.244
R3078 avss.n75 avss.t8 633.244
R3079 avss.n29 avss.t10 633.244
R3080 avss.t20 avss.n30 633.244
R3081 avss.n37 avss.t22 633.244
R3082 avss.t4 avss.n36 412.863
R3083 avss.t0 avss.n38 397.358
R3084 avss.n17 avss.n15 362.704
R3085 avss.n30 avss.n29 362.704
R3086 avss.t6 avss.t4 306.255
R3087 avss.t2 avss.t6 306.255
R3088 avss.t2 avss.t24 306.255
R3089 avss.t24 avss.t0 306.255
R3090 avss.n39 avss.n32 295.807
R3091 avss.n66 avss.n65 289.13
R3092 avss.n87 avss.n3 289.13
R3093 avss.n92 avss.n91 288.753
R3094 avss.n70 avss.n24 288.753
R3095 avss.n89 avss.t18 234.865
R3096 avss.n89 avss.t16 234.865
R3097 avss.n18 avss.t12 234.865
R3098 avss.t14 avss.n18 234.865
R3099 avss.n27 avss.t8 234.865
R3100 avss.t10 avss.n27 234.865
R3101 avss.n68 avss.t20 234.865
R3102 avss.n68 avss.t22 234.865
R3103 avss.n31 avss.n10 152.73
R3104 avss.n73 avss.n72 152.73
R3105 avss.n80 avss.n7 152.73
R3106 avss.n79 avss.n12 152.73
R3107 avss.n39 avss.n33 118.081
R3108 avss.n91 avss.n4 103.529
R3109 avss.n64 avss.n31 103.529
R3110 avss.n72 avss.n71 103.529
R3111 avss.n66 avss.n64 103.529
R3112 avss.n71 avss.n70 103.529
R3113 avss.n86 avss.n7 103.529
R3114 avss.n12 avss.n4 103.529
R3115 avss.n87 avss.n86 103.529
R3116 avss.n88 avss.n87 97.5005
R3117 avss.n89 avss.n88 97.5005
R3118 avss.n91 avss.n90 97.5005
R3119 avss.n90 avss.n89 97.5005
R3120 avss.n13 avss.n7 97.5005
R3121 avss.n18 avss.n13 97.5005
R3122 avss.n14 avss.n12 97.5005
R3123 avss.n18 avss.n14 97.5005
R3124 avss.n31 avss.n21 97.5005
R3125 avss.n27 avss.n21 97.5005
R3126 avss.n72 avss.n22 97.5005
R3127 avss.n27 avss.n22 97.5005
R3128 avss.n70 avss.n69 97.5005
R3129 avss.n69 avss.n68 97.5005
R3130 avss.n67 avss.n66 97.5005
R3131 avss.n68 avss.n67 97.5005
R3132 avss.n42 avss.n33 69.8003
R3133 avss.n38 avss.n35 54.5071
R3134 avss.n5 avss.n3 48.7505
R3135 avss.n19 avss.n5 48.7505
R3136 avss.n8 avss.n6 48.7505
R3137 avss.n15 avss.n6 48.7505
R3138 avss.n16 avss.n8 48.7505
R3139 avss.n17 avss.n16 48.7505
R3140 avss.n79 avss.n78 48.7505
R3141 avss.n78 avss.n77 48.7505
R3142 avss.n74 avss.n73 48.7505
R3143 avss.n75 avss.n74 48.7505
R3144 avss.n28 avss.n23 48.7505
R3145 avss.n29 avss.n28 48.7505
R3146 avss.n25 avss.n23 48.7505
R3147 avss.n30 avss.n25 48.7505
R3148 avss.n65 avss.n26 48.7505
R3149 avss.n37 avss.n26 48.7505
R3150 avss.n40 avss.n39 45.0005
R3151 avss.t2 avss.n40 45.0005
R3152 avss.n42 avss.n41 45.0005
R3153 avss.n41 avss.t2 45.0005
R3154 avss.n64 avss.n63 40.3697
R3155 avss.n71 avss.n23 40.3697
R3156 avss.n86 avss.n85 40.3697
R3157 avss.n8 avss.n4 40.3697
R3158 avss.n94 avss.n1 39.7977
R3159 avss.n34 avss.n33 39.0005
R3160 avss.n36 avss.n34 39.0005
R3161 avss.n35 avss.n32 39.0005
R3162 avss.n94 avss 33.7505
R3163 avss.n84 avss.t13 29.9199
R3164 avss.n62 avss.t21 29.9199
R3165 avss.n62 avss.t11 29.9199
R3166 avss.n84 avss.t17 29.9199
R3167 avss.n2 avss.t19 29.798
R3168 avss.n57 avss.t23 29.798
R3169 avss.n11 avss.t15 29.798
R3170 avss.n11 avss.t9 29.798
R3171 avss.n32 avss.t1 20.9512
R3172 avss.n46 avss.n45 18.8362
R3173 avss.n46 avss.n44 18.6458
R3174 avss.n44 avss.t3 4.133
R3175 avss.n44 avss.t25 4.133
R3176 avss.n45 avss.t5 4.133
R3177 avss.n45 avss.t7 4.133
R3178 avss.n47 avss.n43 1.61679
R3179 avss.n55 avss 1.33946
R3180 avss.n58 avss.n24 1.21803
R3181 avss.n93 avss.n92 1.21803
R3182 avss.n54 avss.n47 0.8655
R3183 avss.n63 avss.n62 0.664786
R3184 avss.n81 avss.n10 0.664786
R3185 avss.n81 avss.n80 0.664786
R3186 avss.n85 avss.n84 0.664786
R3187 avss.n55 avss.n54 0.53175
R3188 avss.n56 avss.n9 0.434977
R3189 avss.n95 avss.n0 0.433066
R3190 avss.n61 avss.n59 0.433066
R3191 avss.n61 avss.n60 0.433066
R3192 avss.n60 avss.n0 0.433066
R3193 avss.n65 avss.n24 0.376971
R3194 avss.n92 avss.n3 0.376971
R3195 avss.n84 avss.n0 0.299413
R3196 avss.n62 avss.n61 0.299413
R3197 avss.n62 avss.n9 0.247783
R3198 avss.n84 avss.n83 0.247783
R3199 avss.n83 avss 0.245943
R3200 avss.n59 avss.n58 0.231236
R3201 avss.n82 avss.n9 0.201672
R3202 avss.n83 avss.n82 0.201672
R3203 avss.n2 avss.n1 0.2005
R3204 avss.n95 avss.n94 0.2005
R3205 avss.n47 avss.n46 0.1855
R3206 avss.n49 avss.n48 0.122162
R3207 avss.n82 avss.n81 0.120904
R3208 avss.n50 avss.n49 0.105544
R3209 avss.n51 avss.n50 0.101695
R3210 avss.n73 avss.n10 0.1005
R3211 avss.n80 avss.n79 0.1005
R3212 avss.n60 avss.n11 0.0997647
R3213 avss.n53 avss.n48 0.0989292
R3214 avss.n56 avss.n55 0.096886
R3215 avss.n54 avss.n53 0.0847138
R3216 avss.n63 avss.n23 0.0825513
R3217 avss.n85 avss.n8 0.0825513
R3218 avss.n51 avss.n48 0.0586846
R3219 avss.n57 avss.n56 0.0480171
R3220 avss avss.n95 0.0332586
R3221 avss.n59 avss 0.0330342
R3222 avss.n94 avss.n93 0.0328276
R3223 avss.n43 avss.n32 0.0328232
R3224 avss.n53 avss.n52 0.0277801
R3225 avss.n50 avss.t28 0.0083125
R3226 avss.n49 avss.t29 0.0083125
R3227 avss.n48 avss.t26 0.0083125
R3228 avss.n52 avss.t27 0.0083125
R3229 avss avss.n1 0.00342969
R3230 avss.n93 avss.n2 0.000931034
R3231 avss.n58 avss.n57 0.000928082
R3232 avss.n81 avss.n11 0.000683824
R3233 avss.n52 avss.n51 0.000622332
R3234 avdd.n92 avdd.n91 15807.9
R3235 avdd.n93 avdd.n92 15807.9
R3236 avdd.n93 avdd.n28 15807.9
R3237 avdd.n91 avdd.n28 15807.9
R3238 avdd.n90 avdd.n27 8112.97
R3239 avdd.n94 avdd.n27 8112.97
R3240 avdd.n94 avdd.n26 8112.97
R3241 avdd.n90 avdd.n26 8112.97
R3242 avdd.n98 avdd.n6 2166
R3243 avdd.n97 avdd.n6 2166
R3244 avdd.n98 avdd.n7 2166
R3245 avdd.n97 avdd.n7 2166
R3246 avdd.n78 avdd.n77 1643.17
R3247 avdd.n77 avdd.n76 1643.17
R3248 avdd.n74 avdd.n69 1643.17
R3249 avdd.n80 avdd.n69 1643.17
R3250 avdd.n52 avdd.n37 1643.17
R3251 avdd.n60 avdd.n37 1643.17
R3252 avdd.n55 avdd.n54 1643.17
R3253 avdd.n58 avdd.n55 1643.17
R3254 avdd.n89 avdd.n88 1439.4
R3255 avdd.n89 avdd.n29 1352.37
R3256 avdd.n66 avdd.n25 1313.54
R3257 avdd.n71 avdd.n70 1106.59
R3258 avdd.n70 avdd.n68 1106.59
R3259 avdd.n40 avdd.n39 1106.59
R3260 avdd.n39 avdd.n36 1106.59
R3261 avdd.n78 avdd.n68 536.587
R3262 avdd.n76 avdd.n71 536.587
R3263 avdd.n74 avdd.n71 536.587
R3264 avdd.n80 avdd.n68 536.587
R3265 avdd.n52 avdd.n40 536.587
R3266 avdd.n54 avdd.n40 536.587
R3267 avdd.n58 avdd.n36 536.587
R3268 avdd.n60 avdd.n36 536.587
R3269 avdd.n75 avdd.t7 382.582
R3270 avdd.n79 avdd.t7 382.582
R3271 avdd.n53 avdd.t0 382.582
R3272 avdd.n59 avdd.t0 382.582
R3273 avdd.n73 avdd.n30 319.248
R3274 avdd.n57 avdd.n56 319.248
R3275 avdd.n88 avdd.n31 287.265
R3276 avdd.n38 avdd.n29 287.265
R3277 avdd.n88 avdd.n30 276.295
R3278 avdd.n56 avdd.n29 276.295
R3279 avdd.n86 avdd.t8 227.377
R3280 avdd.n1 avdd.t19 227.377
R3281 avdd.n34 avdd.t2 227.377
R3282 avdd.n43 avdd.t1 227.377
R3283 avdd.n66 avdd.n3 205.554
R3284 avdd.n72 avdd.n31 189.742
R3285 avdd.n38 avdd.n35 189.742
R3286 avdd.n101 avdd.n3 186.73
R3287 avdd.t17 avdd.n6 157.492
R3288 avdd.t5 avdd.n7 157.492
R3289 avdd.n25 avdd.n4 118.862
R3290 avdd.n100 avdd.n4 115.031
R3291 avdd.n73 avdd.n72 108.569
R3292 avdd.n57 avdd.n35 108.569
R3293 avdd.t3 avdd.t17 107.677
R3294 avdd.t11 avdd.t3 107.677
R3295 avdd.t11 avdd.t9 107.677
R3296 avdd.t9 avdd.t5 107.677
R3297 avdd.n62 avdd.n5 63.4672
R3298 avdd.n23 avdd.t18 60.1061
R3299 avdd.n21 avdd.n20 54.9038
R3300 avdd.n21 avdd.n19 54.9038
R3301 avdd.n72 avdd.n2 32.2138
R3302 avdd.n61 avdd.n35 32.2138
R3303 avdd.n101 avdd.n100 31.7005
R3304 avdd.n102 avdd.n101 30.3938
R3305 avdd.n76 avdd.n73 26.4291
R3306 avdd.n76 avdd.n75 26.4291
R3307 avdd.n74 avdd.n2 26.4291
R3308 avdd.n75 avdd.n74 26.4291
R3309 avdd.n78 avdd.n32 26.4291
R3310 avdd.n79 avdd.n78 26.4291
R3311 avdd.n81 avdd.n80 26.4291
R3312 avdd.n80 avdd.n79 26.4291
R3313 avdd.n58 avdd.n57 26.4291
R3314 avdd.n59 avdd.n58 26.4291
R3315 avdd.n61 avdd.n60 26.4291
R3316 avdd.n60 avdd.n59 26.4291
R3317 avdd.n54 avdd.n41 26.4291
R3318 avdd.n54 avdd.n53 26.4291
R3319 avdd.n52 avdd.n51 26.4291
R3320 avdd.n53 avdd.n52 26.4291
R3321 avdd.n96 avdd.n24 15.6997
R3322 avdd.n97 avdd.n96 14.2313
R3323 avdd.t11 avdd.n97 14.2313
R3324 avdd.n99 avdd.n98 14.2313
R3325 avdd.n98 avdd.t11 14.2313
R3326 avdd.n77 avdd.n30 13.2148
R3327 avdd.n77 avdd.t7 13.2148
R3328 avdd.n70 avdd.n31 13.2148
R3329 avdd.n70 avdd.t7 13.2148
R3330 avdd.n69 avdd.n3 13.2148
R3331 avdd.t7 avdd.n69 13.2148
R3332 avdd.n39 avdd.n38 13.2148
R3333 avdd.n39 avdd.t0 13.2148
R3334 avdd.n56 avdd.n55 13.2148
R3335 avdd.n55 avdd.t0 13.2148
R3336 avdd.n49 avdd.n37 13.2148
R3337 avdd.t0 avdd.n37 13.2148
R3338 avdd.n7 avdd.n4 12.3338
R3339 avdd.n47 avdd.n6 12.3338
R3340 avdd.n100 avdd.n99 8.13132
R3341 avdd.n95 avdd.n25 7.54184
R3342 avdd.n82 avdd.n32 7.30037
R3343 avdd.n46 avdd.n41 7.22016
R3344 avdd.n20 avdd.t4 6.92425
R3345 avdd.n20 avdd.t12 6.92425
R3346 avdd.n19 avdd.t10 6.92425
R3347 avdd.n19 avdd.t6 6.92425
R3348 avdd.n48 avdd.n47 6.88003
R3349 avdd.n99 avdd.n5 6.16704
R3350 avdd.n67 avdd.n66 3.51587
R3351 avdd.n50 avdd.n49 3.30818
R3352 avdd.n82 avdd.n81 2.8599
R3353 avdd.n90 avdd.n89 2.84665
R3354 avdd.n91 avdd.n90 2.84665
R3355 avdd.n95 avdd.n94 2.84665
R3356 avdd.n94 avdd.n93 2.84665
R3357 avdd.n51 avdd.n46 2.78239
R3358 avdd.n48 avdd.n5 2.51338
R3359 avdd.n49 avdd.n48 2.33395
R3360 avdd.n67 avdd.n27 2.28445
R3361 avdd.n92 avdd.n27 2.28445
R3362 avdd.n50 avdd.n26 2.28445
R3363 avdd.n28 avdd.n26 2.28445
R3364 avdd.n84 avdd 1.89829
R3365 avdd.n23 avdd.n22 1.87575
R3366 avdd.n102 avdd.n2 1.70717
R3367 avdd.n62 avdd.n61 1.70717
R3368 avdd.n81 avdd.n67 1.56476
R3369 avdd.n51 avdd.n50 1.54047
R3370 avdd.n85 avdd.n1 1.11161
R3371 avdd.n96 avdd.n95 1.03878
R3372 avdd.n65 avdd.n33 0.909856
R3373 avdd.n87 avdd.n65 0.871595
R3374 avdd.n42 avdd.n29 0.517167
R3375 avdd.n63 avdd.n62 0.517167
R3376 avdd.n103 avdd.n102 0.517167
R3377 avdd.n88 avdd.n87 0.517167
R3378 avdd.n83 avdd.n1 0.457832
R3379 avdd.n88 avdd.n32 0.30326
R3380 avdd.n41 avdd.n29 0.29856
R3381 avdd.n44 avdd.n34 0.277965
R3382 avdd.n44 avdd.n43 0.242141
R3383 avdd.n13 avdd.n12 0.221624
R3384 avdd.n45 avdd.n44 0.191202
R3385 avdd.n15 avdd.n8 0.171
R3386 avdd.n64 avdd 0.165618
R3387 avdd.n18 avdd.n8 0.158572
R3388 avdd.n45 avdd.n33 0.155105
R3389 avdd.n22 avdd.n18 0.129984
R3390 avdd.n65 avdd.n64 0.124867
R3391 avdd.n24 avdd.n23 0.0960224
R3392 avdd.n18 avdd.n17 0.0860931
R3393 avdd.n16 avdd.n15 0.0718577
R3394 avdd.n15 avdd.n14 0.0677409
R3395 avdd.n46 avdd.n45 0.058264
R3396 avdd.n83 avdd.n82 0.058264
R3397 avdd.n86 avdd.n85 0.0482015
R3398 avdd avdd.n63 0.0421667
R3399 avdd avdd.n0 0.035342
R3400 avdd.n12 avdd.n0 0.0293462
R3401 avdd.n22 avdd.n21 0.0285269
R3402 avdd.n17 avdd.n16 0.0255438
R3403 avdd.n14 avdd.n13 0.0253723
R3404 avdd.n12 avdd.n8 0.0246031
R3405 avdd.n85 avdd.n84 0.0240664
R3406 avdd.n11 avdd.t15 0.0122401
R3407 avdd avdd.n103 0.0122337
R3408 avdd.n17 avdd.t13 0.0122173
R3409 avdd.n10 avdd.t16 0.0113908
R3410 avdd.n9 avdd.t14 0.011362
R3411 avdd.n63 avdd.n34 0.0105575
R3412 avdd.n103 avdd.n1 0.0105575
R3413 avdd.n17 avdd.n9 0.00991802
R3414 avdd.n11 avdd.n10 0.00930403
R3415 avdd.n47 avdd.n24 0.00805162
R3416 avdd.n64 avdd 0.00600766
R3417 avdd.n43 avdd.n42 0.00573256
R3418 avdd.n42 avdd.n33 0.00515116
R3419 avdd.n87 avdd.n86 0.00333375
R3420 avdd.n14 avdd.n9 0.00220261
R3421 avdd.n16 avdd.n10 0.00176706
R3422 avdd.n84 avdd.n83 0.00111075
R3423 avdd.n64 avdd.n0 0.00109866
R3424 avdd.n13 avdd.n11 0.000671533
R3425 a_10620_n9666.t0 a_10620_n9666.t1 83.9243
R3426 a_20567_n1869.t1 a_20567_n1869.t0 198.571
R3427 a_20733_n1881.t0 a_20733_n1881.t1 60.0005
R3428 a_15539_n2791.n1 a_15539_n2791.t6 530.01
R3429 a_15539_n2791.t0 a_15539_n2791.n5 421.021
R3430 a_15539_n2791.n0 a_15539_n2791.t5 337.142
R3431 a_15539_n2791.n3 a_15539_n2791.t1 280.223
R3432 a_15539_n2791.n4 a_15539_n2791.t2 263.173
R3433 a_15539_n2791.n4 a_15539_n2791.t4 227.826
R3434 a_15539_n2791.n0 a_15539_n2791.t7 199.762
R3435 a_15539_n2791.n2 a_15539_n2791.n1 170.81
R3436 a_15539_n2791.n2 a_15539_n2791.n0 167.321
R3437 a_15539_n2791.n5 a_15539_n2791.n4 152
R3438 a_15539_n2791.n1 a_15539_n2791.t3 141.923
R3439 a_15539_n2791.n3 a_15539_n2791.n2 10.8376
R3440 a_15539_n2791.n5 a_15539_n2791.n3 2.50485
R3441 a_15705_n2791.t0 a_15705_n2791.n3 370.026
R3442 a_15705_n2791.n0 a_15705_n2791.t5 351.356
R3443 a_15705_n2791.n1 a_15705_n2791.t3 334.717
R3444 a_15705_n2791.n3 a_15705_n2791.t1 325.971
R3445 a_15705_n2791.n1 a_15705_n2791.t4 309.935
R3446 a_15705_n2791.n0 a_15705_n2791.t2 305.683
R3447 a_15705_n2791.n2 a_15705_n2791.n0 16.879
R3448 a_15705_n2791.n3 a_15705_n2791.n2 10.8867
R3449 a_15705_n2791.n2 a_15705_n2791.n1 9.3005
R3450 a_16782_n2425.t0 a_16782_n2425.t1 126.644
R3451 standby.n1 standby.t0 260.322
R3452 standby.n0 standby.t1 194.635
R3453 standby.n1 standby.t2 175.169
R3454 standby.n2 standby.n1 152
R3455 standby.n2 standby.n0 69.674
R3456 standby standby.n2 1.55726
R3457 standby.n0 standby 0.748625
R3458 a_4857_n1521.t0 a_4857_n1521.n1 405.735
R3459 a_4857_n1521.n1 a_4857_n1521.t1 294.611
R3460 a_4857_n1521.n0 a_4857_n1521.t2 254.389
R3461 a_4857_n1521.n0 a_4857_n1521.t3 211.01
R3462 a_4857_n1521.n1 a_4857_n1521.n0 152
R3463 x3.out_b.n5 x3.out_b.t8 397.163
R3464 x3.out_b.n3 x3.out_b.t4 397.163
R3465 x3.out_b.n6 x3.out_b.t8 396.286
R3466 x3.out_b.n4 x3.out_b.t4 396.286
R3467 x3.out_b.t3 x3.out_b.n5 375.649
R3468 x3.out_b.n6 x3.out_b.t3 375.649
R3469 x3.out_b.n0 x3.out_b.t6 375.649
R3470 x3.out_b.n7 x3.out_b.t6 375.649
R3471 x3.out_b.t7 x3.out_b.n3 375.649
R3472 x3.out_b.n4 x3.out_b.t7 375.649
R3473 x3.out_b.n2 x3.out_b.t0 227.887
R3474 x3.out_b.n2 x3.out_b.n8 25.0905
R3475 x3.out_b.n5 x3.out_b.n0 21.5154
R3476 x3.out_b.n3 x3.out_b.n0 21.1069
R3477 x3.out_b.n7 x3.out_b.n4 20.6372
R3478 x3.out_b.n7 x3.out_b.n6 20.6372
R3479 x3.out_b.n2 x3.out_b.t5 12.777
R3480 x3.out_b.n8 x3.out_b.t1 5.5105
R3481 x3.out_b.n8 x3.out_b.t2 5.5105
R3482 x3.out_b.n1 x3.out_b.n0 5.32901
R3483 x3.out_b.n1 x3.out_b.n7 2.74252
R3484 x3.out_b.n2 x3.out_b.n1 1.06508
R3485 a_19955_n2791.n1 a_19955_n2791.t4 530.01
R3486 a_19955_n2791.t1 a_19955_n2791.n5 421.021
R3487 a_19955_n2791.n0 a_19955_n2791.t3 337.142
R3488 a_19955_n2791.n3 a_19955_n2791.t0 280.223
R3489 a_19955_n2791.n4 a_19955_n2791.t6 263.173
R3490 a_19955_n2791.n4 a_19955_n2791.t2 227.826
R3491 a_19955_n2791.n0 a_19955_n2791.t5 199.762
R3492 a_19955_n2791.n2 a_19955_n2791.n1 170.81
R3493 a_19955_n2791.n2 a_19955_n2791.n0 167.321
R3494 a_19955_n2791.n5 a_19955_n2791.n4 152
R3495 a_19955_n2791.n1 a_19955_n2791.t7 141.923
R3496 a_19955_n2791.n3 a_19955_n2791.n2 10.8376
R3497 a_19955_n2791.n5 a_19955_n2791.n3 2.50485
R3498 a_20121_n2791.t0 a_20121_n2791.n3 370.026
R3499 a_20121_n2791.n0 a_20121_n2791.t4 351.356
R3500 a_20121_n2791.n1 a_20121_n2791.t3 334.717
R3501 a_20121_n2791.n3 a_20121_n2791.t1 325.971
R3502 a_20121_n2791.n1 a_20121_n2791.t2 309.935
R3503 a_20121_n2791.n0 a_20121_n2791.t5 305.683
R3504 a_20121_n2791.n2 a_20121_n2791.n0 16.879
R3505 a_20121_n2791.n3 a_20121_n2791.n2 10.8867
R3506 a_20121_n2791.n2 a_20121_n2791.n1 9.3005
R3507 a_19567_n2247.t1 a_19567_n2247.n1 386.31
R3508 a_19567_n2247.n1 a_19567_n2247.t0 249.956
R3509 a_19567_n2247.n0 a_19567_n2247.t3 239.04
R3510 a_19567_n2247.n1 a_19567_n2247.n0 175.661
R3511 a_19567_n2247.n0 a_19567_n2247.t2 166.739
R3512 ena.n0 ena.t2 260.322
R3513 ena.n2 ena.t0 194.63
R3514 ena.n0 ena.t1 175.169
R3515 ena.n1 ena.n0 152
R3516 ena.n3 ena.n2 51.6747
R3517 ena ena.n3 4.94983
R3518 ena.n3 ena.n1 3.45996
R3519 ena.n1 ena 1.55726
R3520 ena.n2 ena 0.746125
R3521 a_19003_n2817.n6 a_19003_n2817.n5 746.659
R3522 a_19003_n2817.n0 a_19003_n2817.t5 389.183
R3523 a_19003_n2817.n2 a_19003_n2817.t3 256.988
R3524 a_19003_n2817.n1 a_19003_n2817.n0 251.167
R3525 a_19003_n2817.n1 a_19003_n2817.t1 223.571
R3526 a_19003_n2817.n4 a_19003_n2817.t8 212.081
R3527 a_19003_n2817.n5 a_19003_n2817.n4 181.942
R3528 a_19003_n2817.n0 a_19003_n2817.t4 174.891
R3529 a_19003_n2817.n2 a_19003_n2817.t6 163.803
R3530 a_19003_n2817.n3 a_19003_n2817.t7 139.78
R3531 a_19003_n2817.n3 a_19003_n2817.n2 129.264
R3532 a_19003_n2817.n6 a_19003_n2817.t2 63.3219
R3533 a_19003_n2817.t0 a_19003_n2817.n6 63.3219
R3534 a_19003_n2817.n5 a_19003_n2817.n1 24.6993
R3535 a_19003_n2817.n4 a_19003_n2817.n3 22.6399
R3536 a_19567_n2791.t0 a_19567_n2791.n1 386.31
R3537 a_19567_n2791.n1 a_19567_n2791.t1 249.956
R3538 a_19567_n2791.n0 a_19567_n2791.t3 239.04
R3539 a_19567_n2791.n1 a_19567_n2791.n0 175.661
R3540 a_19567_n2791.n0 a_19567_n2791.t2 166.739
R3541 vg1.n10 vg1.t0 85.228
R3542 vg1.n0 vg1.t3 61.1305
R3543 vg1.n7 vg1.t5 54.828
R3544 vg1.n7 vg1.t0 54.828
R3545 vg1.n5 vg1.t2 42.6599
R3546 vg1.n8 vg1.n7 32.9015
R3547 vg1.n10 vg1.n9 30.9745
R3548 vg1.n9 vg1.t1 20.9512
R3549 vg1.n6 vg1.n5 3.63479
R3550 vg1.n11 vg1.n10 2.3255
R3551 vg1.n12 vg1.n0 0.471594
R3552 vg1.n5 vg1.n4 0.390524
R3553 vg1.n9 vg1.n8 0.238607
R3554 vg1.n11 vg1.n6 0.176742
R3555 vg1 vg1.n12 0.133236
R3556 vg1.n1 vg1.t9 0.0767969
R3557 vg1.n2 vg1.n1 0.0752537
R3558 vg1.n3 vg1.n2 0.0752537
R3559 vg1.n4 vg1.t8 0.0717511
R3560 vg1.n0 vg1 0.0387813
R3561 vg1.n12 vg1.n11 0.0257152
R3562 vg1.n8 vg1.n6 0.0123355
R3563 vg1.n4 vg1.n3 0.00554581
R3564 vg1.n1 vg1.t4 0.00204321
R3565 vg1.n2 vg1.t7 0.00204321
R3566 vg1.n3 vg1.t6 0.00204321
R3567 a_21145_n1869.n0 a_21145_n1869.t1 68.3338
R3568 a_21145_n1869.n0 a_21145_n1869.t0 26.3935
R3569 a_21145_n1869.n1 a_21145_n1869.n0 14.4005
R3570 a_21211_n2817.n6 a_21211_n2817.n5 746.659
R3571 a_21211_n2817.n0 a_21211_n2817.t8 389.183
R3572 a_21211_n2817.n2 a_21211_n2817.t6 256.988
R3573 a_21211_n2817.n1 a_21211_n2817.n0 251.167
R3574 a_21211_n2817.n1 a_21211_n2817.t1 223.571
R3575 a_21211_n2817.n4 a_21211_n2817.t5 212.081
R3576 a_21211_n2817.n5 a_21211_n2817.n4 181.942
R3577 a_21211_n2817.n0 a_21211_n2817.t7 174.891
R3578 a_21211_n2817.n2 a_21211_n2817.t3 163.803
R3579 a_21211_n2817.n3 a_21211_n2817.t4 139.78
R3580 a_21211_n2817.n3 a_21211_n2817.n2 129.264
R3581 a_21211_n2817.n6 a_21211_n2817.t2 63.3219
R3582 a_21211_n2817.t0 a_21211_n2817.n6 63.3219
R3583 a_21211_n2817.n5 a_21211_n2817.n1 24.6993
R3584 a_21211_n2817.n4 a_21211_n2817.n3 22.6399
R3585 xin.n36 xin.t8 594.832
R3586 xin.t18 xin.n5 380.808
R3587 xin.n6 xin.t18 380.808
R3588 xin.n6 xin.t15 380.611
R3589 xin.t15 xin.n5 380.611
R3590 xin.t13 xin.n7 380.611
R3591 xin.n8 xin.t13 380.611
R3592 xin.t19 xin.n4 380.611
R3593 xin.n9 xin.t19 380.611
R3594 xin.n11 xin.t16 380.611
R3595 xin.t16 xin.n10 380.611
R3596 xin.n12 xin.t11 380.611
R3597 xin.t11 xin.n3 380.611
R3598 xin.t10 xin.n13 380.611
R3599 xin.n14 xin.t10 380.611
R3600 xin.t17 xin.n2 380.611
R3601 xin.n15 xin.t17 380.611
R3602 xin.n17 xin.t14 380.611
R3603 xin.t14 xin.n16 380.611
R3604 xin.n18 xin.t12 380.611
R3605 xin.t12 xin.n1 380.611
R3606 xin.t9 xin.n19 380.611
R3607 xin.n20 xin.t9 380.611
R3608 xin.n21 xin.t6 380.611
R3609 xin.t6 xin.n0 380.611
R3610 xin.n36 xin.t21 194.639
R3611 xin.n25 xin.t20 124.457
R3612 xin.n25 xin.t7 106.793
R3613 xin.t7 xin.n23 86.3125
R3614 xin.t20 xin.n24 86.3125
R3615 xin.n24 xin.n23 58.6245
R3616 xin.n30 xin.t5 45.927
R3617 xin.n28 xin.n27 20.1298
R3618 xin.n27 xin.n23 12.2455
R3619 xin.n35 xin.n34 4.04311
R3620 xin.n26 xin.n24 3.56553
R3621 xin.n34 xin.n29 3.51336
R3622 xin.n30 xin.n29 3.51061
R3623 xin.n28 xin.n22 1.95915
R3624 xin.n35 xin.n28 1.1106
R3625 xin.n22 xin.n21 0.8105
R3626 xin.n22 xin.n0 0.7905
R3627 xin.n27 xin.n26 0.741791
R3628 xin.n26 xin.n25 0.715885
R3629 xin.n36 xin.n35 0.4755
R3630 xin xin.n36 0.377063
R3631 xin.n8 xin.n5 0.198
R3632 xin.n9 xin.n8 0.198
R3633 xin.n10 xin.n9 0.198
R3634 xin.n10 xin.n3 0.198
R3635 xin.n14 xin.n3 0.198
R3636 xin.n15 xin.n14 0.198
R3637 xin.n16 xin.n15 0.198
R3638 xin.n16 xin.n1 0.198
R3639 xin.n20 xin.n1 0.198
R3640 xin.n21 xin.n20 0.198
R3641 xin.n7 xin.n6 0.198
R3642 xin.n7 xin.n4 0.198
R3643 xin.n11 xin.n4 0.198
R3644 xin.n12 xin.n11 0.198
R3645 xin.n13 xin.n12 0.198
R3646 xin.n13 xin.n2 0.198
R3647 xin.n17 xin.n2 0.198
R3648 xin.n18 xin.n17 0.198
R3649 xin.n19 xin.n18 0.198
R3650 xin.n19 xin.n0 0.198
R3651 xin.t3 xin.t1 0.0760058
R3652 xin.n31 xin.n30 0.0410952
R3653 xin.n32 xin.n29 0.0410952
R3654 xin.n34 xin.n33 0.0410952
R3655 xin.n32 xin.t4 0.0264927
R3656 xin.n31 xin.t0 0.0264885
R3657 xin.n33 xin.t3 0.0264703
R3658 xin.n33 xin.t2 0.0264296
R3659 xin.t2 xin.n32 0.0264114
R3660 xin.t4 xin.n31 0.0264072
R3661 a_19182_n2791.t0 a_19182_n2791.t1 87.1434
R3662 a_2132_n17250.t0 a_2132_n17250.t1 82.3314
R3663 a_24220_n9500.t0 a_24220_n9500.t1 83.56
R3664 a_17913_n2241.t0 a_17913_n2241.n3 370.026
R3665 a_17913_n2241.n0 a_17913_n2241.t3 351.356
R3666 a_17913_n2241.n1 a_17913_n2241.t2 334.717
R3667 a_17913_n2241.n3 a_17913_n2241.t1 325.971
R3668 a_17913_n2241.n1 a_17913_n2241.t4 309.935
R3669 a_17913_n2241.n0 a_17913_n2241.t5 305.683
R3670 a_17913_n2241.n2 a_17913_n2241.n0 16.879
R3671 a_17913_n2241.n3 a_17913_n2241.n2 10.8867
R3672 a_17913_n2241.n2 a_17913_n2241.n1 9.3005
R3673 a_18263_n1869.n3 a_18263_n1869.n2 674.338
R3674 a_18263_n1869.n1 a_18263_n1869.t4 332.58
R3675 a_18263_n1869.n2 a_18263_n1869.n0 284.012
R3676 a_18263_n1869.n2 a_18263_n1869.n1 253.648
R3677 a_18263_n1869.n1 a_18263_n1869.t5 168.701
R3678 a_18263_n1869.n3 a_18263_n1869.t2 96.1553
R3679 a_18263_n1869.t1 a_18263_n1869.n3 65.6672
R3680 a_18263_n1869.n0 a_18263_n1869.t3 65.0005
R3681 a_18263_n1869.n0 a_18263_n1869.t0 45.0005
R3682 a_18359_n1869.t0 a_18359_n1869.t1 198.571
R3683 vg2.n2 vg2.t9 87.8852
R3684 vg2.n9 vg2.t5 87.8852
R3685 vg2.n5 vg2.t6 85.228
R3686 vg2.n12 vg2.t7 85.228
R3687 vg2.n15 vg2.t8 67.0783
R3688 vg2.n4 vg2.t9 54.828
R3689 vg2.t6 vg2.n4 54.828
R3690 vg2.n11 vg2.t5 54.828
R3691 vg2.t7 vg2.n11 54.828
R3692 vg2.n16 vg2.t0 42.6015
R3693 vg2.n4 vg2.n3 30.4005
R3694 vg2.n11 vg2.n10 30.4005
R3695 vg2.n3 vg2.n1 29.1205
R3696 vg2.n5 vg2.n1 29.1205
R3697 vg2.n10 vg2.n8 29.1205
R3698 vg2.n12 vg2.n8 29.1205
R3699 vg2.n6 vg2.n5 2.3255
R3700 vg2.n13 vg2.n12 2.3255
R3701 vg2.n3 vg2.n2 2.13477
R3702 vg2.n10 vg2.n9 2.13477
R3703 vg2 vg2.n14 0.742464
R3704 vg2.n16 vg2.n15 0.714193
R3705 vg2.n14 vg2.n6 0.474719
R3706 vg2.n14 vg2.n13 0.474719
R3707 vg2.n1 vg2.n0 0.423227
R3708 vg2.n8 vg2.n7 0.423227
R3709 vg2.n2 vg2.n0 0.308459
R3710 vg2.n9 vg2.n7 0.308459
R3711 vg2.n6 vg2.n0 0.284875
R3712 vg2.n13 vg2.n7 0.284875
R3713 vg2.n15 vg2.t3 0.170134
R3714 vg2 vg2.n16 0.119455
R3715 vg2.t1 vg2.t2 0.0652716
R3716 vg2.t4 vg2.t1 0.0652716
R3717 vg2.t3 vg2.t4 0.0652716
R3718 vrb.n2 vrb.t4 43.1048
R3719 vrb.n0 vrb.t3 22.3777
R3720 vrb.n1 vrb.t0 22.1989
R3721 vrb.n1 vrb.t2 21.3671
R3722 vrb.n0 vrb.t1 21.3663
R3723 vrb.n3 vrb.n2 1.11856
R3724 vrb.n3 vrb.n0 0.759192
R3725 vrb.n2 vrb.n1 0.758408
R3726 vrb vrb.n3 0.0491111
R3727 a_18359_n2791.t0 a_18359_n2791.t1 198.571
R3728 a_18525_n2791.t0 a_18525_n2791.t1 60.0005
R3729 a_2130_n20844.t0 a_2130_n20844.t1 82.0028
R3730 a_24530_n21010.t0 a_24530_n21010.t1 81.9478
R3731 a_15083_n2791.t0 a_15083_n2791.t1 60.0005
R3732 a_18932_n15424.t0 a_18932_n15424.t1 83.5579
R3733 a_14285_n2281.n1 a_14285_n2281.n0 953.039
R3734 a_14285_n2281.n0 a_14285_n2281.t3 33.4905
R3735 a_14285_n2281.n0 a_14285_n2281.t2 31.5205
R3736 a_14285_n2281.t0 a_14285_n2281.n1 26.5955
R3737 a_14285_n2281.n1 a_14285_n2281.t1 26.5955
R3738 a_14285_n2079.n0 a_14285_n2079.t1 1201.3
R3739 a_14285_n2079.n0 a_14285_n2079.t2 26.5955
R3740 a_14285_n2079.t0 a_14285_n2079.n0 26.5955
R3741 a_18828_n1869.n3 a_18828_n1869.n2 636.953
R3742 a_18828_n1869.n1 a_18828_n1869.t4 366.856
R3743 a_18828_n1869.n2 a_18828_n1869.n0 300.2
R3744 a_18828_n1869.n2 a_18828_n1869.n1 225.036
R3745 a_18828_n1869.n1 a_18828_n1869.t5 174.056
R3746 a_18828_n1869.n0 a_18828_n1869.t2 70.0005
R3747 a_18828_n1869.t1 a_18828_n1869.n3 68.0124
R3748 a_18828_n1869.n3 a_18828_n1869.t3 63.3219
R3749 a_18828_n1869.n0 a_18828_n1869.t0 61.6672
R3750 a_19182_n1881.t0 a_19182_n1881.t1 87.1434
R3751 a_19003_n1943.n5 a_19003_n1943.n1 746.659
R3752 a_19003_n1943.n0 a_19003_n1943.t8 389.183
R3753 a_19003_n1943.n2 a_19003_n1943.t5 256.988
R3754 a_19003_n1943.n6 a_19003_n1943.n0 251.167
R3755 a_19003_n1943.t0 a_19003_n1943.n6 223.571
R3756 a_19003_n1943.n4 a_19003_n1943.t7 212.081
R3757 a_19003_n1943.n5 a_19003_n1943.n4 181.942
R3758 a_19003_n1943.n0 a_19003_n1943.t3 174.891
R3759 a_19003_n1943.n2 a_19003_n1943.t6 163.803
R3760 a_19003_n1943.n3 a_19003_n1943.t4 139.78
R3761 a_19003_n1943.n3 a_19003_n1943.n2 129.264
R3762 a_19003_n1943.n1 a_19003_n1943.t1 63.3219
R3763 a_19003_n1943.n1 a_19003_n1943.t2 63.3219
R3764 a_19003_n1943.n6 a_19003_n1943.n5 24.6993
R3765 a_19003_n1943.n4 a_19003_n1943.n3 22.6399
R3766 vn.t9 vn.n3 182.935
R3767 vn.t0 vn.n0 144.126
R3768 vn.n8 vn.n5 97.2442
R3769 vn.n9 vn.n3 97.2442
R3770 vn.n4 vn.t9 88.2031
R3771 vn.t8 vn.n3 85.228
R3772 vn.n5 vn.t8 85.228
R3773 vn.n9 vn.t3 85.228
R3774 vn.t3 vn.n8 85.228
R3775 vn.n1 vn.t0 85.228
R3776 vn vn.t6 64.2147
R3777 vn.n7 vn.n1 58.8987
R3778 vn vn.n2 56.3112
R3779 vn vn.t2 21.1687
R3780 vn.n8 vn.n7 17.975
R3781 vn.n9 vn.n0 17.975
R3782 vn vn.n6 16.8187
R3783 vn.n2 vn.t7 6.92425
R3784 vn.n2 vn.t5 6.92425
R3785 vn.n6 vn.t4 4.3505
R3786 vn.n6 vn.t1 4.3505
R3787 vn.n4 vn 3.29454
R3788 vn vn.n1 2.80102
R3789 vn.n8 vn 2.44682
R3790 vn.n3 vn 2.3255
R3791 vn vn.n9 2.3255
R3792 vn.n5 vn.n4 2.20282
R3793 vn.n7 vn 2.69718
R3794 vn vn.n0 2.67028
R3795 a_10620_n7674.t0 a_10620_n7674.t1 82.5973
R3796 a_24220_n7840.t0 a_24220_n7840.t1 83.56
R3797 x7.x2.Qb1.n4 x7.x2.Qb1.t1 372.361
R3798 x7.x2.Qb1.n2 x7.x2.Qb1.t5 333.651
R3799 x7.x2.Qb1.n2 x7.x2.Qb1.t2 297.233
R3800 x7.x2.Qb1.n1 x7.x2.Qb1.t3 294.557
R3801 x7.x2.Qb1.n5 x7.x2.Qb1.t0 231.921
R3802 x7.x2.Qb1.n1 x7.x2.Qb1.t4 211.01
R3803 x7.x2.Qb1 x7.x2.Qb1.n2 195.701
R3804 x7.x2.Qb1.n0 x7.x2.Qb1.n1 152
R3805 x7.x2.Qb1.n5 x7.x2.Qb1.n0 40.9605
R3806 x7.x2.Qb1.n5 x7.x2.Qb1.n4 18.1966
R3807 x7.x2.Qb1.n0 x7.x2.Qb1 10.4234
R3808 x7.x2.Qb1.n4 x7.x2.Qb1.n3 9.35675
R3809 x7.x2.Qb1.n3 x7.x2.Qb1 6.49269
R3810 x7.x2.Qb1.n3 x7.x2.Qb1 3.52967
R3811 x7.x2.Qb1 x7.x2.Qb1.n5 2.5605
R3812 x7.x2.Qb1.n0 x7.x2.Qb1 2.01193
R3813 a_15960_n2791.n1 a_15960_n2791.n0 926.024
R3814 a_15960_n2791.t1 a_15960_n2791.n1 82.0838
R3815 a_15960_n2791.n0 a_15960_n2791.t0 63.3338
R3816 a_15960_n2791.n1 a_15960_n2791.t2 63.3219
R3817 a_15960_n2791.n0 a_15960_n2791.t3 29.7268
R3818 a_2130_n19516.t0 a_2130_n19516.t1 82.0028
R3819 a_24530_n19682.t0 a_24530_n19682.t1 81.9478
R3820 a_20579_n2247.t0 a_20579_n2247.n0 1327.82
R3821 a_20579_n2247.n0 a_20579_n2247.t2 194.655
R3822 a_20579_n2247.n0 a_20579_n2247.t1 63.3219
R3823 a_15083_n1881.t0 a_15083_n1881.t1 60.0005
R3824 a_18481_n2273.n3 a_18481_n2273.n2 647.119
R3825 a_18481_n2273.n1 a_18481_n2273.t4 350.253
R3826 a_18481_n2273.n2 a_18481_n2273.n0 260.339
R3827 a_18481_n2273.n2 a_18481_n2273.n1 246.119
R3828 a_18481_n2273.n1 a_18481_n2273.t5 189.588
R3829 a_18481_n2273.n3 a_18481_n2273.t0 89.1195
R3830 a_18481_n2273.n0 a_18481_n2273.t1 63.3338
R3831 a_18481_n2273.t2 a_18481_n2273.n3 41.0422
R3832 a_18481_n2273.n0 a_18481_n2273.t3 31.9797
R3833 a_18525_n1881.t0 a_18525_n1881.t1 60.0005
R3834 x7.x2.Qb2.n4 x7.x2.Qb2.t0 372.361
R3835 x7.x2.Qb2.n2 x7.x2.Qb2.t5 333.651
R3836 x7.x2.Qb2.n2 x7.x2.Qb2.t2 297.233
R3837 x7.x2.Qb2.n1 x7.x2.Qb2.t3 294.557
R3838 x7.x2.Qb2.n5 x7.x2.Qb2.t1 231.921
R3839 x7.x2.Qb2.n1 x7.x2.Qb2.t4 211.01
R3840 x7.x2.Qb2 x7.x2.Qb2.n2 195.701
R3841 x7.x2.Qb2.n0 x7.x2.Qb2.n1 152
R3842 x7.x2.Qb2.n5 x7.x2.Qb2.n0 40.9605
R3843 x7.x2.Qb2.n5 x7.x2.Qb2.n4 18.1966
R3844 x7.x2.Qb2.n0 x7.x2.Qb2 10.4234
R3845 x7.x2.Qb2.n4 x7.x2.Qb2.n3 9.36092
R3846 x7.x2.Qb2.n3 x7.x2.Qb2 6.49269
R3847 x7.x2.Qb2.n3 x7.x2.Qb2 3.52967
R3848 x7.x2.Qb2 x7.x2.Qb2.n5 2.5605
R3849 x7.x2.Qb2.n0 x7.x2.Qb2 2.01193
R3850 a_18168_n2791.n1 a_18168_n2791.n0 926.024
R3851 a_18168_n2791.n1 a_18168_n2791.t3 82.0838
R3852 a_18168_n2791.n0 a_18168_n2791.t0 63.3338
R3853 a_18168_n2791.t1 a_18168_n2791.n1 63.3219
R3854 a_18168_n2791.n0 a_18168_n2791.t2 29.7268
R3855 a_16055_n2791.n3 a_16055_n2791.n2 674.338
R3856 a_16055_n2791.n1 a_16055_n2791.t4 332.58
R3857 a_16055_n2791.n2 a_16055_n2791.n0 284.012
R3858 a_16055_n2791.n2 a_16055_n2791.n1 253.648
R3859 a_16055_n2791.n1 a_16055_n2791.t5 168.701
R3860 a_16055_n2791.t0 a_16055_n2791.n3 96.1553
R3861 a_16055_n2791.n3 a_16055_n2791.t2 65.6672
R3862 a_16055_n2791.n0 a_16055_n2791.t1 65.0005
R3863 a_16055_n2791.n0 a_16055_n2791.t3 45.0005
R3864 x7.x1.x4.Q x7.x1.x4.Q.t0 240.05
R3865 x7.x1.x4.Q x7.x1.x4.Q.t1 155.386
R3866 a_14009_n2404.t1 a_14009_n2404.n3 669.389
R3867 a_14009_n2404.n0 a_14009_n2404.t2 326.493
R3868 a_14009_n2404.n0 a_14009_n2404.t0 249.615
R3869 a_14009_n2404.n1 a_14009_n2404.t3 249.615
R3870 a_14009_n2404.n2 a_14009_n2404.t4 241.536
R3871 a_14009_n2404.n2 a_14009_n2404.t5 169.237
R3872 a_14009_n2404.n3 a_14009_n2404.n2 152
R3873 a_14009_n2404.n3 a_14009_n2404.n1 108.529
R3874 a_14009_n2404.n1 a_14009_n2404.n0 26.6245
R3875 a_24530_n20678.t0 a_24530_n20678.t1 81.9478
R3876 a_15539_n2241.n1 a_15539_n2241.t5 530.01
R3877 a_15539_n2241.t0 a_15539_n2241.n5 421.021
R3878 a_15539_n2241.n0 a_15539_n2241.t3 337.142
R3879 a_15539_n2241.n3 a_15539_n2241.t1 280.223
R3880 a_15539_n2241.n4 a_15539_n2241.t4 263.173
R3881 a_15539_n2241.n4 a_15539_n2241.t6 227.826
R3882 a_15539_n2241.n0 a_15539_n2241.t2 199.762
R3883 a_15539_n2241.n2 a_15539_n2241.n1 170.81
R3884 a_15539_n2241.n2 a_15539_n2241.n0 167.321
R3885 a_15539_n2241.n5 a_15539_n2241.n4 152
R3886 a_15539_n2241.n1 a_15539_n2241.t7 141.923
R3887 a_15539_n2241.n3 a_15539_n2241.n2 10.8376
R3888 a_15539_n2241.n5 a_15539_n2241.n3 2.50485
R3889 a_16729_n1869.n0 a_16729_n1869.t1 68.3338
R3890 a_16729_n1869.n0 a_16729_n1869.t0 26.3935
R3891 a_16729_n1869.n1 a_16729_n1869.n0 14.4005
R3892 a_16055_n1869.n3 a_16055_n1869.n2 674.338
R3893 a_16055_n1869.n1 a_16055_n1869.t4 332.58
R3894 a_16055_n1869.n2 a_16055_n1869.n0 284.012
R3895 a_16055_n1869.n2 a_16055_n1869.n1 253.648
R3896 a_16055_n1869.n1 a_16055_n1869.t5 168.701
R3897 a_16055_n1869.t1 a_16055_n1869.n3 96.1553
R3898 a_16055_n1869.n3 a_16055_n1869.t2 65.6672
R3899 a_16055_n1869.n0 a_16055_n1869.t0 65.0005
R3900 a_16055_n1869.n0 a_16055_n1869.t3 45.0005
R3901 a_2132_n15258.t0 a_2132_n15258.t1 83.9223
R3902 a_18990_n2425.t0 a_18990_n2425.t1 126.644
R3903 a_24530_n19350.t0 a_24530_n19350.t1 81.9478
R3904 a_16163_n2247.n0 a_16163_n2247.t1 1327.82
R3905 a_16163_n2247.t0 a_16163_n2247.n0 194.655
R3906 a_16163_n2247.n0 a_16163_n2247.t2 63.3219
R3907 a_2132_n16918.t0 a_2132_n16918.t1 82.3314
R3908 a_18932_n17084.t0 a_18932_n17084.t1 83.5579
R3909 a_10620_n9334.t0 a_10620_n9334.t1 83.9243
R3910 a_3134_n13324.t0 a_3134_n13324.t1 83.9223
R3911 x7.x1.x2.Q x7.x1.x2.Q.t0 240.05
R3912 x7.x1.x2.Q x7.x1.x2.Q.t1 155.386
R3913 a_18932_n17748.t0 a_18932_n17748.t1 83.5579
R3914 a_18937_n2791.t1 a_18937_n2791.t0 94.7268
R3915 x3.out.n3 x3.out.t6 393.144
R3916 x3.out.n5 x3.out.t7 393.144
R3917 x3.out.n4 x3.out.t6 391.815
R3918 x3.out.t7 x3.out.n2 391.815
R3919 x3.out.n5 x3.out.t4 371.31
R3920 x3.out.t4 x3.out.n2 371.31
R3921 x3.out.t3 x3.out.n1 371.31
R3922 x3.out.n6 x3.out.t3 371.31
R3923 x3.out.n4 x3.out.t8 371.31
R3924 x3.out.t8 x3.out.n3 371.31
R3925 x3.out.n0 x3.out.t0 227.886
R3926 x3.out.n0 x3.out.n9 25.0903
R3927 x3.out.n1 x3.out.n5 21.8335
R3928 x3.out.n3 x3.out.n1 21.6959
R3929 x3.out.n6 x3.out.n4 20.5053
R3930 x3.out.n7 x3.out.n2 19.6003
R3931 x3.out.n0 x3.out.t5 12.7763
R3932 x3.out.n9 x3.out.t1 5.5105
R3933 x3.out.n9 x3.out.t2 5.5105
R3934 x3.out.n8 x3.out.n1 5.0449
R3935 x3.out.n8 x3.out.n7 2.71826
R3936 x3.out.n7 x3.out.n6 0.90555
R3937 x3.out x3.out.n8 0.88175
R3938 x3.out x3.out.n0 0.794875
R3939 a_17359_n2247.t0 a_17359_n2247.n1 386.31
R3940 a_17359_n2247.n1 a_17359_n2247.t1 249.956
R3941 a_17359_n2247.n0 a_17359_n2247.t2 239.04
R3942 a_17359_n2247.n1 a_17359_n2247.n0 175.661
R3943 a_17359_n2247.n0 a_17359_n2247.t3 166.739
R3944 a_24530_n22338.t0 a_24530_n22338.t1 81.9492
R3945 dout_filt.n0 dout_filt.t2 687.288
R3946 x7.clkout dout_filt.t0 229.845
R3947 dout_filt.n1 dout_filt.t1 223.571
R3948 dout_filt.n1 dout_filt.n0 139.672
R3949 dout_filt.n2 dout_filt.t4 97.4114
R3950 dout_filt.n2 dout_filt.t3 56.9639
R3951 x7.clkout x7.x5.Z 28.6323
R3952 x7.x5.Z x7.clkout 28.3622
R3953 x7.clkout dout_filt.n2 10.5187
R3954 x7.x5.Z dout_filt.n1 4.70638
R3955 x7.x5.Z dout_filt.n0 4.70638
R3956 x4.out_b.n0 x4.out_b.t0 227.887
R3957 x4.out_b.n0 x4.out_b.n1 25.0905
R3958 x4.out_b.n0 x4.out_b.t3 12.777
R3959 x4.out_b.n1 x4.out_b.t1 5.5105
R3960 x4.out_b.n1 x4.out_b.t2 5.5105
R3961 x4.out_b x4.out_b.n0 0.83175
R3962 a_15960_n1881.n1 a_15960_n1881.n0 926.024
R3963 a_15960_n1881.n1 a_15960_n1881.t3 82.0838
R3964 a_15960_n1881.n0 a_15960_n1881.t2 63.3338
R3965 a_15960_n1881.t0 a_15960_n1881.n1 63.3219
R3966 a_15960_n1881.n0 a_15960_n1881.t1 29.7268
R3967 a_20471_n2791.n3 a_20471_n2791.n2 674.338
R3968 a_20471_n2791.n1 a_20471_n2791.t5 332.58
R3969 a_20471_n2791.n2 a_20471_n2791.n0 284.012
R3970 a_20471_n2791.n2 a_20471_n2791.n1 253.648
R3971 a_20471_n2791.n1 a_20471_n2791.t4 168.701
R3972 a_20471_n2791.t1 a_20471_n2791.n3 96.1553
R3973 a_20471_n2791.n3 a_20471_n2791.t3 65.6672
R3974 a_20471_n2791.n0 a_20471_n2791.t0 65.0005
R3975 a_20471_n2791.n0 a_20471_n2791.t2 45.0005
R3976 a_24220_n9168.t0 a_24220_n9168.t1 83.56
R3977 a_21036_n2791.n3 a_21036_n2791.n2 636.953
R3978 a_21036_n2791.n1 a_21036_n2791.t5 366.856
R3979 a_21036_n2791.n2 a_21036_n2791.n0 300.2
R3980 a_21036_n2791.n2 a_21036_n2791.n1 225.036
R3981 a_21036_n2791.n1 a_21036_n2791.t4 174.056
R3982 a_21036_n2791.n0 a_21036_n2791.t2 70.0005
R3983 a_21036_n2791.t1 a_21036_n2791.n3 68.0124
R3984 a_21036_n2791.n3 a_21036_n2791.t3 63.3219
R3985 a_21036_n2791.n0 a_21036_n2791.t0 61.6672
R3986 a_18937_n1869.n0 a_18937_n1869.t0 68.3338
R3987 a_18937_n1869.n0 a_18937_n1869.t1 26.3935
R3988 a_18937_n1869.n1 a_18937_n1869.n0 14.4005
R3989 a_17747_n2791.n1 a_17747_n2791.t7 530.01
R3990 a_17747_n2791.t0 a_17747_n2791.n5 421.021
R3991 a_17747_n2791.n0 a_17747_n2791.t6 337.142
R3992 a_17747_n2791.n3 a_17747_n2791.t1 280.223
R3993 a_17747_n2791.n4 a_17747_n2791.t3 263.173
R3994 a_17747_n2791.n4 a_17747_n2791.t5 227.826
R3995 a_17747_n2791.n0 a_17747_n2791.t2 199.762
R3996 a_17747_n2791.n2 a_17747_n2791.n1 170.81
R3997 a_17747_n2791.n2 a_17747_n2791.n0 167.321
R3998 a_17747_n2791.n5 a_17747_n2791.n4 152
R3999 a_17747_n2791.n1 a_17747_n2791.t4 141.923
R4000 a_17747_n2791.n3 a_17747_n2791.n2 10.8376
R4001 a_17747_n2791.n5 a_17747_n2791.n3 2.50485
R4002 a_17359_n2791.t0 a_17359_n2791.n1 386.31
R4003 a_17359_n2791.n1 a_17359_n2791.t1 249.956
R4004 a_17359_n2791.n0 a_17359_n2791.t3 239.04
R4005 a_17359_n2791.n1 a_17359_n2791.n0 175.661
R4006 a_17359_n2791.n0 a_17359_n2791.t2 166.739
R4007 a_2130_n20512.t0 a_2130_n20512.t1 82.0028
R4008 a_18263_n2791.n3 a_18263_n2791.n2 674.338
R4009 a_18263_n2791.n1 a_18263_n2791.t4 332.58
R4010 a_18263_n2791.n2 a_18263_n2791.n0 284.012
R4011 a_18263_n2791.n2 a_18263_n2791.n1 253.648
R4012 a_18263_n2791.n1 a_18263_n2791.t5 168.701
R4013 a_18263_n2791.t1 a_18263_n2791.n3 96.1553
R4014 a_18263_n2791.n3 a_18263_n2791.t3 65.6672
R4015 a_18263_n2791.n0 a_18263_n2791.t0 65.0005
R4016 a_18263_n2791.n0 a_18263_n2791.t2 45.0005
R4017 a_2132_n14926.t0 a_2132_n14926.t1 83.9223
R4018 a_18932_n15092.t0 a_18932_n15092.t1 83.5579
R4019 a_14357_n2743.t0 a_14357_n2743.t1 64.6411
R4020 dout.n0 dout.t1 120.561
R4021 dout.n0 dout.t0 61.4115
R4022 dout dout.n0 3.88384
R4023 a_20376_n1881.n1 a_20376_n1881.n0 926.024
R4024 a_20376_n1881.n1 a_20376_n1881.t2 82.0838
R4025 a_20376_n1881.n0 a_20376_n1881.t3 63.3338
R4026 a_20376_n1881.t0 a_20376_n1881.n1 63.3219
R4027 a_20376_n1881.n0 a_20376_n1881.t1 29.7268
R4028 a_20471_n1869.n3 a_20471_n1869.n2 674.338
R4029 a_20471_n1869.n1 a_20471_n1869.t5 332.58
R4030 a_20471_n1869.n2 a_20471_n1869.n0 284.012
R4031 a_20471_n1869.n2 a_20471_n1869.n1 253.648
R4032 a_20471_n1869.n1 a_20471_n1869.t4 168.701
R4033 a_20471_n1869.n3 a_20471_n1869.t3 96.1553
R4034 a_20471_n1869.t1 a_20471_n1869.n3 65.6672
R4035 a_20471_n1869.n0 a_20471_n1869.t2 65.0005
R4036 a_20471_n1869.n0 a_20471_n1869.t0 45.0005
R4037 x7.x1.Qb1.n4 x7.x1.Qb1.t0 372.361
R4038 x7.x1.Qb1.n2 x7.x1.Qb1.t4 333.651
R4039 x7.x1.Qb1.n2 x7.x1.Qb1.t5 297.233
R4040 x7.x1.Qb1.n0 x7.x1.Qb1.t2 294.557
R4041 x7.x1.Qb1.n5 x7.x1.Qb1.t1 231.921
R4042 x7.x1.Qb1.n0 x7.x1.Qb1.t3 211.01
R4043 x7.x1.Qb1 x7.x1.Qb1.n2 195.701
R4044 x7.x1.Qb1.n1 x7.x1.Qb1.n0 152
R4045 x7.x1.Qb1.n5 x7.x1.Qb1.n1 41.5091
R4046 x7.x1.Qb1.n5 x7.x1.Qb1.n4 18.1966
R4047 x7.x1.Qb1.n4 x7.x1.Qb1.n3 9.35675
R4048 x7.x1.Qb1.n3 x7.x1.Qb1 6.49269
R4049 x7.x1.Qb1.n1 x7.x1.Qb1 4.20621
R4050 x7.x1.Qb1.n3 x7.x1.Qb1 3.52967
R4051 x7.x1.Qb1 x7.x1.Qb1.n5 2.5605
R4052 x7.x2.x2.Q x7.x2.x2.Q.t0 246.839
R4053 x7.x2.x2.Q x7.x2.x2.Q.t1 148.597
R4054 a_14035_n2743.t0 a_14035_n2743.t1 60.0005
R4055 a_24530_n20346.t0 a_24530_n20346.t1 81.9478
R4056 a_18932_n14760.t0 a_18932_n14760.t1 83.5579
R4057 x7.x1.x3.Q x7.x1.x3.Q.t0 240.05
R4058 x7.x1.x3.Q x7.x1.x3.Q.t1 155.386
R4059 a_2130_n19184.t0 a_2130_n19184.t1 82.0028
R4060 a_24530_n19018.t0 a_24530_n19018.t1 81.9478
R4061 a_10620_n9002.t0 a_10620_n9002.t1 83.9243
R4062 a_14035_n2281.t0 a_14035_n2281.t1 60.9236
R4063 a_24220_n8836.t0 a_24220_n8836.t1 83.56
R4064 a_2130_n20180.t0 a_2130_n20180.t1 82.0028
R4065 a_2130_n22172.t0 a_2130_n22172.t1 82.0028
R4066 a_24530_n22006.t0 a_24530_n22006.t1 81.9492
R4067 a_2130_n21840.t0 a_2130_n21840.t1 82.0028
R4068 a_2132_n16586.t0 a_2132_n16586.t1 83.9223
R4069 a_18932_n16420.t0 a_18932_n16420.t1 83.5579
R4070 a_10620_n8670.t0 a_10620_n8670.t1 83.9243
R4071 a_22601_n15524.t0 a_22601_n15524.t1 120.212
R4072 a_20579_n2425.n0 a_20579_n2425.t1 1327.82
R4073 a_20579_n2425.t0 a_20579_n2425.n0 194.655
R4074 a_20579_n2425.n0 a_20579_n2425.t2 63.3219
R4075 a_21198_n2247.t0 a_21198_n2247.t1 126.644
R4076 a_17747_n2241.n1 a_17747_n2241.t4 530.01
R4077 a_17747_n2241.t0 a_17747_n2241.n5 421.021
R4078 a_17747_n2241.n0 a_17747_n2241.t2 337.142
R4079 a_17747_n2241.n3 a_17747_n2241.t1 280.223
R4080 a_17747_n2241.n4 a_17747_n2241.t3 263.173
R4081 a_17747_n2241.n4 a_17747_n2241.t6 227.826
R4082 a_17747_n2241.n0 a_17747_n2241.t5 199.762
R4083 a_17747_n2241.n2 a_17747_n2241.n1 170.81
R4084 a_17747_n2241.n2 a_17747_n2241.n0 167.321
R4085 a_17747_n2241.n5 a_17747_n2241.n4 152
R4086 a_17747_n2241.n1 a_17747_n2241.t7 141.923
R4087 a_17747_n2241.n3 a_17747_n2241.n2 10.8376
R4088 a_17747_n2241.n5 a_17747_n2241.n3 2.50485
R4089 a_2132_n14594.t0 a_2132_n14594.t1 82.3314
R4090 a_18932_n14428.t0 a_18932_n14428.t1 83.5579
R4091 a_16163_n2425.n0 a_16163_n2425.t2 1327.82
R4092 a_16163_n2425.n0 a_16163_n2425.t1 194.655
R4093 a_16163_n2425.t0 a_16163_n2425.n0 63.3219
R4094 a_18371_n2247.n0 a_18371_n2247.t2 1327.82
R4095 a_18371_n2247.t0 a_18371_n2247.n0 194.655
R4096 a_18371_n2247.n0 a_18371_n2247.t1 63.3219
R4097 a_24220_n8504.t0 a_24220_n8504.t1 83.56
R4098 x7.x2.x4.Q x7.x2.x4.Q.t0 246.839
R4099 x7.x2.x4.Q x7.x2.x4.Q.t1 148.597
R4100 a_18932_n16752.t0 a_18932_n16752.t1 83.5579
R4101 a_2130_n21508.t0 a_2130_n21508.t1 82.0028
R4102 a_24530_n21674.t0 a_24530_n21674.t1 81.9478
R4103 a_21390_n2791.t0 a_21390_n2791.t1 87.1434
R4104 a_2130_n18852.t0 a_2130_n18852.t1 82.0028
R4105 a_21390_n1881.t0 a_21390_n1881.t1 87.1434
R4106 a_8268_n12482.t1 a_8268_n12482.t0 193.599
R4107 a_21145_n2791.t1 a_21145_n2791.t0 94.7268
R4108 a_16782_n2247.t0 a_16782_n2247.t1 126.644
R4109 x7.x2.x3.Q x7.x2.x3.Q.t0 246.839
R4110 x7.x2.x3.Q x7.x2.x3.Q.t1 148.597
R4111 a_10620_n8006.t0 a_10620_n8006.t1 83.9243
R4112 a_2132_n16254.t0 a_2132_n16254.t1 83.9053
R4113 a_16729_n2791.t0 a_16729_n2791.t1 94.7268
R4114 a_2132_n17914.t0 a_2132_n17914.t1 83.9223
R4115 a_21198_n2425.t0 a_21198_n2425.t1 126.644
R4116 a_18932_n16088.t0 a_18932_n16088.t1 83.5579
R4117 a_18371_n2425.n0 a_18371_n2425.t1 1327.82
R4118 a_18371_n2425.t0 a_18371_n2425.n0 194.655
R4119 a_18371_n2425.n0 a_18371_n2425.t2 63.3219
R4120 a_18990_n2247.t0 a_18990_n2247.t1 126.644
R4121 a_2132_n14262.t0 a_2132_n14262.t1 83.9053
R4122 a_2132_n15922.t0 a_2132_n15922.t1 83.9223
C0 x7.x2.x3.Q x7.x2.Qb2 0.040893f
C1 vg1 xin 0.215332p
C2 x7.ena_done_b x7.x1.Qb1 0.095485f
C3 x7.x1.x3.Q x7.x1.Qb2 0.040893f
C4 vg2 xout 0.938912f
C5 dvss_ip tail 0.416372f
C6 avss_ip xout 26.396301f
C7 avss_ip x3.out 2.42666f
C8 dvdd_ip avdd_ip 3.92913f
C9 ibias_ip dvss_ip 20.3173f
C10 avss avdd 0.11051p
C11 x7.ena_done_b x7.stby_done_b 1.61077f
C12 dvdd_ip inv_in 10.408401f
C13 inv_in vbp 0.265485f
C14 vg1 xout 0.637062f
C15 x7.x1.x2.CLK dvdd 0.406962f
C16 dvdd standby 0.386478f
C17 dvdd standby_33 0.092517f
C18 dvdd x7.x1.Qb2 1.22125f
C19 x7.x2.x4.Q x7.stby_done_b 0.061065f
C20 dvdd_ip dvss_ip 0.502488p
C21 x7.x2.x2.Q x7.stby_done_b 0.012057f
C22 x7.x1.x3.Q x7.ena_done_b 0.012117f
C23 ibias dvdd 0.083154f
C24 dvss_ip vbp 1.28877f
C25 dvdd_ip inv_m1 2.8465f
C26 ibias_ip standby_33 0.622578f
C27 inv_in vn 0.137437f
C28 x3.out avdd 9.26841f
C29 standby_33 x4.out_b 0.696369f
C30 dvdd_ip vrb 0.182588f
C31 x7.x1.x2.CLK x7.x2.x2.CLK 0.011009f
C32 dvdd_ip vg2 0.10449f
C33 x7.ena_done_b x7.x1.x2.Q 0.012057f
C34 ibias_ip ibias 0.846688f
C35 dvdd_ip avss_ip 2.34725f
C36 avdd dvdd 0.151932f
C37 x7.x1.x2.Q x7.x1.Qb1 0.040893f
C38 ena standby 0.095384f
C39 standby_ip standby 0.045124f
C40 dvss_ip ena_ip 0.012218f
C41 dvss_ip vn 6.6789f
C42 dvdd_ip inv_m2 1.90217f
C43 dvdd_ip standby_33 3.32f
C44 x7.ena_done_b dvdd 6.16668f
C45 x7.clk_disable x7.stby_done_b 0.724301f
C46 avdd_ip inv_in 0.669037f
C47 x7.x1.Qb1 dvdd 1.22948f
C48 ibias standby_ip 0.288754f
C49 dvdd_ip vg1 0.707385f
C50 dvdd dout 0.550876f
C51 dvdd_ip ibias 0.012207f
C52 avdd x4.out_b 7.47205f
C53 x3.out avss 5.85073f
C54 x7.ena_done_b x7.x1.x4.Q 0.061065f
C55 x7.x2.x4.Q dvdd 0.118417f
C56 dvdd x7.stby_done_b 5.41509f
C57 dvdd x7.x2.x2.Q 0.11753f
C58 avdd_ip dvss_ip 20.9126f
C59 xin xout 12.4168f
C60 ena avdd 0.026836f
C61 avss dvdd 0.230608f
C62 avdd standby_ip 0.691145f
C63 x7.x1.x2.CLK ena_ip 0.073063f
C64 dvss_ip inv_in 14.9295f
C65 ena_ip standby 0.035742f
C66 x7.x2.x3.Q x7.stby_done_b 0.012117f
C67 dvdd_ip avdd 0.116559f
C68 ena_ip x7.x1.Qb2 0.347451f
C69 inv_in inv_m1 0.243271f
C70 x7.ena_done_b standby_ip 0.121215f
C71 x7.x2.Qb1 x7.x1.Qb1 0.0262f
C72 dvss_ip x7.x2.Qb2 0.073361f
C73 ibias ena_ip 0.172379f
C74 x7.x1.x3.Q dvdd 0.112744f
C75 dvdd_ip x7.ena_done_b 0.022633f
C76 avdd_ip vg2 0.280688f
C77 avdd_ip avss_ip 0.843902p
C78 xin tail 1.6128f
C79 avss x4.out_b 1.60462f
C80 x7.x2.x2.CLK x7.stby_done_b 0.055466f
C81 inv_in vg2 0.137694f
C82 dvdd_ip dout 1.66314f
C83 dvss_ip inv_m1 3.10116f
C84 x7.x2.Qb1 x7.stby_done_b 0.111333f
C85 avss_ip inv_in 1.9489f
C86 x7.x2.Qb1 x7.x2.x2.Q 0.040893f
C87 dvdd x7.clk_disable 0.383458f
C88 dvdd_ip x7.stby_done_b 0.02481f
C89 x7.x1.x2.Q dvdd 0.116301f
C90 ena_ip avdd 0.712717f
C91 avss standby_ip 1.86774f
C92 dvss_ip vrb 1.20334f
C93 inv_in standby_33 0.08455f
C94 avdd_ip vg1 1.83467f
C95 dvdd_ip avss 0.031818f
C96 dvss_ip vg2 3.9276f
C97 dvss_ip avss_ip 24.1368f
C98 x7.ena_done_b ena_ip 0.702741f
C99 xout tail 1.23159f
C100 x7.x1.Qb1 ena_ip 0.347396f
C101 dvss_ip inv_m2 1.69984f
C102 dvdd_ip xin 4.32555f
C103 dvss_ip standby_33 3.43231f
C104 x7.x2.Qb2 x7.x1.Qb2 0.0262f
C105 x7.x2.x3.Q dvdd 0.112734f
C106 inv_m1 inv_m2 0.947856f
C107 vrb vg2 4.64006f
C108 dvss_ip x7.x1.Qb2 0.069883f
C109 x7.clk_disable x7.x2.x2.CLK 0.012819f
C110 avss_ip vrb 6.48162f
C111 avdd_ip avdd 9.334331f
C112 dvdd x7.x1.x4.Q 0.118427f
C113 dvss_ip vg1 6.37401f
C114 ibias_ip dvdd 0.020082f
C115 dvss_ip ibias 0.014158f
C116 avss_ip vg2 0.156018p
C117 inv_in avdd 0.025173f
C118 avss ena_ip 1.87864f
C119 dvdd_ip xout 4.80514f
C120 dvdd x7.x2.x2.CLK 0.367738f
C121 ibias_ip tail 0.011037f
C122 x7.x2.Qb1 dvdd 1.15446f
C123 vg1 vrb 0.454276f
C124 ena dvdd 0.377442f
C125 vn xin 3.09633f
C126 dvdd standby_ip 10.361099f
C127 x7.x1.x3.Q ena_ip 0.035311f
C128 vg1 vg2 1.36272f
C129 dvdd_ip dvdd 14.0421f
C130 avss_ip vg1 20.7774f
C131 dvss_ip x7.ena_done_b 1.48709f
C132 avdd_ip avss 0.574893f
C133 dvdd_ip tail 3.21426f
C134 ibias standby_33 1.11388f
C135 inv_in avss 0.144174f
C136 x7.x1.x2.Q ena_ip 0.035311f
C137 x4.out_b standby_ip 0.931668f
C138 vbp tail 10.143401f
C139 avdd_ip xin 6.15469f
C140 dvss_ip dout 6.66227f
C141 vn xout 0.039662f
C142 ibias_ip dvdd_ip 1.4709f
C143 x7.x2.Qb2 x7.stby_done_b 0.099468f
C144 avss_ip avdd 2.34938f
C145 ibias_ip vbp 1.36181f
C146 inv_in xin 0.302115f
C147 dvss_ip x7.stby_done_b 1.50207f
C148 ena_ip dvdd 7.78514f
C149 avdd standby_33 9.00234f
C150 dvdd_ip standby_ip 3.51143f
C151 x7.ena_done_b x7.x1.x2.CLK 0.044383f
C152 vn tail 0.670061f
C153 avdd_ip xout 7.21813f
C154 dvss_ip xin 1.63056f
C155 avdd_ip x3.out 0.010186f
C156 dvdd_ip vbp 26.197498f
C157 x7.ena_done_b x7.x1.Qb2 0.095442f
C158 inv_in xout 1.1656f
C159 avss_ip avss 7.313931f
C160 inv_in dvdd 0.696511f
C161 ena ena_ip 0.081602f
C162 ena_ip standby_ip 4.64341f
C163 vg2 xin 6.28706f
C164 avss_ip xin 73.1079f
C165 dvss_ip xout 14.2041f
C166 avss standby_33 1.55853f
C167 dvdd_ip vn 1.05192f
C168 inv_in tail 0.604094f
C169 dvdd x7.x2.Qb2 1.2179f
C170 dvss_ip dvdd 20.2592f
C171 ibias_ip inv_in 0.023743f
C172 xout dvss 4.205515f
C173 xin dvss 11.862524f
C174 dout dvss 4.99223f
C175 standby dvss 1.31811f
C176 ena dvss 1.29717f
C177 avss dvss 9.38759f
C178 ibias dvss 5.68171f
C179 dvdd dvss 0.138268p
C180 avdd dvss 93.42453f
C181 vg1 dvss -0.243245f
C182 vrb dvss 0.16284f
C183 vg2 dvss 4.395665f
C184 tail dvss 12.477897f
C185 inv_m2 dvss 0.561945f
C186 inv_m1 dvss 1.14191f
C187 inv_in dvss 6.33693f
C188 vn dvss 7.76391f
C189 vbp dvss 19.58865f
C190 x4.out_b dvss 1.060934f
C191 x3.out dvss 2.07711f
C192 x7.x2.x4.Q dvss 0.099773f
C193 x7.x2.x3.Q dvss 0.092032f
C194 x7.x2.Qb2 dvss 0.510343f
C195 x7.x2.x2.Q dvss 0.092454f
C196 x7.x2.Qb1 dvss 0.539804f
C197 x7.x2.x2.CLK dvss 0.389657f
C198 x7.clk_disable dvss 4.59421f
C199 x7.x1.x4.Q dvss 0.099773f
C200 x7.x1.x3.Q dvss 0.092032f
C201 x7.x1.x2.Q dvss 0.092454f
C202 x7.stby_done_b dvss 3.879532f
C203 ibias_ip dvss 12.69437f
C204 standby_33 dvss 11.1604f
C205 x7.x1.Qb2 dvss 0.511115f
C206 x7.x1.Qb1 dvss 0.528314f
C207 x7.x1.x2.CLK dvss 0.382316f
C208 x7.ena_done_b dvss 5.915554f
C209 standby_ip dvss 22.070288f
C210 ena_ip dvss 24.167025f
C211 avss_ip dvss 11.3398f
C212 dvss_ip dvss 36.609398f
C213 avdd_ip dvss 0.929763p
C214 dvdd_ip dvss 0.361469p
C215 a_8268_n12482.t1 dvss 0.033931f
C216 a_8268_n12482.t0 dvss 3.56607f
C217 a_22601_n15524.t1 dvss 1.2f
C218 a_22601_n15524.t0 dvss 1.2f
C219 dout.t1 dvss 0.040138f
C220 dout.t0 dvss 0.223213f
C221 dout.n0 dvss 3.29562f
C222 x4.out_b.n0 dvss 5.53652f
C223 x4.out_b.t3 dvss 1.30743f
C224 x4.out_b.t1 dvss 0.044437f
C225 x4.out_b.t2 dvss 0.044437f
C226 x4.out_b.n1 dvss 0.140668f
C227 x4.out_b.t0 dvss 0.055178f
C228 x7.clkout dvss 5.76435f
C229 dout_filt.t2 dvss 0.033084f
C230 dout_filt.n0 dvss 0.063466f
C231 dout_filt.t1 dvss 0.020119f
C232 dout_filt.n1 dvss 0.064349f
C233 x7.x5.Z dvss 0.084653f
C234 dout_filt.t0 dvss 0.028544f
C235 dout_filt.t3 dvss 0.296603f
C236 dout_filt.t4 dvss 0.738515f
C237 dout_filt.n2 dvss 6.50632f
C238 x3.out.n0 dvss 7.39524f
C239 x3.out.n1 dvss 0.893601f
C240 x3.out.n2 dvss 0.392503f
C241 x3.out.t6 dvss 0.479128f
C242 x3.out.n3 dvss 0.382459f
C243 x3.out.t8 dvss 0.458669f
C244 x3.out.n4 dvss 0.394877f
C245 x3.out.t7 dvss 0.479113f
C246 x3.out.t4 dvss 0.458669f
C247 x3.out.n5 dvss 0.382543f
C248 x3.out.t3 dvss 0.458669f
C249 x3.out.n6 dvss 0.161457f
C250 x3.out.n7 dvss 0.521199f
C251 x3.out.n8 dvss 1.69978f
C252 x3.out.t5 dvss 1.7568f
C253 x3.out.t1 dvss 0.059712f
C254 x3.out.t2 dvss 0.059712f
C255 x3.out.n9 dvss 0.188953f
C256 x3.out.t0 dvss 0.074144f
C257 vn.n0 dvss 0.636215f
C258 vn.n1 dvss 0.311146f
C259 vn.t7 dvss 0.039422f
C260 vn.t5 dvss 0.039422f
C261 vn.n2 dvss 0.106375f
C262 vn.t6 dvss 0.171883f
C263 vn.n3 dvss 0.444704f
C264 vn.t8 dvss 0.871134f
C265 vn.t9 dvss 1.02426f
C266 vn.n4 dvss 0.591267f
C267 vn.n5 dvss 0.320978f
C268 vn.t0 dvss 0.973785f
C269 vn.t4 dvss 0.039422f
C270 vn.t1 dvss 0.039422f
C271 vn.n6 dvss 0.078843f
C272 vn.t2 dvss 0.133384f
C273 vn.n7 dvss 0.489753f
C274 vn.n8 dvss 0.299827f
C275 vn.t3 dvss 0.871134f
C276 vn.n9 dvss 0.296493f
C277 vrb.t1 dvss 0.274519f
C278 vrb.t3 dvss 0.33602f
C279 vrb.n0 dvss 3.02505f
C280 vrb.t2 dvss 0.274548f
C281 vrb.t0 dvss 0.333171f
C282 vrb.n1 dvss 3.02989f
C283 vrb.t4 dvss 0.080693f
C284 vrb.n2 dvss 2.40037f
C285 vrb.n3 dvss 1.30448f
C286 vg2.n0 dvss 0.282949f
C287 vg2.n1 dvss 0.261019f
C288 vg2.t9 dvss 0.640509f
C289 vg2.n2 dvss 1.17147f
C290 vg2.n3 dvss 0.244906f
C291 vg2.n4 dvss 0.522037f
C292 vg2.t6 dvss 0.628646f
C293 vg2.n5 dvss 0.314177f
C294 vg2.n6 dvss 0.32051f
C295 vg2.n7 dvss 0.282949f
C296 vg2.n8 dvss 0.261019f
C297 vg2.t5 dvss 0.640544f
C298 vg2.n9 dvss 1.17258f
C299 vg2.n10 dvss 0.244906f
C300 vg2.n11 dvss 0.522037f
C301 vg2.t7 dvss 0.628646f
C302 vg2.n12 dvss 0.313029f
C303 vg2.n13 dvss 0.32051f
C304 vg2.n14 dvss 0.051368f
C305 vg2.t0 dvss 0.031316f
C306 vg2.t8 dvss 0.505469f
C307 vg2.t2 dvss 39.125f
C308 vg2.t1 dvss 39.3426f
C309 vg2.t4 dvss 39.3426f
C310 vg2.t3 dvss 39.11f
C311 vg2.n15 dvss 9.00528f
C312 vg2.n16 dvss 2.91513f
C313 xin.t21 dvss 0.023931f
C314 xin.t8 dvss 0.023302f
C315 xin.n0 dvss 0.172553f
C316 xin.n1 dvss 0.096625f
C317 xin.n2 dvss 0.096625f
C318 xin.n3 dvss 0.096625f
C319 xin.n4 dvss 0.096625f
C320 xin.n5 dvss 0.183862f
C321 xin.t18 dvss 0.191901f
C322 xin.t15 dvss 0.191811f
C323 xin.n6 dvss 0.183862f
C324 xin.n7 dvss 0.096625f
C325 xin.t13 dvss 0.191811f
C326 xin.n8 dvss 0.096625f
C327 xin.t19 dvss 0.191811f
C328 xin.n9 dvss 0.096625f
C329 xin.n10 dvss 0.096625f
C330 xin.t16 dvss 0.191811f
C331 xin.n11 dvss 0.096625f
C332 xin.t11 dvss 0.191811f
C333 xin.n12 dvss 0.096625f
C334 xin.n13 dvss 0.096625f
C335 xin.t10 dvss 0.191811f
C336 xin.n14 dvss 0.096625f
C337 xin.t17 dvss 0.191811f
C338 xin.n15 dvss 0.096625f
C339 xin.n16 dvss 0.096625f
C340 xin.t14 dvss 0.191811f
C341 xin.n17 dvss 0.096625f
C342 xin.t12 dvss 0.191811f
C343 xin.n18 dvss 0.096625f
C344 xin.n19 dvss 0.096625f
C345 xin.t9 dvss 0.191811f
C346 xin.n20 dvss 0.096625f
C347 xin.t6 dvss 0.191811f
C348 xin.n21 dvss 0.17495f
C349 xin.n22 dvss 0.783747f
C350 xin.n23 dvss 0.308143f
C351 xin.n24 dvss 0.374177f
C352 xin.t20 dvss 0.826777f
C353 xin.t7 dvss 0.795041f
C354 xin.n25 dvss 0.5132f
C355 xin.n26 dvss 0.386346f
C356 xin.n27 dvss 3.78897f
C357 xin.n28 dvss 4.51207f
C358 xin.n29 dvss 3.60717f
C359 xin.t1 dvss 56.9351f
C360 xin.t3 dvss 44.1175f
C361 xin.t0 dvss 43.9435f
C362 xin.t5 dvss 0.124032f
C363 xin.n30 dvss 4.76717f
C364 xin.n31 dvss 27.2312f
C365 xin.t4 dvss 31.1439f
C366 xin.n32 dvss 27.2243f
C367 xin.t2 dvss 31.1129f
C368 xin.n33 dvss 27.2277f
C369 xin.n34 dvss 3.77116f
C370 xin.n35 dvss 1.85382f
C371 xin.n36 dvss 0.499796f
C372 vg1.t3 dvss 0.056949f
C373 vg1.n0 dvss 0.44953f
C374 vg1.t8 dvss 46.057503f
C375 vg1.t9 dvss 46.8352f
C376 vg1.t4 dvss 23.996801f
C377 vg1.n1 dvss 23.9575f
C378 vg1.t7 dvss 23.996801f
C379 vg1.n2 dvss 23.4861f
C380 vg1.t6 dvss 23.996801f
C381 vg1.n3 dvss 12.9859f
C382 vg1.n4 dvss 15.228601f
C383 vg1.t2 dvss 0.01371f
C384 vg1.n5 dvss 3.04049f
C385 vg1.n6 dvss 1.50262f
C386 vg1.t0 dvss 0.271659f
C387 vg1.t5 dvss 0.353472f
C388 vg1.n7 dvss 0.229145f
C389 vg1.n8 dvss 0.08087f
C390 vg1.t1 dvss 0.049005f
C391 vg1.n9 dvss 0.281876f
C392 vg1.n10 dvss 0.146945f
C393 vg1.n11 dvss 0.153437f
C394 vg1.n12 dvss 0.372304f
C395 x3.out_b.t6 dvss 0.402581f
C396 x3.out_b.n0 dvss 0.790285f
C397 x3.out_b.n1 dvss 1.5584f
C398 x3.out_b.n2 dvss 6.60541f
C399 x3.out_b.t4 dvss 0.420289f
C400 x3.out_b.n3 dvss 0.339622f
C401 x3.out_b.t7 dvss 0.402581f
C402 x3.out_b.n4 dvss 0.342378f
C403 x3.out_b.t8 dvss 0.420331f
C404 x3.out_b.n5 dvss 0.338349f
C405 x3.out_b.t3 dvss 0.402581f
C406 x3.out_b.n6 dvss 0.345348f
C407 x3.out_b.n7 dvss 0.58218f
C408 x3.out_b.t5 dvss 1.5189f
C409 x3.out_b.t1 dvss 0.051624f
C410 x3.out_b.t2 dvss 0.051624f
C411 x3.out_b.n8 dvss 0.163419f
C412 x3.out_b.t0 dvss 0.064102f
C413 avdd.n0 dvss 0.492818f
C414 avdd.t19 dvss 0.034087f
C415 avdd.n1 dvss 1.6981f
C416 avdd.n2 dvss 0.060856f
C417 avdd.n3 dvss 0.056499f
C418 avdd.n4 dvss 0.266474f
C419 avdd.n5 dvss 0.585389f
C420 avdd.n6 dvss 1.03476f
C421 avdd.n7 dvss 1.03476f
C422 avdd.t17 dvss 0.894926f
C423 avdd.t3 dvss 0.702496f
C424 avdd.t5 dvss 0.894926f
C425 avdd.t9 dvss 0.702496f
C426 avdd.n8 dvss 0.46232f
C427 avdd.t14 dvss 7.53658f
C428 avdd.n9 dvss 7.5153f
C429 avdd.t13 dvss 9.12027f
C430 avdd.t16 dvss 7.25381f
C431 avdd.n10 dvss 7.71793f
C432 avdd.t15 dvss 9.163919f
C433 avdd.n11 dvss 3.68652f
C434 avdd.n12 dvss 0.768588f
C435 avdd.n13 dvss 0.579746f
C436 avdd.n14 dvss 0.560241f
C437 avdd.n15 dvss 0.353066f
C438 avdd.n16 dvss 0.487874f
C439 avdd.n17 dvss 3.7478f
C440 avdd.n18 dvss 0.731215f
C441 avdd.t10 dvss 0.036998f
C442 avdd.t6 dvss 0.036998f
C443 avdd.n19 dvss 0.090684f
C444 avdd.t4 dvss 0.036998f
C445 avdd.t12 dvss 0.036998f
C446 avdd.n20 dvss 0.090684f
C447 avdd.n21 dvss 1.93441f
C448 avdd.n22 dvss 0.967373f
C449 avdd.t18 dvss 0.135207f
C450 avdd.n23 dvss 0.34342f
C451 avdd.n24 dvss 5.68989f
C452 avdd.n25 dvss 1.05169f
C453 avdd.n26 dvss 1.1887f
C454 avdd.n27 dvss 1.1887f
C455 avdd.n28 dvss 4.46094f
C456 avdd.n29 dvss 1.35368f
C457 avdd.n30 dvss 0.090671f
C458 avdd.n31 dvss 0.071983f
C459 avdd.n32 dvss 0.548551f
C460 avdd.n33 dvss 1.56238f
C461 avdd.t2 dvss 0.034087f
C462 avdd.n34 dvss 1.46595f
C463 avdd.n35 dvss 0.107384f
C464 avdd.n36 dvss 0.107943f
C465 avdd.n37 dvss 0.158157f
C466 avdd.t0 dvss 2.51038f
C467 avdd.n38 dvss 0.071983f
C468 avdd.n39 dvss 0.10415f
C469 avdd.n40 dvss 0.107943f
C470 avdd.n41 dvss 0.559667f
C471 avdd.t1 dvss 0.034087f
C472 avdd.n42 dvss 0.023315f
C473 avdd.n43 dvss 0.687088f
C474 avdd.n44 dvss 1.48367f
C475 avdd.n45 dvss 1.13727f
C476 avdd.n46 dvss 0.744579f
C477 avdd.n47 dvss 2.46523f
C478 avdd.n48 dvss 3.43088f
C479 avdd.n49 dvss 1.15288f
C480 avdd.n50 dvss 0.362301f
C481 avdd.n51 dvss 0.321745f
C482 avdd.n52 dvss 0.106191f
C483 avdd.n53 dvss 1.67879f
C484 avdd.n54 dvss 0.106191f
C485 avdd.n55 dvss 0.158157f
C486 avdd.n56 dvss 0.090671f
C487 avdd.n57 dvss 0.062903f
C488 avdd.n58 dvss 0.106191f
C489 avdd.n59 dvss 1.67879f
C490 avdd.n60 dvss 0.106191f
C491 avdd.n61 dvss 0.060856f
C492 avdd.n62 dvss 0.116928f
C493 avdd.n63 dvss 0.719248f
C494 avdd.n64 dvss 1.37927f
C495 avdd.n65 dvss 1.47231f
C496 avdd.t8 dvss 0.034087f
C497 avdd.n66 dvss 1.45902f
C498 avdd.n67 dvss 0.366507f
C499 avdd.n68 dvss 0.107943f
C500 avdd.n69 dvss 0.158157f
C501 avdd.t7 dvss 2.51038f
C502 avdd.n70 dvss 0.10415f
C503 avdd.n71 dvss 0.107943f
C504 avdd.n72 dvss 0.107384f
C505 avdd.n73 dvss 0.062903f
C506 avdd.n74 dvss 0.106191f
C507 avdd.n75 dvss 1.67879f
C508 avdd.n76 dvss 0.106191f
C509 avdd.n77 dvss 0.158157f
C510 avdd.n78 dvss 0.106191f
C511 avdd.n79 dvss 1.67879f
C512 avdd.n80 dvss 0.106191f
C513 avdd.n81 dvss 0.319178f
C514 avdd.n82 dvss 0.73302f
C515 avdd.n83 dvss 1.95073f
C516 avdd.n84 dvss 4.13419f
C517 avdd.n85 dvss 0.707422f
C518 avdd.n86 dvss 0.479606f
C519 avdd.n87 dvss 1.32047f
C520 avdd.n88 dvss 1.35617f
C521 avdd.n89 dvss 0.536684f
C522 avdd.n90 dvss 1.19042f
C523 avdd.n91 dvss 4.48227f
C524 avdd.n92 dvss 4.46094f
C525 avdd.n93 dvss 4.48227f
C526 avdd.n94 dvss 1.19042f
C527 avdd.n95 dvss 0.66577f
C528 avdd.n96 dvss 3.27742f
C529 avdd.n97 dvss 0.20944f
C530 avdd.t11 dvss 0.702496f
C531 avdd.n98 dvss 0.20944f
C532 avdd.n99 dvss 0.731637f
C533 avdd.n100 dvss 0.757787f
C534 avdd.n101 dvss 0.146948f
C535 avdd.n102 dvss 0.057614f
C536 avdd.n103 dvss 0.303016f
C537 avss.n0 dvss 0.274689f
C538 avss.n1 dvss 0.256432f
C539 avss.t19 dvss 0.062902f
C540 avss.n2 dvss 0.199691f
C541 avss.n3 dvss 0.027139f
C542 avss.n4 dvss 0.10291f
C543 avss.n5 dvss 0.092262f
C544 avss.n6 dvss 0.092262f
C545 avss.t18 dvss 0.441575f
C546 avss.t16 dvss 0.441575f
C547 avss.n7 dvss 0.044347f
C548 avss.n8 dvss 0.078584f
C549 avss.t17 dvss 0.063155f
C550 avss.t13 dvss 0.063155f
C551 avss.n9 dvss 0.832446f
C552 avss.n10 dvss 0.117588f
C553 avss.t9 dvss 0.062902f
C554 avss.t15 dvss 0.062902f
C555 avss.n11 dvss 0.501337f
C556 avss.n12 dvss 0.044307f
C557 avss.n13 dvss 0.093826f
C558 avss.n14 dvss 0.093826f
C559 avss.n15 dvss 0.506602f
C560 avss.n16 dvss 0.092262f
C561 avss.n17 dvss 0.506602f
C562 avss.t12 dvss 0.441575f
C563 avss.n18 dvss 0.238935f
C564 avss.t14 dvss 0.441575f
C565 avss.n19 dvss 3.28532f
C566 avss.n20 dvss 7.3481f
C567 avss.t8 dvss 0.441575f
C568 avss.n21 dvss 0.093826f
C569 avss.n22 dvss 0.093826f
C570 avss.n23 dvss 0.078584f
C571 avss.n24 dvss 0.152326f
C572 avss.n25 dvss 0.092262f
C573 avss.n26 dvss 0.092262f
C574 avss.n27 dvss 0.238935f
C575 avss.t10 dvss 0.441575f
C576 avss.n28 dvss 0.092262f
C577 avss.n29 dvss 0.506602f
C578 avss.n30 dvss 0.506602f
C579 avss.t20 dvss 0.441575f
C580 avss.t22 dvss 0.441575f
C581 avss.n31 dvss 0.044347f
C582 avss.t11 dvss 0.063155f
C583 avss.t21 dvss 0.063155f
C584 avss.t23 dvss 0.062902f
C585 avss.t1 dvss 0.080794f
C586 avss.n32 dvss 0.370586f
C587 avss.n33 dvss 0.325025f
C588 avss.n34 dvss 0.132878f
C589 avss.n35 dvss 0.404741f
C590 avss.n36 dvss 2.98049f
C591 avss.t4 dvss 0.860518f
C592 avss.t6 dvss 0.732948f
C593 avss.n37 dvss 2.16357f
C594 avss.n38 dvss 1.84584f
C595 avss.t0 dvss 0.841962f
C596 avss.t24 dvss 0.732948f
C597 avss.n39 dvss 0.3741f
C598 avss.n40 dvss 0.133098f
C599 avss.t2 dvss 0.732948f
C600 avss.n41 dvss 0.133098f
C601 avss.n42 dvss 1.68799f
C602 avss.n43 dvss 0.462717f
C603 avss.t3 dvss 0.023705f
C604 avss.t25 dvss 0.023705f
C605 avss.n44 dvss 0.079436f
C606 avss.t5 dvss 0.023705f
C607 avss.t7 dvss 0.023705f
C608 avss.n45 dvss 0.086235f
C609 avss.n46 dvss 1.36147f
C610 avss.n47 dvss 1.03577f
C611 avss.t26 dvss 8.17429f
C612 avss.n48 dvss 7.701231f
C613 avss.t29 dvss 8.17429f
C614 avss.n49 dvss 8.01034f
C615 avss.t28 dvss 8.17429f
C616 avss.n50 dvss 7.90618f
C617 avss.n51 dvss 4.01706f
C618 avss.t27 dvss 8.17429f
C619 avss.n52 dvss 2.18128f
C620 avss.n53 dvss 4.97729f
C621 avss.n54 dvss 1.85282f
C622 avss.n55 dvss 1.94389f
C623 avss.n56 dvss 1.85115f
C624 avss.n57 dvss 0.09532f
C625 avss.n58 dvss 0.227287f
C626 avss.n59 dvss 0.265186f
C627 avss.n60 dvss 0.643717f
C628 avss.n61 dvss 0.274689f
C629 avss.n62 dvss 0.354568f
C630 avss.n63 dvss 0.078584f
C631 avss.n64 dvss 0.102951f
C632 avss.n65 dvss 0.027139f
C633 avss.n66 dvss 0.036993f
C634 avss.n67 dvss 0.093826f
C635 avss.n68 dvss 0.238935f
C636 avss.n69 dvss 0.093826f
C637 avss.n70 dvss 0.036957f
C638 avss.n71 dvss 0.10291f
C639 avss.n72 dvss 0.044307f
C640 avss.n73 dvss 0.117505f
C641 avss.n74 dvss 0.092262f
C642 avss.n75 dvss 0.79544f
C643 avss.n76 dvss 1.9882f
C644 avss.n77 dvss 0.79544f
C645 avss.n78 dvss 0.092262f
C646 avss.n79 dvss 0.117505f
C647 avss.n80 dvss 0.117588f
C648 avss.n81 dvss 0.455799f
C649 avss.n82 dvss 1.20688f
C650 avss.n83 dvss 0.606761f
C651 avss.n84 dvss 0.354568f
C652 avss.n85 dvss 0.078584f
C653 avss.n86 dvss 0.102951f
C654 avss.n87 dvss 0.036993f
C655 avss.n88 dvss 0.093826f
C656 avss.n89 dvss 0.238935f
C657 avss.n90 dvss 0.093826f
C658 avss.n91 dvss 0.036957f
C659 avss.n92 dvss 0.152326f
C660 avss.n93 dvss 0.088692f
C661 avss.n94 dvss 0.162188f
C662 avss.n95 dvss 0.241706f
C663 standby_ip.n0 dvss 0.442006f
C664 standby_ip.n1 dvss 2.94931f
C665 standby_ip.n2 dvss 0.096644f
C666 standby_ip.t1 dvss 0.020548f
C667 standby_ip.t0 dvss 0.029549f
C668 standby_ip.t3 dvss 0.019059f
C669 standby_ip.t14 dvss 0.011911f
C670 standby_ip.n4 dvss 0.034123f
C671 standby_ip.n5 dvss 0.060427f
C672 standby_ip.t10 dvss 0.937707f
C673 standby_ip.n6 dvss 0.647213f
C674 standby_ip.n7 dvss 0.112804f
C675 standby_ip.n8 dvss 0.20956f
C676 standby_ip.t15 dvss 0.303892f
C677 standby_ip.t9 dvss 0.288571f
C678 standby_ip.n9 dvss 0.20956f
C679 standby_ip.n10 dvss 0.112804f
C680 standby_ip.t8 dvss 0.288571f
C681 standby_ip.n11 dvss 0.112804f
C682 standby_ip.t12 dvss 0.288571f
C683 standby_ip.n12 dvss 0.112804f
C684 standby_ip.n13 dvss 0.102826f
C685 standby_ip.t11 dvss 0.288571f
C686 standby_ip.n14 dvss 0.102826f
C687 standby_ip.n15 dvss 0.112804f
C688 standby_ip.n16 dvss 0.21492f
C689 standby_ip.t4 dvss 0.304656f
C690 standby_ip.t6 dvss 0.288571f
C691 standby_ip.n17 dvss 0.213848f
C692 standby_ip.n18 dvss 0.112804f
C693 standby_ip.t17 dvss 0.288571f
C694 standby_ip.n19 dvss 0.112804f
C695 standby_ip.t18 dvss 0.288571f
C696 standby_ip.n20 dvss 0.112804f
C697 standby_ip.n21 dvss 0.099933f
C698 standby_ip.t5 dvss 0.288571f
C699 standby_ip.n22 dvss 0.099933f
C700 standby_ip.t2 dvss 0.264174f
C701 standby_ip.n23 dvss 0.228673f
C702 standby_ip.t13 dvss 0.23888f
C703 standby_ip.t7 dvss 0.238694f
C704 standby_ip.n24 dvss 0.200628f
C705 standby_ip.n25 dvss 0.922727f
C706 standby_ip.t16 dvss 0.273054f
C707 standby_ip.n26 dvss 0.12393f
C708 xin_buf.t0 dvss 0.205358p
C709 xin_buf.t1 dvss 0.22283f
C710 xin_buf.t2 dvss 0.075836f
C711 xin_buf.n0 dvss 0.129036f
C712 xin_buf.t4 dvss 0.263405f
C713 xin_buf.t3 dvss 0.089459f
C714 xin_buf.n1 dvss 0.161326f
C715 x7.x1.x1.A dvss 0.017818f
C716 x7.x1.clkin dvss 0.290534f
C717 x7.x2.x1.A dvss 0.017818f
C718 x7.x2.clkin dvss 0.174689f
C719 x7.x5.A dvss 0.084584f
C720 dout_ip.n0 dvss 3.72627f
C721 x7.clkin dvss 5.05976f
C722 dout_ip.t9 dvss 0.01616f
C723 dout_ip.n1 dvss 0.038785f
C724 dout_ip.t6 dvss 0.012534f
C725 dout_ip.n2 dvss 0.033243f
C726 dout_ip.n3 dvss 0.027616f
C727 dout_ip.n4 dvss 0.027616f
C728 dout_ip.t5 dvss 0.012534f
C729 dout_ip.n5 dvss 0.033243f
C730 dout_ip.n6 dvss 0.35872f
C731 dout_ip.n7 dvss 0.352547f
C732 dout_ip.t3 dvss 0.021945f
C733 dout_ip.t2 dvss 0.021852f
C734 dout_ip.t0 dvss 0.022644f
C735 dout_ip.t1 dvss 0.022607f
C736 inv_m1.t0 dvss 0.046767f
C737 inv_m1.n0 dvss 1.05525f
C738 inv_m1.n1 dvss 0.129812f
C739 inv_m1.t5 dvss 0.363826f
C740 inv_m1.t2 dvss 0.363827f
C741 inv_m1.n2 dvss 0.117923f
C742 inv_m1.t4 dvss 0.341649f
C743 inv_m1.t3 dvss 0.34165f
C744 inv_m1.n3 dvss 2.65565f
C745 inv_m1.t1 dvss 0.045634f
C746 inv_in.t3 dvss 0.657711f
C747 inv_in.t11 dvss 5.68012f
C748 inv_in.n0 dvss 5.17707f
C749 inv_in.t5 dvss 5.52894f
C750 inv_in.n1 dvss 2.62426f
C751 inv_in.t6 dvss 5.52894f
C752 inv_in.n2 dvss 2.66147f
C753 inv_in.n3 dvss 2.79669f
C754 inv_in.t14 dvss 5.52894f
C755 inv_in.n4 dvss 5.29306f
C756 inv_in.t12 dvss 5.55261f
C757 inv_in.n5 dvss 5.28615f
C758 inv_in.t13 dvss 5.52894f
C759 inv_in.n6 dvss 2.66147f
C760 inv_in.t9 dvss 5.5836f
C761 inv_in.n7 dvss 5.39875f
C762 inv_in.t10 dvss 5.5836f
C763 inv_in.t2 dvss 5.5836f
C764 inv_in.n8 dvss 5.26653f
C765 inv_in.n9 dvss 5.40864f
C766 inv_in.t4 dvss 5.52894f
C767 inv_in.n10 dvss 2.66147f
C768 inv_in.n11 dvss 2.90209f
C769 inv_in.n12 dvss 2.75998f
C770 inv_in.t8 dvss 5.52894f
C771 inv_in.n13 dvss 2.62426f
C772 inv_in.n14 dvss 2.76492f
C773 inv_in.n15 dvss 2.76492f
C774 inv_in.n16 dvss 2.76201f
C775 inv_in.t7 dvss 5.52894f
C776 inv_in.n17 dvss 5.4592f
C777 inv_in.n18 dvss 0.82306f
C778 inv_in.t0 dvss 0.104143f
C779 inv_in.t1 dvss 0.647866f
C780 inv_in.n19 dvss 2.16816f
C781 xout.t26 dvss 0.047347f
C782 xout.t24 dvss 0.048657f
C783 xout.t18 dvss 0.243993f
C784 xout.t16 dvss 0.243993f
C785 xout.n0 dvss 2.4243f
C786 xout.t17 dvss 0.243993f
C787 xout.t15 dvss 0.243993f
C788 xout.n1 dvss 1.60432f
C789 xout.n2 dvss 6.32987f
C790 xout.t14 dvss 0.256529f
C791 xout.t19 dvss 0.243993f
C792 xout.n3 dvss 1.22843f
C793 xout.t12 dvss 0.256529f
C794 xout.t20 dvss 0.243993f
C795 xout.n4 dvss 1.23308f
C796 xout.n5 dvss 2.18555f
C797 xout.n6 dvss 8.527769f
C798 xout.n7 dvss 3.77761f
C799 xout.t9 dvss 0.243993f
C800 xout.t10 dvss 0.243993f
C801 xout.n8 dvss 1.27442f
C802 xout.n9 dvss 1.83376f
C803 xout.t11 dvss 0.243993f
C804 xout.t13 dvss 0.243993f
C805 xout.n10 dvss 1.43377f
C806 xout.n11 dvss 1.68066f
C807 xout.n12 dvss 1.24537f
C808 xout.t5 dvss 0.066767f
C809 xout.t7 dvss 0.066767f
C810 xout.n13 dvss 0.227228f
C811 xout.t3 dvss 0.066767f
C812 xout.t6 dvss 0.066767f
C813 xout.n14 dvss 0.217681f
C814 xout.t2 dvss 0.066767f
C815 xout.t4 dvss 0.066767f
C816 xout.n15 dvss 0.229174f
C817 xout.n16 dvss 4.49086f
C818 xout.t21 dvss 0.066767f
C819 xout.t22 dvss 0.066767f
C820 xout.n17 dvss 0.217681f
C821 xout.t1 dvss 0.066767f
C822 xout.t8 dvss 0.066767f
C823 xout.n18 dvss 0.149204f
C824 xout.n19 dvss 2.97025f
C825 xout.n20 dvss 3.47714f
C826 xout.n21 dvss 4.15788f
C827 xout.t0 dvss 0.091048f
C828 xout.n22 dvss 4.02374f
C829 xout.n23 dvss 0.626416f
C830 xout.n24 dvss 0.760656f
C831 xout.t25 dvss 1.61622f
C832 xout.t23 dvss 1.68073f
C833 xout.n25 dvss 1.04327f
C834 xout.n26 dvss 0.785936f
C835 xout.n27 dvss 8.087669f
C836 xout.n28 dvss 9.65943f
C837 xout.n29 dvss 1.9924f
C838 avdd_ip.t4 dvss 0.076964f
C839 avdd_ip.t3 dvss 0.076964f
C840 avdd_ip.n0 dvss 0.188642f
C841 avdd_ip.t6 dvss 0.076964f
C842 avdd_ip.t0 dvss 0.076964f
C843 avdd_ip.n1 dvss 0.199053f
C844 avdd_ip.t1 dvss 0.322205f
C845 avdd_ip.n2 dvss 26.4789f
C846 avdd_ip.t33 dvss 0.207758p
C847 avdd_ip.n3 dvss 43.6415f
C848 avdd_ip.n4 dvss 32.1711f
C849 avdd_ip.t30 dvss 13.0044f
C850 avdd_ip.n5 dvss 8.302629f
C851 avdd_ip.t31 dvss 13.0044f
C852 avdd_ip.n6 dvss 8.004399f
C853 avdd_ip.n7 dvss 10.5476f
C854 avdd_ip.t29 dvss 13.0044f
C855 avdd_ip.n8 dvss 11.6712f
C856 avdd_ip.t32 dvss 13.0044f
C857 avdd_ip.n9 dvss 11.647f
C858 avdd_ip.n10 dvss 11.3857f
C859 avdd_ip.n11 dvss 26.6555f
C860 avdd_ip.n12 dvss 7.31264f
C861 avdd_ip.n13 dvss 0.515994f
C862 avdd_ip.n14 dvss 4.47303f
C863 avdd_ip.n15 dvss 15.6554f
C864 avdd_ip.n16 dvss 15.6554f
C865 avdd_ip.t7 dvss 19.9269f
C866 avdd_ip.n17 dvss 1.66473f
C867 avdd_ip.t12 dvss 0.281261f
C868 avdd_ip.n18 dvss 5.57691f
C869 avdd_ip.t17 dvss 0.281261f
C870 avdd_ip.t18 dvss 0.281261f
C871 avdd_ip.n19 dvss 2.84698f
C872 avdd_ip.t14 dvss 0.281261f
C873 avdd_ip.t16 dvss 0.281261f
C874 avdd_ip.n20 dvss 1.65413f
C875 avdd_ip.n21 dvss 2.53602f
C876 avdd_ip.n22 dvss 6.96979f
C877 avdd_ip.t8 dvss 0.281261f
C878 avdd_ip.t9 dvss 0.281261f
C879 avdd_ip.t10 dvss 0.281261f
C880 avdd_ip.n23 dvss 2.35113f
C881 avdd_ip.n24 dvss 6.93137f
C882 avdd_ip.n25 dvss 4.04083f
C883 avdd_ip.n26 dvss 16.1821f
C884 avdd_ip.t22 dvss 0.281261f
C885 avdd_ip.t28 dvss 0.281261f
C886 avdd_ip.n27 dvss 2.77031f
C887 avdd_ip.t19 dvss 0.281261f
C888 avdd_ip.t27 dvss 0.281261f
C889 avdd_ip.n28 dvss 1.65277f
C890 avdd_ip.n29 dvss 2.61066f
C891 avdd_ip.n30 dvss 1.06102f
C892 avdd_ip.t20 dvss 0.281261f
C893 avdd_ip.n31 dvss 1.10166f
C894 avdd_ip.n32 dvss 1.22761f
C895 avdd_ip.t21 dvss 0.281261f
C896 avdd_ip.n33 dvss 0.364113f
C897 avdd_ip.t26 dvss 0.281261f
C898 avdd_ip.n34 dvss 0.527532f
C899 avdd_ip.n35 dvss 0.321659f
C900 avdd_ip.n36 dvss 0.936889f
C901 avdd_ip.t24 dvss 0.281261f
C902 avdd_ip.n37 dvss 1.28394f
C903 avdd_ip.t25 dvss 0.281261f
C904 avdd_ip.n38 dvss 1.40677f
C905 avdd_ip.t23 dvss 0.293118f
C906 avdd_ip.n39 dvss 1.03578f
C907 avdd_ip.n40 dvss 1.65219f
C908 avdd_ip.n41 dvss 12.23f
C909 avdd_ip.n42 dvss 6.74729f
C910 avdd_ip.n43 dvss 5.54535f
C911 avdd_ip.n44 dvss 12.9266f
C912 avdd_ip.n45 dvss 7.920741f
C913 avdd_ip.n46 dvss 8.73601f
C914 avdd_ip.n47 dvss 8.79801f
C915 avdd_ip.n48 dvss 8.79801f
C916 avdd_ip.n49 dvss 33.810898f
C917 avdd_ip.n50 dvss 7.28254f
C918 avdd_ip.n51 dvss 2.98117f
C919 avdd_ip.n52 dvss 8.78597f
C920 avdd_ip.n53 dvss 33.6251f
C921 avdd_ip.n54 dvss 33.810898f
C922 avdd_ip.n55 dvss 33.6251f
C923 avdd_ip.n56 dvss 8.78597f
C924 avdd_ip.n57 dvss 2.90114f
C925 avdd_ip.n58 dvss 0.083546f
C926 avdd_ip.n59 dvss 0.057941f
C927 avdd_ip.n60 dvss 0.058384f
C928 avdd_ip.n61 dvss 0.058384f
C929 avdd_ip.n62 dvss 0.067492f
C930 avdd_ip.n63 dvss 0.059867f
C931 avdd_ip.n64 dvss 0.283817f
C932 avdd_ip.t5 dvss 0.438989f
C933 avdd_ip.n67 dvss 0.283817f
C934 avdd_ip.n68 dvss 0.06656f
C935 avdd_ip.n69 dvss 0.062001f
C936 avdd_ip.n70 dvss 2.71257f
C937 avdd_ip.n71 dvss 0.079796f
C938 avdd_ip.n72 dvss 0.057936f
C939 avdd_ip.n73 dvss 0.058384f
C940 avdd_ip.t2 dvss 0.377338f
C941 avdd_ip.n74 dvss 0.06837f
C942 avdd_ip.n75 dvss 0.060427f
C943 avdd_ip.n76 dvss -23.5782f
C944 avdd_ip.n77 dvss 23.864698f
C945 avdd_ip.n78 dvss 0.058921f
C946 avdd_ip.n79 dvss 0.058384f
C947 avdd_ip.n81 dvss 0.283817f
C948 avdd_ip.n82 dvss 0.06656f
C949 avdd_ip.n83 dvss 0.062001f
C950 avdd_ip.n84 dvss 2.41392f
C951 avdd_ip.n85 dvss 3.17873f
C952 avdd_ip.n86 dvss 6.26191f
C953 avdd_ip.n87 dvss 28.2098f
C954 avdd_ip.n88 dvss 11.163099f
C955 avdd_ip.n89 dvss 2.27252f
C956 avdd_ip.n90 dvss 5.94738f
C957 avdd_ip.t13 dvss 0.281261f
C958 avdd_ip.t15 dvss 0.281261f
C959 avdd_ip.n91 dvss 2.34378f
C960 avdd_ip.n92 dvss 0.801311f
C961 avdd_ip.n93 dvss 1.44437f
C962 avdd_ip.t11 dvss 19.9269f
C963 avdd_ip.n94 dvss 17.055302f
C964 avdd_ip.n95 dvss 1.44437f
C965 avdd_ip.n96 dvss 2.92893f
C966 avdd_ip.n97 dvss 1.20647f
C967 avdd_ip.n98 dvss 0.016222f
C968 avdd_ip.n99 dvss 24.4049f
C969 ibias_ip.n0 dvss 4.75326f
C970 ibias_ip.n1 dvss 0.974101f
C971 ibias_ip.t13 dvss 0.653909f
C972 ibias_ip.t3 dvss 0.646782f
C973 ibias_ip.t4 dvss 0.082653f
C974 ibias_ip.t8 dvss 0.081898f
C975 ibias_ip.t7 dvss 0.644915f
C976 ibias_ip.t2 dvss 0.077591f
C977 ibias_ip.t1 dvss 0.650434f
C978 ibias_ip.t5 dvss 0.647233f
C979 ibias_ip.t11 dvss 0.653916f
C980 ibias_ip.t6 dvss 0.082116f
C981 ibias_ip.t10 dvss 0.082367f
C982 ibias_ip.t9 dvss 0.645067f
C983 ibias_ip.t12 dvss 0.646314f
C984 ibias_ip.t0 dvss 0.184945f
C985 standby_33.n0 dvss 7.35104f
C986 standby_33.t3 dvss 0.807828f
C987 standby_33.t4 dvss 1.63225f
C988 standby_33.t1 dvss 0.055479f
C989 standby_33.t2 dvss 0.055479f
C990 standby_33.n1 dvss 0.175556f
C991 standby_33.t0 dvss 0.068888f
C992 x7.ena_done_b.t1 dvss 0.054284f
C993 x7.ena_done_b.t0 dvss 0.068732f
C994 x7.ena_done_b.t3 dvss 0.033951f
C995 x7.ena_done_b.t2 dvss 0.02132f
C996 x7.ena_done_b.n0 dvss 0.045927f
C997 x7.ena_done_b.n1 dvss 0.058447f
C998 x7.ena_done_b.t4 dvss 0.018591f
C999 x7.ena_done_b.n2 dvss 0.053311f
C1000 x7.ena_done_b.t7 dvss 0.018802f
C1001 x7.ena_done_b.n3 dvss 0.05789f
C1002 x7.ena_done_b.n4 dvss 0.011573f
C1003 x7.ena_done_b.n5 dvss 0.060019f
C1004 x7.ena_done_b.t6 dvss 0.025304f
C1005 x7.ena_done_b.t5 dvss 0.027855f
C1006 x7.ena_done_b.n6 dvss 0.079658f
C1007 x7.ena_done_b.n7 dvss 1.96309f
C1008 x7.ena_done_b.n8 dvss 0.077694f
C1009 a_9120_n9346.t4 dvss 0.036089f
C1010 a_9120_n9346.t3 dvss 1.47746f
C1011 a_9120_n9346.n0 dvss 3.32132f
C1012 a_9120_n9346.t1 dvss 1.67898f
C1013 a_9120_n9346.t2 dvss 0.027167f
C1014 a_9120_n9346.n1 dvss 2.97825f
C1015 a_9120_n9346.n2 dvss 1.80939f
C1016 a_9120_n9346.t0 dvss 0.071336f
C1017 x7.x2.x4.RESET_B dvss 1.471743f
C1018 x7.x3.A1 dvss 0.02912f
C1019 standby_b.t1 dvss 2.65544f
C1020 standby_b.n0 dvss 0.147325f
C1021 x7.x2.x2.RESET_B dvss 0.028793f
C1022 x7.x2.x3.RESET_B dvss 0.028793f
C1023 standby_b.n1 dvss 3.12348f
C1024 x7.stby_b dvss 1.34845f
C1025 standby_b.t14 dvss 0.185493f
C1026 standby_b.t6 dvss 0.185354f
C1027 standby_b.n2 dvss 0.084915f
C1028 standby_b.n3 dvss 0.157601f
C1029 standby_b.t21 dvss 0.228815f
C1030 standby_b.t19 dvss 0.217171f
C1031 standby_b.n4 dvss 0.157601f
C1032 standby_b.n5 dvss 0.084915f
C1033 standby_b.t9 dvss 0.217171f
C1034 standby_b.n6 dvss 0.084915f
C1035 standby_b.t25 dvss 0.217171f
C1036 standby_b.n7 dvss 0.084915f
C1037 standby_b.n8 dvss 0.077844f
C1038 standby_b.t23 dvss 0.217171f
C1039 standby_b.n9 dvss 0.077734f
C1040 standby_b.n10 dvss 0.084915f
C1041 standby_b.n11 dvss 0.162102f
C1042 standby_b.t8 dvss 0.229503f
C1043 standby_b.t18 dvss 0.217171f
C1044 standby_b.n12 dvss 0.161693f
C1045 standby_b.n13 dvss 0.084915f
C1046 standby_b.t20 dvss 0.217171f
C1047 standby_b.n14 dvss 0.084915f
C1048 standby_b.t2 dvss 0.217171f
C1049 standby_b.n15 dvss 0.084915f
C1050 standby_b.n16 dvss 0.074529f
C1051 standby_b.t5 dvss 0.217171f
C1052 standby_b.n17 dvss 0.07464f
C1053 standby_b.t16 dvss 0.014102f
C1054 standby_b.n18 dvss 0.025012f
C1055 standby_b.t27 dvss 0.014102f
C1056 standby_b.n20 dvss 0.025012f
C1057 standby_b.t13 dvss 0.014102f
C1058 standby_b.n22 dvss 0.025012f
C1059 standby_b.t4 dvss 0.012275f
C1060 standby_b.n24 dvss 0.023944f
C1061 standby_b.t17 dvss 0.012275f
C1062 standby_b.n25 dvss 0.023944f
C1063 standby_b.t15 dvss 0.012275f
C1064 standby_b.n26 dvss 0.023944f
C1065 standby_b.t26 dvss 0.014675f
C1066 standby_b.n27 dvss 0.022499f
C1067 standby_b.t0 dvss 0.03467f
C1068 tail.n0 dvss 0.76343f
C1069 tail.n1 dvss 2.82244f
C1070 tail.t0 dvss 0.054705f
C1071 tail.t1 dvss 0.054705f
C1072 tail.n2 dvss 0.119757f
C1073 tail.t2 dvss 0.102772f
C1074 tail.t7 dvss 0.102893f
C1075 tail.t9 dvss 0.102832f
C1076 tail.t4 dvss 0.102832f
C1077 tail.t6 dvss 0.103102f
C1078 tail.t11 dvss 0.102562f
C1079 tail.t5 dvss 0.103102f
C1080 tail.t10 dvss 0.102562f
C1081 tail.n3 dvss 0.753923f
C1082 tail.t8 dvss 0.102998f
C1083 tail.t3 dvss 0.102668f
C1084 dvdd_ip.n0 dvss 0.04438f
C1085 dvdd_ip.n1 dvss 1.69588f
C1086 dvdd_ip.n2 dvss 9.84588f
C1087 dvdd_ip.n3 dvss 1.74493f
C1088 dvdd_ip.n4 dvss 0.43405f
C1089 dvdd_ip.n5 dvss 6.8385f
C1090 dvdd_ip.n6 dvss 0.547569f
C1091 dvdd_ip.n7 dvss 0.511986f
C1092 dvdd_ip.n8 dvss 16.501402f
C1093 dvdd_ip.n9 dvss 5.38917f
C1094 dvdd_ip.n10 dvss 0.857623f
C1095 dvdd_ip.n11 dvss 0.059854f
C1096 dvdd_ip.t56 dvss 0.407966p
C1097 dvdd_ip.n12 dvss 0.923802f
C1098 dvdd_ip.n13 dvss 0.626632f
C1099 dvdd_ip.n14 dvss 2.12851f
C1100 dvdd_ip.n15 dvss 1.11147f
C1101 dvdd_ip.n16 dvss 0.753616f
C1102 dvdd_ip.n17 dvss 0.856242f
C1103 dvdd_ip.n18 dvss 6.76846f
C1104 dvdd_ip.n19 dvss 0.352823f
C1105 dvdd_ip.n20 dvss 1.29174f
C1106 dvdd_ip.n21 dvss 0.411312f
C1107 dvdd_ip.n22 dvss 0.257212f
C1108 dvdd_ip.n23 dvss 1.14899f
C1109 dvdd_ip.n24 dvss 2.28269f
C1110 dvdd_ip.n25 dvss 0.853257f
C1111 dvdd_ip.n26 dvss 0.30361f
C1112 dvdd_ip.n27 dvss 1.71807f
C1113 dvdd_ip.n28 dvss 0.7202f
C1114 dvdd_ip.n30 dvss 0.162868f
C1115 dvdd_ip.n31 dvss 0.098289f
C1116 dvdd_ip.n32 dvss 0.098289f
C1117 dvdd_ip.t16 dvss 1.16977f
C1118 dvdd_ip.n33 dvss 0.088581f
C1119 dvdd_ip.n35 dvss 0.836093f
C1120 dvdd_ip.n36 dvss 0.098289f
C1121 dvdd_ip.n38 dvss 0.836093f
C1122 dvdd_ip.n39 dvss 0.105976f
C1123 dvdd_ip.n40 dvss 1.54065f
C1124 dvdd_ip.n41 dvss 2.06853f
C1125 dvdd_ip.n42 dvss 2.06853f
C1126 dvdd_ip.n43 dvss 7.93383f
C1127 dvdd_ip.t21 dvss 0.104505f
C1128 dvdd_ip.n45 dvss 0.067374f
C1129 dvdd_ip.n46 dvss 0.058872f
C1130 dvdd_ip.n47 dvss 0.058872f
C1131 dvdd_ip.n48 dvss 0.506053f
C1132 dvdd_ip.t14 dvss 0.013379f
C1133 dvdd_ip.n49 dvss 0.242497f
C1134 dvdd_ip.n50 dvss 0.332713f
C1135 dvdd_ip.t51 dvss 0.053917f
C1136 dvdd_ip.t35 dvss 0.053871f
C1137 dvdd_ip.t33 dvss 0.053983f
C1138 dvdd_ip.t45 dvss 0.05381f
C1139 dvdd_ip.t43 dvss 0.081434f
C1140 dvdd_ip.t44 dvss 0.051849f
C1141 dvdd_ip.n51 dvss 0.496721f
C1142 dvdd_ip.t48 dvss 0.053917f
C1143 dvdd_ip.t52 dvss 0.051849f
C1144 dvdd_ip.t28 dvss 0.051849f
C1145 dvdd_ip.t46 dvss 0.05446f
C1146 dvdd_ip.t30 dvss 0.051849f
C1147 dvdd_ip.n52 dvss 0.366284f
C1148 dvdd_ip.t31 dvss 0.051849f
C1149 dvdd_ip.n53 dvss 0.279183f
C1150 dvdd_ip.t39 dvss 0.05446f
C1151 dvdd_ip.t49 dvss 0.051849f
C1152 dvdd_ip.n54 dvss 0.366284f
C1153 dvdd_ip.t50 dvss 0.051849f
C1154 dvdd_ip.n55 dvss 0.279183f
C1155 dvdd_ip.t17 dvss 0.013379f
C1156 dvdd_ip.n57 dvss 0.889873f
C1157 dvdd_ip.n58 dvss 0.249178f
C1158 dvdd_ip.n59 dvss 0.659876f
C1159 dvdd_ip.t1 dvss 0.013379f
C1160 dvdd_ip.n61 dvss 0.501881f
C1161 dvdd_ip.n62 dvss 0.776954f
C1162 dvdd_ip.t0 dvss 1.29168f
C1163 dvdd_ip.n64 dvss 0.09647f
C1164 dvdd_ip.n65 dvss 0.776954f
C1165 dvdd_ip.n66 dvss 0.106044f
C1166 dvdd_ip.n67 dvss 0.674388f
C1167 dvdd_ip.n68 dvss 0.755374f
C1168 dvdd_ip.n69 dvss 0.092376f
C1169 dvdd_ip.n70 dvss 1.14551f
C1170 dvdd_ip.n71 dvss 1.14551f
C1171 dvdd_ip.t23 dvss 1.45965f
C1172 dvdd_ip.t19 dvss 1.18355f
C1173 dvdd_ip.n72 dvss 0.235608f
C1174 dvdd_ip.t18 dvss 1.45965f
C1175 dvdd_ip.t22 dvss 1.18355f
C1176 dvdd_ip.n73 dvss 0.789036f
C1177 dvdd_ip.n74 dvss 0.235608f
C1178 dvdd_ip.t41 dvss 0.05446f
C1179 dvdd_ip.t26 dvss 0.051849f
C1180 dvdd_ip.n75 dvss 0.366284f
C1181 dvdd_ip.t25 dvss 0.051849f
C1182 dvdd_ip.n76 dvss 0.279183f
C1183 dvdd_ip.t47 dvss 0.054399f
C1184 dvdd_ip.t37 dvss 0.051849f
C1185 dvdd_ip.n77 dvss 0.364367f
C1186 dvdd_ip.t36 dvss 0.051849f
C1187 dvdd_ip.n78 dvss 0.279183f
C1188 dvdd_ip.n79 dvss 0.975269f
C1189 dvdd_ip.t24 dvss 1.57973f
C1190 dvdd_ip.t40 dvss 1.93128f
C1191 dvdd_ip.t32 dvss 1.93128f
C1192 dvdd_ip.t34 dvss 1.44846f
C1193 dvdd_ip.n80 dvss 0.96564f
C1194 dvdd_ip.t42 dvss 1.44846f
C1195 dvdd_ip.t27 dvss 1.93128f
C1196 dvdd_ip.t38 dvss 1.93128f
C1197 dvdd_ip.t29 dvss 1.57973f
C1198 dvdd_ip.n81 dvss 0.973802f
C1199 dvdd_ip.n82 dvss 0.463049f
C1200 dvdd_ip.n85 dvss 0.458062f
C1201 dvdd_ip.n86 dvss 0.568458f
C1202 dvdd_ip.n87 dvss 0.300827f
C1203 dvdd_ip.n88 dvss 0.077314f
C1204 dvdd_ip.n89 dvss 0.033341f
C1205 dvdd_ip.n90 dvss 0.362868f
C1206 dvdd_ip.t7 dvss 0.378798f
C1207 dvdd_ip.n91 dvss 0.24424f
C1208 dvdd_ip.t9 dvss 0.378798f
C1209 dvdd_ip.n92 dvss 0.362868f
C1210 dvdd_ip.n93 dvss 0.54101f
C1211 dvdd_ip.t20 dvss 0.866692f
C1212 dvdd_ip.n95 dvss 0.067374f
C1213 dvdd_ip.n96 dvss 0.54101f
C1214 dvdd_ip.n97 dvss 1.79645f
C1215 dvdd_ip.n98 dvss 0.822077f
C1216 dvdd_ip.n99 dvss 2.06224f
C1217 dvdd_ip.n100 dvss 7.83594f
C1218 dvdd_ip.n101 dvss 7.93383f
C1219 dvdd_ip.n102 dvss 7.83594f
C1220 dvdd_ip.n103 dvss 2.06224f
C1221 dvdd_ip.n104 dvss 0.976313f
C1222 dvdd_ip.n105 dvss 0.638912f
C1223 dvdd_ip.t11 dvss 0.028672f
C1224 dvdd_ip.t53 dvss 0.028672f
C1225 dvdd_ip.n106 dvss 0.068783f
C1226 dvdd_ip.t6 dvss 0.028672f
C1227 dvdd_ip.t54 dvss 0.028672f
C1228 dvdd_ip.n107 dvss 0.068762f
C1229 dvdd_ip.t3 dvss 0.028672f
C1230 dvdd_ip.t55 dvss 0.028672f
C1231 dvdd_ip.n108 dvss 0.068783f
C1232 dvdd_ip.t5 dvss 0.028672f
C1233 dvdd_ip.t12 dvss 0.028672f
C1234 dvdd_ip.n109 dvss 0.068762f
C1235 dvdd_ip.t4 dvss 0.028672f
C1236 dvdd_ip.t2 dvss 0.028672f
C1237 dvdd_ip.n110 dvss 0.068762f
C1238 dvdd_ip.n111 dvss 12.7858f
C1239 vbp.n0 dvss 0.179072f
C1240 vbp.n1 dvss 0.347213f
C1241 vbp.n2 dvss 0.361375f
C1242 vbp.n3 dvss 6.70539f
C1243 vbp.n4 dvss 0.178688f
C1244 vbp.n5 dvss 0.347213f
C1245 vbp.n6 dvss 0.345626f
C1246 vbp.n7 dvss 0.353693f
C1247 vbp.t13 dvss 0.876014f
C1248 vbp.t5 dvss 0.946258f
C1249 vbp.t2 dvss 0.114991f
C1250 vbp.t9 dvss 0.880979f
C1251 vbp.t7 dvss 0.853138f
C1252 vbp.t12 dvss 0.876026f
C1253 vbp.t17 dvss 0.946667f
C1254 vbp.t11 dvss 1.12602f
C1255 vbp.t14 dvss 0.854726f
C1256 vbp.t4 dvss 0.854724f
C1257 vbp.t1 dvss 0.908023f
C1258 vbp.t15 dvss 1.12462f
C1259 vbp.t8 dvss 0.853138f
C1260 vbp.t16 dvss 0.891507f
C1261 vbp.t6 dvss 0.891734f
C1262 vbp.t10 dvss 0.871833f
C1263 vbp.t3 dvss 0.8852f
C1264 vbp.t0 dvss 0.123277f
C1265 vbreg.n0 dvss 3.5606f
C1266 vbreg.n1 dvss 0.713612f
C1267 vbreg.n2 dvss 0.583542f
C1268 vbreg.n3 dvss 3.65749f
C1269 vbreg.n4 dvss 1.34473f
C1270 vbreg.n5 dvss 3.556f
C1271 vbreg.n6 dvss 0.687636f
C1272 vbreg.n7 dvss 0.582626f
C1273 vbreg.n8 dvss 1.213f
C1274 vbreg.n9 dvss 2.841f
C1275 vbreg.n10 dvss 0.583359f
C1276 vbreg.n11 dvss 2.61721f
C1277 vbreg.n12 dvss 0.592924f
C1278 vbreg.n14 dvss 0.594449f
C1279 vbreg.n15 dvss 0.931401f
C1280 vbreg.n16 dvss 0.933049f
C1281 vbreg.n17 dvss 0.404251f
C1282 vbreg.n18 dvss 0.933049f
C1283 vbreg.t11 dvss 1.20117f
C1284 vbreg.n19 dvss 0.931401f
C1285 vbreg.t4 dvss 0.23921f
C1286 vbreg.n20 dvss 1.79539f
C1287 vbreg.n21 dvss 12.184299f
C1288 vbreg.t6 dvss 0.228907f
C1289 vbreg.n22 dvss 1.25884f
C1290 vbreg.n23 dvss 0.616431f
C1291 vbreg.t7 dvss 1.20117f
C1292 vbreg.n24 dvss 0.662505f
C1293 vbreg.t19 dvss 1.20117f
C1294 vbreg.n25 dvss 0.404251f
C1295 vbreg.n26 dvss 0.400957f
C1296 vbreg.t20 dvss 1.20117f
C1297 vbreg.t18 dvss 1.20117f
C1298 vbreg.t15 dvss 1.20117f
C1299 vbreg.n27 dvss 1.00001f
C1300 vbreg.t16 dvss 1.20117f
C1301 vbreg.n28 dvss 0.685977f
C1302 vbreg.n29 dvss 0.530447f
C1303 vbreg.n30 dvss 0.404251f
C1304 vbreg.n31 dvss 0.710976f
C1305 vbreg.t10 dvss 1.21612f
C1306 vbreg.t13 dvss 1.20117f
C1307 vbreg.n32 dvss 1.00001f
C1308 vbreg.n33 dvss 0.085368f
C1309 vbreg.t12 dvss 1.20117f
C1310 vbreg.n34 dvss 1.00001f
C1311 vbreg.t14 dvss 1.20117f
C1312 vbreg.n35 dvss 0.692695f
C1313 vbreg.n36 dvss 1.00001f
C1314 vbreg.t9 dvss 1.20117f
C1315 vbreg.n37 dvss 0.530447f
C1316 vbreg.n38 dvss 0.661796f
C1317 vbreg.t17 dvss 1.20117f
C1318 vbreg.n39 dvss 1.00001f
C1319 vbreg.n40 dvss 0.168268f
C1320 vbreg.n41 dvss 1.00001f
C1321 vbreg.t8 dvss 0.228404f
C1322 vbreg.n42 dvss 0.815331f
C1323 vbreg.n43 dvss 0.528798f
C1324 vbreg.n44 dvss 0.404251f
C1325 vbreg.n45 dvss 1.00001f
C1326 vbreg.t22 dvss 1.20117f
C1327 vbreg.t24 dvss 1.20117f
C1328 vbreg.t25 dvss 1.20117f
C1329 vbreg.n46 dvss 1.00001f
C1330 vbreg.t21 dvss 1.20117f
C1331 vbreg.n47 dvss 0.531546f
C1332 vbreg.t23 dvss 1.21618f
C1333 vbreg.n48 dvss 1.00001f
C1334 vbreg.n49 dvss 0.085917f
C1335 vbreg.n50 dvss 1.30967f
C1336 vbreg.n51 dvss 0.705366f
C1337 vbreg.n52 dvss 0.531546f
C1338 vbreg.n53 dvss 0.404251f
C1339 vbreg.n54 dvss 0.527699f
C1340 vbreg.n55 dvss 0.527699f
C1341 vbreg.n56 dvss 0.404251f
C1342 vbreg.n57 dvss 0.55298f
C1343 vbreg.t0 dvss 0.214967f
C1344 vbreg.t5 dvss 0.228223f
C1345 vbreg.t1 dvss 0.268952f
C1346 vbreg.t3 dvss 0.218294f
C1347 vbreg.t2 dvss 0.138373f
C1348 icnode.t1 dvss 80.4574f
C1349 icnode.t0 dvss 0.042604f
C1350 ena_ip.n0 dvss 0.052729f
C1351 ena_ip.t0 dvss 0.038646f
C1352 ena_ip.n1 dvss 0.299073f
C1353 ena_ip.t14 dvss 0.312422f
C1354 ena_ip.t17 dvss 0.312179f
C1355 ena_ip.n2 dvss 0.262394f
C1356 ena_ip.n3 dvss 1.2068f
C1357 ena_ip.t2 dvss 0.357117f
C1358 ena_ip.t12 dvss 0.343909f
C1359 ena_ip.t18 dvss 0.013233f
C1360 ena_ip.t16 dvss 0.021012f
C1361 ena_ip.n4 dvss 0.040986f
C1362 ena_ip.t15 dvss 0.010303f
C1363 ena_ip.t4 dvss 0.024139f
C1364 ena_ip.n7 dvss 0.042815f
C1365 ena_ip.t10 dvss 0.013233f
C1366 ena_ip.t8 dvss 0.021012f
C1367 ena_ip.n8 dvss 0.040986f
C1368 ena_ip.t5 dvss 0.010303f
C1369 ena_ip.t13 dvss 0.024139f
C1370 ena_ip.n11 dvss 0.042815f
C1371 ena_ip.t9 dvss 0.013233f
C1372 ena_ip.t6 dvss 0.021012f
C1373 ena_ip.n12 dvss 0.040986f
C1374 ena_ip.t3 dvss 0.010303f
C1375 ena_ip.t7 dvss 0.024139f
C1376 ena_ip.n15 dvss 0.042815f
C1377 ena_ip.t19 dvss 0.025235f
C1378 ena_ip.t11 dvss 0.015832f
C1379 ena_ip.n16 dvss 0.036079f
C1380 ena_ip.n17 dvss 0.024525f
C1381 ena_ip.n18 dvss 0.153572f
C1382 ena_ip.t1 dvss 0.026873f
C1383 dvdd.t37 dvss 0.010234f
C1384 dvdd.t39 dvss 0.010234f
C1385 dvdd.n0 dvss 0.232259f
C1386 dvdd.n1 dvss 0.072245f
C1387 dvdd.n3 dvss 0.016615f
C1388 dvdd.n4 dvss 0.115145f
C1389 dvdd.n5 dvss 0.115145f
C1390 dvdd.t108 dvss 0.054261f
C1391 dvdd.t148 dvss 0.018343f
C1392 dvdd.n9 dvss 0.013679f
C1393 dvdd.n11 dvss 0.04491f
C1394 dvdd.n14 dvss 0.023525f
C1395 dvdd.n15 dvss 0.02803f
C1396 dvdd.n16 dvss 0.018576f
C1397 dvdd.t127 dvss 0.054261f
C1398 dvdd.t114 dvss 0.018343f
C1399 dvdd.n18 dvss 0.04491f
C1400 dvdd.n23 dvss 0.013679f
C1401 dvdd.n25 dvss 0.028928f
C1402 dvdd.n26 dvss 0.011776f
C1403 dvdd.n27 dvss 0.115145f
C1404 dvdd.n28 dvss 0.016615f
C1405 dvdd.n29 dvss 0.115145f
C1406 dvdd.n30 dvss 0.016628f
C1407 dvdd.t38 dvss 0.165693f
C1408 dvdd.n33 dvss 0.016628f
C1409 dvdd.n34 dvss 0.011776f
C1410 dvdd.n38 dvss 0.474106f
C1411 dvdd.n39 dvss 0.250318f
C1412 dvdd.n41 dvss 0.011776f
C1413 dvdd.n42 dvss 0.016628f
C1414 dvdd.t36 dvss 0.165693f
C1415 dvdd.n45 dvss 0.016628f
C1416 dvdd.n46 dvss 0.011776f
C1417 dvdd.n48 dvss 0.09808f
C1418 dvdd.n49 dvss 1.84984f
C1419 dvdd.t175 dvss 3.84176f
C1420 dvdd.n50 dvss 3.23391f
C1421 dvdd.n51 dvss 0.770276f
C1422 dvdd.n53 dvss 0.031969f
C1423 dvdd.n54 dvss 0.031969f
C1424 dvdd.n55 dvss 0.031969f
C1425 dvdd.n56 dvss 0.013375f
C1426 dvdd.n69 dvss 0.018583f
C1427 dvdd.n73 dvss 0.012437f
C1428 dvdd.n90 dvss 0.018583f
C1429 dvdd.n94 dvss 0.012437f
C1430 dvdd.n111 dvss 0.018583f
C1431 dvdd.n115 dvss 0.012437f
C1432 dvdd.n125 dvss 0.015342f
C1433 dvdd.n131 dvss 0.025982f
C1434 dvdd.n144 dvss 0.013272f
C1435 dvdd.n151 dvss 0.013047f
C1436 dvdd.n156 dvss 0.016487f
C1437 dvdd.n163 dvss 0.015342f
C1438 dvdd.n169 dvss 0.025982f
C1439 dvdd.n182 dvss 0.013272f
C1440 dvdd.n189 dvss 0.013047f
C1441 dvdd.n194 dvss 0.016487f
C1442 dvdd.n201 dvss 0.015342f
C1443 dvdd.n207 dvss 0.025982f
C1444 dvdd.n220 dvss 0.013272f
C1445 dvdd.n227 dvss 0.013047f
C1446 dvdd.n232 dvss 0.016487f
C1447 dvdd.n239 dvss 0.037534f
C1448 dvdd.t76 dvss 0.052411f
C1449 dvdd.t45 dvss 0.026976f
C1450 dvdd.t47 dvss 0.021118f
C1451 dvdd.t10 dvss 0.039f
C1452 dvdd.t137 dvss 0.029134f
C1453 dvdd.t14 dvss 0.043779f
C1454 dvdd.t92 dvss 0.041929f
C1455 dvdd.t124 dvss 0.025897f
C1456 dvdd.t44 dvss 0.017573f
C1457 dvdd.n246 dvss 0.045107f
C1458 dvdd.n254 dvss 0.010792f
C1459 dvdd.n257 dvss 0.013038f
C1460 dvdd.n265 dvss 0.013229f
C1461 dvdd.n267 dvss 0.032824f
C1462 dvdd.n269 dvss 0.071001f
C1463 dvdd.t74 dvss 0.045391f
C1464 dvdd.t26 dvss 0.065777f
C1465 dvdd.t33 dvss 0.084259f
C1466 dvdd.n270 dvss 0.072157f
C1467 dvdd.t2 dvss 0.040499f
C1468 dvdd.t12 dvss 0.095403f
C1469 dvdd.t18 dvss 0.097578f
C1470 dvdd.t98 dvss 0.051915f
C1471 dvdd.t63 dvss 0.064961f
C1472 dvdd.t31 dvss 0.064418f
C1473 dvdd.t106 dvss 0.07991f
C1474 dvdd.t8 dvss 0.080454f
C1475 dvdd.t110 dvss 0.050284f
C1476 dvdd.t97 dvss 0.046207f
C1477 dvdd.t117 dvss 0.052187f
C1478 dvdd.t90 dvss 0.052187f
C1479 dvdd.t125 dvss 0.067408f
C1480 dvdd.t66 dvss 0.104101f
C1481 dvdd.t64 dvss 0.08589f
C1482 dvdd.t133 dvss 0.067408f
C1483 dvdd.n271 dvss 0.070798f
C1484 dvdd.t20 dvss 0.040499f
C1485 dvdd.t4 dvss 0.095403f
C1486 dvdd.t22 dvss 0.097578f
C1487 dvdd.t159 dvss 0.051915f
C1488 dvdd.t7 dvss 0.064961f
C1489 dvdd.t152 dvss 0.064418f
C1490 dvdd.t16 dvss 0.07991f
C1491 dvdd.t0 dvss 0.080454f
C1492 dvdd.t6 dvss 0.050284f
C1493 dvdd.t96 dvss 0.046207f
C1494 dvdd.t120 dvss 0.052187f
C1495 dvdd.t72 dvss 0.052187f
C1496 dvdd.t111 dvss 0.067408f
C1497 dvdd.t145 dvss 0.104101f
C1498 dvdd.t135 dvss 0.08589f
C1499 dvdd.t129 dvss 0.067408f
C1500 dvdd.n272 dvss 0.070798f
C1501 dvdd.t93 dvss 0.040499f
C1502 dvdd.t81 dvss 0.095403f
C1503 dvdd.t24 dvss 0.097578f
C1504 dvdd.t158 dvss 0.051915f
C1505 dvdd.t142 dvss 0.064961f
C1506 dvdd.t49 dvss 0.064418f
C1507 dvdd.t61 dvss 0.07991f
C1508 dvdd.t28 dvss 0.080454f
C1509 dvdd.t57 dvss 0.050284f
C1510 dvdd.t83 dvss 0.046207f
C1511 dvdd.t84 dvss 0.052187f
C1512 dvdd.t102 dvss 0.052187f
C1513 dvdd.t86 dvss 0.067408f
C1514 dvdd.t58 dvss 0.104101f
C1515 dvdd.t100 dvss 0.08589f
C1516 dvdd.t52 dvss 0.095845f
C1517 dvdd.n273 dvss 0.098023f
C1518 dvdd.n274 dvss 6.549109f
C1519 dvdd.n275 dvss 9.83819f
C1520 dvdd.t178 dvss 3.84176f
C1521 dvdd.n276 dvss 6.8075f
C1522 dvdd.t177 dvss 3.84176f
C1523 dvdd.n277 dvss 3.73525f
C1524 dvdd.t176 dvss 3.84176f
C1525 dvdd.n278 dvss 3.61309f
C1526 dvdd.n279 dvss 2.5797f
C1527 dvdd.n280 dvss 0.391121f
C1528 dvdd.t172 dvss 0.011141f
C1529 dvdd.t56 dvss 0.011141f
C1530 dvdd.n281 dvss 0.026719f
C1531 dvdd.t41 dvss 0.011141f
C1532 dvdd.t71 dvss 0.011141f
C1533 dvdd.n282 dvss 0.026719f
C1534 dvdd.n283 dvss 0.052335f
C1535 dvdd.t170 dvss 0.040608f
C1536 dvdd.n284 dvss 0.048007f
C1537 dvdd.n285 dvss 0.047867f
C1538 dvdd.n286 dvss 0.047867f
C1539 dvdd.t69 dvss 0.040608f
C1540 dvdd.t80 dvss 0.011141f
C1541 dvdd.t78 dvss 0.011141f
C1542 dvdd.n287 dvss 0.026719f
C1543 dvdd.t168 dvss 0.011141f
C1544 dvdd.t43 dvss 0.011141f
C1545 dvdd.n288 dvss 0.026719f
C1546 dvdd.n289 dvss 0.466772f
C1547 dvdd.n290 dvss 0.870378f
C1548 dvdd.n291 dvss 0.243449f
C1549 dvdd.n292 dvss 0.211336f
C1550 dvdd.t68 dvss 0.223235f
C1551 dvdd.t79 dvss 0.187866f
C1552 dvdd.t77 dvss 0.187866f
C1553 dvdd.t167 dvss 0.187866f
C1554 dvdd.t42 dvss 0.140899f
C1555 dvdd.n293 dvss 0.093933f
C1556 dvdd.t171 dvss 0.140899f
C1557 dvdd.t55 dvss 0.187866f
C1558 dvdd.t40 dvss 0.187866f
C1559 dvdd.t70 dvss 0.187866f
C1560 dvdd.t169 dvss 0.223235f
C1561 dvdd.n294 dvss 0.211336f
C1562 dvdd.n295 dvss 0.256347f
C1563 dvdd.n296 dvss 0.77501f
C1564 dvdd.n297 dvss 0.375275f
C1565 dvdd.n298 dvss 0.088595f
C1566 x7.stby_done_b.t1 dvss 0.057884f
C1567 x7.stby_done_b.n0 dvss 1.92933f
C1568 x7.stby_done_b.t5 dvss 0.028593f
C1569 x7.stby_done_b.t7 dvss 0.017955f
C1570 x7.stby_done_b.n1 dvss 0.038437f
C1571 x7.stby_done_b.n2 dvss 0.05998f
C1572 x7.stby_done_b.t4 dvss 0.015834f
C1573 x7.stby_done_b.n3 dvss 0.048959f
C1574 x7.stby_done_b.t3 dvss 0.015657f
C1575 x7.stby_done_b.n4 dvss 0.044896f
C1576 x7.stby_done_b.n5 dvss 0.047435f
C1577 x7.stby_done_b.t2 dvss 0.02131f
C1578 x7.stby_done_b.t6 dvss 0.023458f
C1579 x7.stby_done_b.n6 dvss 0.067085f
C1580 x7.stby_done_b.n7 dvss 1.67028f
C1581 x7.stby_done_b.n8 dvss 0.069954f
C1582 x7.stby_done_b.t0 dvss 0.043534f
.ends

