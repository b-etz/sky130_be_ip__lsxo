magic
tech sky130A
magscale 1 2
timestamp 1712854380
<< nwell >>
rect -996 -383 996 383
<< pmos >>
rect -800 64 800 164
rect -800 -164 800 -64
<< pdiff >>
rect -858 152 -800 164
rect -858 76 -846 152
rect -812 76 -800 152
rect -858 64 -800 76
rect 800 152 858 164
rect 800 76 812 152
rect 846 76 858 152
rect 800 64 858 76
rect -858 -76 -800 -64
rect -858 -152 -846 -76
rect -812 -152 -800 -76
rect -858 -164 -800 -152
rect 800 -76 858 -64
rect 800 -152 812 -76
rect 846 -152 858 -76
rect 800 -164 858 -152
<< pdiffc >>
rect -846 76 -812 152
rect 812 76 846 152
rect -846 -152 -812 -76
rect 812 -152 846 -76
<< nsubdiff >>
rect -960 313 -864 347
rect 864 313 960 347
rect -960 251 -926 313
rect 926 251 960 313
rect -960 -313 -926 -251
rect 926 -313 960 -251
rect -960 -347 -864 -313
rect 864 -347 960 -313
<< nsubdiffcont >>
rect -864 313 864 347
rect -960 -251 -926 251
rect 926 -251 960 251
rect -864 -347 864 -313
<< poly >>
rect -800 245 800 261
rect -800 211 -784 245
rect 784 211 800 245
rect -800 164 800 211
rect -800 17 800 64
rect -800 -17 -784 17
rect 784 -17 800 17
rect -800 -64 800 -17
rect -800 -211 800 -164
rect -800 -245 -784 -211
rect 784 -245 800 -211
rect -800 -261 800 -245
<< polycont >>
rect -784 211 784 245
rect -784 -17 784 17
rect -784 -245 784 -211
<< locali >>
rect -960 313 -864 347
rect 864 313 960 347
rect -960 251 -926 313
rect 926 251 960 313
rect -800 211 -784 245
rect 784 211 800 245
rect -846 152 -812 168
rect -846 60 -812 76
rect 812 152 846 168
rect 812 60 846 76
rect -800 -17 -784 17
rect 784 -17 800 17
rect -846 -76 -812 -60
rect -846 -168 -812 -152
rect 812 -76 846 -60
rect 812 -168 846 -152
rect -800 -245 -784 -211
rect 784 -245 800 -211
rect -960 -313 -926 -251
rect 926 -313 960 -251
rect -960 -347 -864 -313
rect 864 -347 960 -313
<< viali >>
rect -784 211 784 245
rect -846 76 -812 152
rect 812 76 846 152
rect -784 -17 784 17
rect -846 -152 -812 -76
rect 812 -152 846 -76
rect -784 -245 784 -211
<< metal1 >>
rect -796 245 796 251
rect -796 211 -784 245
rect 784 211 796 245
rect -796 205 796 211
rect -852 152 -806 164
rect -852 76 -846 152
rect -812 76 -806 152
rect -852 64 -806 76
rect 806 152 852 164
rect 806 76 812 152
rect 846 76 852 152
rect 806 64 852 76
rect -796 17 796 23
rect -796 -17 -784 17
rect 784 -17 796 17
rect -796 -23 796 -17
rect -852 -76 -806 -64
rect -852 -152 -846 -76
rect -812 -152 -806 -76
rect -852 -164 -806 -152
rect 806 -76 852 -64
rect 806 -152 812 -76
rect 846 -152 852 -76
rect 806 -164 852 -152
rect -796 -211 796 -205
rect -796 -245 -784 -211
rect 784 -245 796 -211
rect -796 -251 796 -245
<< properties >>
string FIXED_BBOX -943 -330 943 330
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 8 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
