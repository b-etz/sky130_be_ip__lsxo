magic
tech sky130A
magscale 1 2
timestamp 1712853061
<< nwell >>
rect -1312 -737 1312 737
<< pmos >>
rect -1116 118 -716 518
rect -658 118 -258 518
rect -200 118 200 518
rect 258 118 658 518
rect 716 118 1116 518
rect -1116 -518 -716 -118
rect -658 -518 -258 -118
rect -200 -518 200 -118
rect 258 -518 658 -118
rect 716 -518 1116 -118
<< pdiff >>
rect -1174 506 -1116 518
rect -1174 130 -1162 506
rect -1128 130 -1116 506
rect -1174 118 -1116 130
rect -716 506 -658 518
rect -716 130 -704 506
rect -670 130 -658 506
rect -716 118 -658 130
rect -258 506 -200 518
rect -258 130 -246 506
rect -212 130 -200 506
rect -258 118 -200 130
rect 200 506 258 518
rect 200 130 212 506
rect 246 130 258 506
rect 200 118 258 130
rect 658 506 716 518
rect 658 130 670 506
rect 704 130 716 506
rect 658 118 716 130
rect 1116 506 1174 518
rect 1116 130 1128 506
rect 1162 130 1174 506
rect 1116 118 1174 130
rect -1174 -130 -1116 -118
rect -1174 -506 -1162 -130
rect -1128 -506 -1116 -130
rect -1174 -518 -1116 -506
rect -716 -130 -658 -118
rect -716 -506 -704 -130
rect -670 -506 -658 -130
rect -716 -518 -658 -506
rect -258 -130 -200 -118
rect -258 -506 -246 -130
rect -212 -506 -200 -130
rect -258 -518 -200 -506
rect 200 -130 258 -118
rect 200 -506 212 -130
rect 246 -506 258 -130
rect 200 -518 258 -506
rect 658 -130 716 -118
rect 658 -506 670 -130
rect 704 -506 716 -130
rect 658 -518 716 -506
rect 1116 -130 1174 -118
rect 1116 -506 1128 -130
rect 1162 -506 1174 -130
rect 1116 -518 1174 -506
<< pdiffc >>
rect -1162 130 -1128 506
rect -704 130 -670 506
rect -246 130 -212 506
rect 212 130 246 506
rect 670 130 704 506
rect 1128 130 1162 506
rect -1162 -506 -1128 -130
rect -704 -506 -670 -130
rect -246 -506 -212 -130
rect 212 -506 246 -130
rect 670 -506 704 -130
rect 1128 -506 1162 -130
<< nsubdiff >>
rect -1276 667 -1180 701
rect 1180 667 1276 701
rect -1276 605 -1242 667
rect 1242 605 1276 667
rect -1276 -667 -1242 -605
rect 1242 -667 1276 -605
rect -1276 -701 -1180 -667
rect 1180 -701 1276 -667
<< nsubdiffcont >>
rect -1180 667 1180 701
rect -1276 -605 -1242 605
rect 1242 -605 1276 605
rect -1180 -701 1180 -667
<< poly >>
rect -1116 599 -716 615
rect -1116 565 -1100 599
rect -732 565 -716 599
rect -1116 518 -716 565
rect -658 599 -258 615
rect -658 565 -642 599
rect -274 565 -258 599
rect -658 518 -258 565
rect -200 599 200 615
rect -200 565 -184 599
rect 184 565 200 599
rect -200 518 200 565
rect 258 599 658 615
rect 258 565 274 599
rect 642 565 658 599
rect 258 518 658 565
rect 716 599 1116 615
rect 716 565 732 599
rect 1100 565 1116 599
rect 716 518 1116 565
rect -1116 71 -716 118
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -1116 21 -716 37
rect -658 71 -258 118
rect -658 37 -642 71
rect -274 37 -258 71
rect -658 21 -258 37
rect -200 71 200 118
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect 258 71 658 118
rect 258 37 274 71
rect 642 37 658 71
rect 258 21 658 37
rect 716 71 1116 118
rect 716 37 732 71
rect 1100 37 1116 71
rect 716 21 1116 37
rect -1116 -37 -716 -21
rect -1116 -71 -1100 -37
rect -732 -71 -716 -37
rect -1116 -118 -716 -71
rect -658 -37 -258 -21
rect -658 -71 -642 -37
rect -274 -71 -258 -37
rect -658 -118 -258 -71
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -118 200 -71
rect 258 -37 658 -21
rect 258 -71 274 -37
rect 642 -71 658 -37
rect 258 -118 658 -71
rect 716 -37 1116 -21
rect 716 -71 732 -37
rect 1100 -71 1116 -37
rect 716 -118 1116 -71
rect -1116 -565 -716 -518
rect -1116 -599 -1100 -565
rect -732 -599 -716 -565
rect -1116 -615 -716 -599
rect -658 -565 -258 -518
rect -658 -599 -642 -565
rect -274 -599 -258 -565
rect -658 -615 -258 -599
rect -200 -565 200 -518
rect -200 -599 -184 -565
rect 184 -599 200 -565
rect -200 -615 200 -599
rect 258 -565 658 -518
rect 258 -599 274 -565
rect 642 -599 658 -565
rect 258 -615 658 -599
rect 716 -565 1116 -518
rect 716 -599 732 -565
rect 1100 -599 1116 -565
rect 716 -615 1116 -599
<< polycont >>
rect -1100 565 -732 599
rect -642 565 -274 599
rect -184 565 184 599
rect 274 565 642 599
rect 732 565 1100 599
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect -1100 -71 -732 -37
rect -642 -71 -274 -37
rect -184 -71 184 -37
rect 274 -71 642 -37
rect 732 -71 1100 -37
rect -1100 -599 -732 -565
rect -642 -599 -274 -565
rect -184 -599 184 -565
rect 274 -599 642 -565
rect 732 -599 1100 -565
<< locali >>
rect -1276 667 -1180 701
rect 1180 667 1276 701
rect -1276 605 -1242 667
rect 1242 605 1276 667
rect -1116 565 -1100 599
rect -732 565 -716 599
rect -658 565 -642 599
rect -274 565 -258 599
rect -200 565 -184 599
rect 184 565 200 599
rect 258 565 274 599
rect 642 565 658 599
rect 716 565 732 599
rect 1100 565 1116 599
rect -1162 506 -1128 522
rect -1162 114 -1128 130
rect -704 506 -670 522
rect -704 114 -670 130
rect -246 506 -212 522
rect -246 114 -212 130
rect 212 506 246 522
rect 212 114 246 130
rect 670 506 704 522
rect 670 114 704 130
rect 1128 506 1162 522
rect 1128 114 1162 130
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -658 37 -642 71
rect -274 37 -258 71
rect -200 37 -184 71
rect 184 37 200 71
rect 258 37 274 71
rect 642 37 658 71
rect 716 37 732 71
rect 1100 37 1116 71
rect -1116 -71 -1100 -37
rect -732 -71 -716 -37
rect -658 -71 -642 -37
rect -274 -71 -258 -37
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect 258 -71 274 -37
rect 642 -71 658 -37
rect 716 -71 732 -37
rect 1100 -71 1116 -37
rect -1162 -130 -1128 -114
rect -1162 -522 -1128 -506
rect -704 -130 -670 -114
rect -704 -522 -670 -506
rect -246 -130 -212 -114
rect -246 -522 -212 -506
rect 212 -130 246 -114
rect 212 -522 246 -506
rect 670 -130 704 -114
rect 670 -522 704 -506
rect 1128 -130 1162 -114
rect 1128 -522 1162 -506
rect -1116 -599 -1100 -565
rect -732 -599 -716 -565
rect -658 -599 -642 -565
rect -274 -599 -258 -565
rect -200 -599 -184 -565
rect 184 -599 200 -565
rect 258 -599 274 -565
rect 642 -599 658 -565
rect 716 -599 732 -565
rect 1100 -599 1116 -565
rect -1276 -667 -1242 -605
rect 1242 -667 1276 -605
rect -1276 -701 -1180 -667
rect 1180 -701 1276 -667
<< viali >>
rect -1100 565 -732 599
rect -642 565 -274 599
rect -184 565 184 599
rect 274 565 642 599
rect 732 565 1100 599
rect -1162 130 -1128 506
rect -704 130 -670 506
rect -246 130 -212 506
rect 212 130 246 506
rect 670 130 704 506
rect 1128 130 1162 506
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect -1100 -71 -732 -37
rect -642 -71 -274 -37
rect -184 -71 184 -37
rect 274 -71 642 -37
rect 732 -71 1100 -37
rect -1162 -506 -1128 -130
rect -704 -506 -670 -130
rect -246 -506 -212 -130
rect 212 -506 246 -130
rect 670 -506 704 -130
rect 1128 -506 1162 -130
rect -1100 -599 -732 -565
rect -642 -599 -274 -565
rect -184 -599 184 -565
rect 274 -599 642 -565
rect 732 -599 1100 -565
<< metal1 >>
rect -1112 599 -720 605
rect -1112 565 -1100 599
rect -732 565 -720 599
rect -1112 559 -720 565
rect -654 599 -262 605
rect -654 565 -642 599
rect -274 565 -262 599
rect -654 559 -262 565
rect -196 599 196 605
rect -196 565 -184 599
rect 184 565 196 599
rect -196 559 196 565
rect 262 599 654 605
rect 262 565 274 599
rect 642 565 654 599
rect 262 559 654 565
rect 720 599 1112 605
rect 720 565 732 599
rect 1100 565 1112 599
rect 720 559 1112 565
rect -1168 506 -1122 518
rect -1168 130 -1162 506
rect -1128 130 -1122 506
rect -1168 118 -1122 130
rect -710 506 -664 518
rect -710 130 -704 506
rect -670 130 -664 506
rect -710 118 -664 130
rect -252 506 -206 518
rect -252 130 -246 506
rect -212 130 -206 506
rect -252 118 -206 130
rect 206 506 252 518
rect 206 130 212 506
rect 246 130 252 506
rect 206 118 252 130
rect 664 506 710 518
rect 664 130 670 506
rect 704 130 710 506
rect 664 118 710 130
rect 1122 506 1168 518
rect 1122 130 1128 506
rect 1162 130 1168 506
rect 1122 118 1168 130
rect -1112 71 -720 77
rect -1112 37 -1100 71
rect -732 37 -720 71
rect -1112 31 -720 37
rect -654 71 -262 77
rect -654 37 -642 71
rect -274 37 -262 71
rect -654 31 -262 37
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect 262 71 654 77
rect 262 37 274 71
rect 642 37 654 71
rect 262 31 654 37
rect 720 71 1112 77
rect 720 37 732 71
rect 1100 37 1112 71
rect 720 31 1112 37
rect -1112 -37 -720 -31
rect -1112 -71 -1100 -37
rect -732 -71 -720 -37
rect -1112 -77 -720 -71
rect -654 -37 -262 -31
rect -654 -71 -642 -37
rect -274 -71 -262 -37
rect -654 -77 -262 -71
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect 262 -37 654 -31
rect 262 -71 274 -37
rect 642 -71 654 -37
rect 262 -77 654 -71
rect 720 -37 1112 -31
rect 720 -71 732 -37
rect 1100 -71 1112 -37
rect 720 -77 1112 -71
rect -1168 -130 -1122 -118
rect -1168 -506 -1162 -130
rect -1128 -506 -1122 -130
rect -1168 -518 -1122 -506
rect -710 -130 -664 -118
rect -710 -506 -704 -130
rect -670 -506 -664 -130
rect -710 -518 -664 -506
rect -252 -130 -206 -118
rect -252 -506 -246 -130
rect -212 -506 -206 -130
rect -252 -518 -206 -506
rect 206 -130 252 -118
rect 206 -506 212 -130
rect 246 -506 252 -130
rect 206 -518 252 -506
rect 664 -130 710 -118
rect 664 -506 670 -130
rect 704 -506 710 -130
rect 664 -518 710 -506
rect 1122 -130 1168 -118
rect 1122 -506 1128 -130
rect 1162 -506 1168 -130
rect 1122 -518 1168 -506
rect -1112 -565 -720 -559
rect -1112 -599 -1100 -565
rect -732 -599 -720 -565
rect -1112 -605 -720 -599
rect -654 -565 -262 -559
rect -654 -599 -642 -565
rect -274 -599 -262 -565
rect -654 -605 -262 -599
rect -196 -565 196 -559
rect -196 -599 -184 -565
rect 184 -599 196 -565
rect -196 -605 196 -599
rect 262 -565 654 -559
rect 262 -599 274 -565
rect 642 -599 654 -565
rect 262 -605 654 -599
rect 720 -565 1112 -559
rect 720 -599 732 -565
rect 1100 -599 1112 -565
rect 720 -605 1112 -599
<< properties >>
string FIXED_BBOX -1259 -684 1259 684
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 2.0 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
