magic
tech sky130A
magscale 1 2
timestamp 1713144909
<< metal3 >>
rect -3798 3610 -1716 4520
rect -1186 3610 894 4520
rect -3798 3310 894 3610
rect -3798 2440 -1716 3310
rect -1186 2440 894 3310
rect -2916 2200 -2618 2440
rect -304 2200 -6 2440
rect -3798 1312 -1716 2200
rect -1186 1312 894 2200
rect -3798 1012 894 1312
rect -3798 120 -1716 1012
rect -1186 120 894 1012
rect -2916 -120 -2618 120
rect -304 -120 -6 120
rect -3798 -988 -1716 -120
rect -1186 -988 894 -120
rect 1426 -988 3506 -120
rect 3990 -988 6070 -116
rect -3798 -1286 6070 -988
rect -3798 -2200 -1716 -1286
rect -1186 -2200 894 -1286
rect 1426 -2200 3506 -1286
rect 3990 -2196 6070 -1286
rect -2916 -2440 -2618 -2200
rect -304 -2440 -6 -2200
rect 2294 -2440 2592 -2200
rect -3798 -3324 -1716 -2440
rect -1186 -3324 894 -2440
rect 1426 -3324 3506 -2440
rect 4874 -2442 5172 -2196
rect 3986 -3324 6066 -2442
rect -3798 -3622 6066 -3324
rect -3798 -4520 -1716 -3622
rect -1186 -4520 894 -3622
rect 1426 -4520 3506 -3622
rect 3986 -4522 6066 -3622
<< mimcap >>
rect -3758 4440 -1758 4480
rect -3758 2520 -3718 4440
rect -1798 2520 -1758 4440
rect -3758 2480 -1758 2520
rect -1146 4440 854 4480
rect -1146 2520 -1106 4440
rect 814 2520 854 4440
rect -1146 2480 854 2520
rect -3758 2120 -1758 2160
rect -3758 200 -3718 2120
rect -1798 200 -1758 2120
rect -3758 160 -1758 200
rect -1146 2120 854 2160
rect -1146 200 -1106 2120
rect 814 200 854 2120
rect -1146 160 854 200
rect -3758 -200 -1758 -160
rect -3758 -2120 -3718 -200
rect -1798 -2120 -1758 -200
rect -3758 -2160 -1758 -2120
rect -1146 -200 854 -160
rect -1146 -2120 -1106 -200
rect 814 -2120 854 -200
rect -1146 -2160 854 -2120
rect 1466 -200 3466 -160
rect 1466 -2120 1506 -200
rect 3426 -2120 3466 -200
rect 1466 -2160 3466 -2120
rect 4030 -196 6030 -156
rect 4030 -2116 4070 -196
rect 5990 -2116 6030 -196
rect 4030 -2156 6030 -2116
rect -3758 -2520 -1758 -2480
rect -3758 -4440 -3718 -2520
rect -1798 -4440 -1758 -2520
rect -3758 -4480 -1758 -4440
rect -1146 -2520 854 -2480
rect -1146 -4440 -1106 -2520
rect 814 -4440 854 -2520
rect -1146 -4480 854 -4440
rect 1466 -2520 3466 -2480
rect 1466 -4440 1506 -2520
rect 3426 -4440 3466 -2520
rect 1466 -4480 3466 -4440
rect 4030 -2516 6030 -2476
rect 4030 -4436 4070 -2516
rect 5990 -4436 6030 -2516
rect 4030 -4476 6030 -4436
<< mimcapcontact >>
rect -3718 2520 -1798 4440
rect -1106 2520 814 4440
rect -3718 200 -1798 2120
rect -1106 200 814 2120
rect -3718 -2120 -1798 -200
rect -1106 -2120 814 -200
rect 1506 -2120 3426 -200
rect 4070 -2116 5990 -196
rect -3718 -4440 -1798 -2520
rect -1106 -4440 814 -2520
rect 1506 -4440 3426 -2520
rect 4070 -4436 5990 -2516
<< metal4 >>
rect -2810 4441 -2706 4534
rect -198 4441 -94 4534
rect -3719 4440 -1797 4441
rect -3719 2520 -3718 4440
rect -1798 3610 -1797 4440
rect -1107 4440 815 4441
rect -1107 3610 -1106 4440
rect -1798 3310 -1106 3610
rect -1798 2520 -1797 3310
rect -3719 2519 -1797 2520
rect -1107 2520 -1106 3310
rect 814 2520 815 4440
rect -1107 2519 815 2520
rect -2916 2121 -2618 2519
rect -304 2121 -6 2519
rect -3719 2120 -1797 2121
rect -3719 200 -3718 2120
rect -1798 1312 -1797 2120
rect -1107 2120 815 2121
rect -1107 1312 -1106 2120
rect -1798 1012 -1106 1312
rect -1798 200 -1797 1012
rect -3719 199 -1797 200
rect -1107 200 -1106 1012
rect 814 200 815 2120
rect -1107 199 815 200
rect -2916 -199 -2618 199
rect -304 -199 -6 199
rect 2414 -199 2518 -114
rect 4978 -195 5082 -102
rect 4069 -196 5991 -195
rect -3719 -200 -1797 -199
rect -3719 -2120 -3718 -200
rect -1798 -988 -1797 -200
rect -1107 -200 815 -199
rect -1107 -988 -1106 -200
rect -1798 -1286 -1106 -988
rect -1798 -2120 -1797 -1286
rect -3719 -2121 -1797 -2120
rect -1107 -2120 -1106 -1286
rect 814 -988 815 -200
rect 1505 -200 3427 -199
rect 1505 -988 1506 -200
rect 814 -1286 1506 -988
rect 814 -2120 815 -1286
rect -1107 -2121 815 -2120
rect 1505 -2120 1506 -1286
rect 3426 -988 3427 -200
rect 4069 -988 4070 -196
rect 3426 -1286 4070 -988
rect 3426 -2120 3427 -1286
rect 4069 -2116 4070 -1286
rect 5990 -2116 5991 -196
rect 4069 -2117 5991 -2116
rect 1505 -2121 3427 -2120
rect -2916 -2519 -2618 -2121
rect -304 -2519 -6 -2121
rect 2294 -2519 2592 -2121
rect 4874 -2515 5172 -2117
rect 4069 -2516 5991 -2515
rect -3719 -2520 -1797 -2519
rect -3719 -4440 -3718 -2520
rect -1798 -3324 -1797 -2520
rect -1107 -2520 815 -2519
rect -1107 -3324 -1106 -2520
rect -1798 -3622 -1106 -3324
rect -1798 -4440 -1797 -3622
rect -3719 -4441 -1797 -4440
rect -1107 -4440 -1106 -3622
rect 814 -3324 815 -2520
rect 1505 -2520 3427 -2519
rect 1505 -3324 1506 -2520
rect 814 -3622 1506 -3324
rect 814 -4440 815 -3622
rect -1107 -4441 815 -4440
rect 1505 -4440 1506 -3622
rect 3426 -3324 3427 -2520
rect 4069 -3324 4070 -2516
rect 3426 -3622 4070 -3324
rect 3426 -4440 3427 -3622
rect 4069 -4436 4070 -3622
rect 5990 -4436 5991 -2516
rect 4069 -4437 5991 -4436
rect 1505 -4441 3427 -4440
rect -2810 -4532 -2706 -4441
rect -198 -4532 -94 -4441
rect 2414 -4532 2518 -4441
rect 4978 -4522 5082 -4437
<< properties >>
string FIXED_BBOX 1426 2440 3506 4520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10 l 10 val 207.6 carea 2.00 cperi 0.19 nx 3 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
