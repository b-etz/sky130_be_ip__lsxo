magic
tech sky130A
magscale 1 2
timestamp 1712250795
<< metal3 >>
rect -10328 4492 -7956 4520
rect -10328 2468 -8040 4492
rect -7976 2468 -7956 4492
rect -10328 2440 -7956 2468
rect -7716 4492 -5344 4520
rect -7716 2468 -5428 4492
rect -5364 2468 -5344 4492
rect -7716 2440 -5344 2468
rect -5104 4492 -2732 4520
rect -5104 2468 -2816 4492
rect -2752 2468 -2732 4492
rect -5104 2440 -2732 2468
rect -2492 4492 -120 4520
rect -2492 2468 -204 4492
rect -140 2468 -120 4492
rect -2492 2440 -120 2468
rect 120 4492 2492 4520
rect 120 2468 2408 4492
rect 2472 2468 2492 4492
rect 120 2440 2492 2468
rect 2732 4492 5104 4520
rect 2732 2468 5020 4492
rect 5084 2468 5104 4492
rect 2732 2440 5104 2468
rect 5344 4492 7716 4520
rect 5344 2468 7632 4492
rect 7696 2468 7716 4492
rect 5344 2440 7716 2468
rect 7956 4492 10328 4520
rect 7956 2468 10244 4492
rect 10308 2468 10328 4492
rect 7956 2440 10328 2468
rect -10328 2172 -7956 2200
rect -10328 148 -8040 2172
rect -7976 148 -7956 2172
rect -10328 120 -7956 148
rect -7716 2172 -5344 2200
rect -7716 148 -5428 2172
rect -5364 148 -5344 2172
rect -7716 120 -5344 148
rect -5104 2172 -2732 2200
rect -5104 148 -2816 2172
rect -2752 148 -2732 2172
rect -5104 120 -2732 148
rect -2492 2172 -120 2200
rect -2492 148 -204 2172
rect -140 148 -120 2172
rect -2492 120 -120 148
rect 120 2172 2492 2200
rect 120 148 2408 2172
rect 2472 148 2492 2172
rect 120 120 2492 148
rect 2732 2172 5104 2200
rect 2732 148 5020 2172
rect 5084 148 5104 2172
rect 2732 120 5104 148
rect 5344 2172 7716 2200
rect 5344 148 7632 2172
rect 7696 148 7716 2172
rect 5344 120 7716 148
rect 7956 2172 10328 2200
rect 7956 148 10244 2172
rect 10308 148 10328 2172
rect 7956 120 10328 148
rect -10328 -148 -7956 -120
rect -10328 -2172 -8040 -148
rect -7976 -2172 -7956 -148
rect -10328 -2200 -7956 -2172
rect -7716 -148 -5344 -120
rect -7716 -2172 -5428 -148
rect -5364 -2172 -5344 -148
rect -7716 -2200 -5344 -2172
rect -5104 -148 -2732 -120
rect -5104 -2172 -2816 -148
rect -2752 -2172 -2732 -148
rect -5104 -2200 -2732 -2172
rect -2492 -148 -120 -120
rect -2492 -2172 -204 -148
rect -140 -2172 -120 -148
rect -2492 -2200 -120 -2172
rect 120 -148 2492 -120
rect 120 -2172 2408 -148
rect 2472 -2172 2492 -148
rect 120 -2200 2492 -2172
rect 2732 -148 5104 -120
rect 2732 -2172 5020 -148
rect 5084 -2172 5104 -148
rect 2732 -2200 5104 -2172
rect 5344 -148 7716 -120
rect 5344 -2172 7632 -148
rect 7696 -2172 7716 -148
rect 5344 -2200 7716 -2172
rect 7956 -148 10328 -120
rect 7956 -2172 10244 -148
rect 10308 -2172 10328 -148
rect 7956 -2200 10328 -2172
rect -10328 -2468 -7956 -2440
rect -10328 -4492 -8040 -2468
rect -7976 -4492 -7956 -2468
rect -10328 -4520 -7956 -4492
rect -7716 -2468 -5344 -2440
rect -7716 -4492 -5428 -2468
rect -5364 -4492 -5344 -2468
rect -7716 -4520 -5344 -4492
rect -5104 -2468 -2732 -2440
rect -5104 -4492 -2816 -2468
rect -2752 -4492 -2732 -2468
rect -5104 -4520 -2732 -4492
rect -2492 -2468 -120 -2440
rect -2492 -4492 -204 -2468
rect -140 -4492 -120 -2468
rect -2492 -4520 -120 -4492
rect 120 -2468 2492 -2440
rect 120 -4492 2408 -2468
rect 2472 -4492 2492 -2468
rect 120 -4520 2492 -4492
rect 2732 -2468 5104 -2440
rect 2732 -4492 5020 -2468
rect 5084 -4492 5104 -2468
rect 2732 -4520 5104 -4492
rect 5344 -2468 7716 -2440
rect 5344 -4492 7632 -2468
rect 7696 -4492 7716 -2468
rect 5344 -4520 7716 -4492
rect 7956 -2468 10328 -2440
rect 7956 -4492 10244 -2468
rect 10308 -4492 10328 -2468
rect 7956 -4520 10328 -4492
<< via3 >>
rect -8040 2468 -7976 4492
rect -5428 2468 -5364 4492
rect -2816 2468 -2752 4492
rect -204 2468 -140 4492
rect 2408 2468 2472 4492
rect 5020 2468 5084 4492
rect 7632 2468 7696 4492
rect 10244 2468 10308 4492
rect -8040 148 -7976 2172
rect -5428 148 -5364 2172
rect -2816 148 -2752 2172
rect -204 148 -140 2172
rect 2408 148 2472 2172
rect 5020 148 5084 2172
rect 7632 148 7696 2172
rect 10244 148 10308 2172
rect -8040 -2172 -7976 -148
rect -5428 -2172 -5364 -148
rect -2816 -2172 -2752 -148
rect -204 -2172 -140 -148
rect 2408 -2172 2472 -148
rect 5020 -2172 5084 -148
rect 7632 -2172 7696 -148
rect 10244 -2172 10308 -148
rect -8040 -4492 -7976 -2468
rect -5428 -4492 -5364 -2468
rect -2816 -4492 -2752 -2468
rect -204 -4492 -140 -2468
rect 2408 -4492 2472 -2468
rect 5020 -4492 5084 -2468
rect 7632 -4492 7696 -2468
rect 10244 -4492 10308 -2468
<< mimcap >>
rect -10288 4440 -8288 4480
rect -10288 2520 -10248 4440
rect -8328 2520 -8288 4440
rect -10288 2480 -8288 2520
rect -7676 4440 -5676 4480
rect -7676 2520 -7636 4440
rect -5716 2520 -5676 4440
rect -7676 2480 -5676 2520
rect -5064 4440 -3064 4480
rect -5064 2520 -5024 4440
rect -3104 2520 -3064 4440
rect -5064 2480 -3064 2520
rect -2452 4440 -452 4480
rect -2452 2520 -2412 4440
rect -492 2520 -452 4440
rect -2452 2480 -452 2520
rect 160 4440 2160 4480
rect 160 2520 200 4440
rect 2120 2520 2160 4440
rect 160 2480 2160 2520
rect 2772 4440 4772 4480
rect 2772 2520 2812 4440
rect 4732 2520 4772 4440
rect 2772 2480 4772 2520
rect 5384 4440 7384 4480
rect 5384 2520 5424 4440
rect 7344 2520 7384 4440
rect 5384 2480 7384 2520
rect 7996 4440 9996 4480
rect 7996 2520 8036 4440
rect 9956 2520 9996 4440
rect 7996 2480 9996 2520
rect -10288 2120 -8288 2160
rect -10288 200 -10248 2120
rect -8328 200 -8288 2120
rect -10288 160 -8288 200
rect -7676 2120 -5676 2160
rect -7676 200 -7636 2120
rect -5716 200 -5676 2120
rect -7676 160 -5676 200
rect -5064 2120 -3064 2160
rect -5064 200 -5024 2120
rect -3104 200 -3064 2120
rect -5064 160 -3064 200
rect -2452 2120 -452 2160
rect -2452 200 -2412 2120
rect -492 200 -452 2120
rect -2452 160 -452 200
rect 160 2120 2160 2160
rect 160 200 200 2120
rect 2120 200 2160 2120
rect 160 160 2160 200
rect 2772 2120 4772 2160
rect 2772 200 2812 2120
rect 4732 200 4772 2120
rect 2772 160 4772 200
rect 5384 2120 7384 2160
rect 5384 200 5424 2120
rect 7344 200 7384 2120
rect 5384 160 7384 200
rect 7996 2120 9996 2160
rect 7996 200 8036 2120
rect 9956 200 9996 2120
rect 7996 160 9996 200
rect -10288 -200 -8288 -160
rect -10288 -2120 -10248 -200
rect -8328 -2120 -8288 -200
rect -10288 -2160 -8288 -2120
rect -7676 -200 -5676 -160
rect -7676 -2120 -7636 -200
rect -5716 -2120 -5676 -200
rect -7676 -2160 -5676 -2120
rect -5064 -200 -3064 -160
rect -5064 -2120 -5024 -200
rect -3104 -2120 -3064 -200
rect -5064 -2160 -3064 -2120
rect -2452 -200 -452 -160
rect -2452 -2120 -2412 -200
rect -492 -2120 -452 -200
rect -2452 -2160 -452 -2120
rect 160 -200 2160 -160
rect 160 -2120 200 -200
rect 2120 -2120 2160 -200
rect 160 -2160 2160 -2120
rect 2772 -200 4772 -160
rect 2772 -2120 2812 -200
rect 4732 -2120 4772 -200
rect 2772 -2160 4772 -2120
rect 5384 -200 7384 -160
rect 5384 -2120 5424 -200
rect 7344 -2120 7384 -200
rect 5384 -2160 7384 -2120
rect 7996 -200 9996 -160
rect 7996 -2120 8036 -200
rect 9956 -2120 9996 -200
rect 7996 -2160 9996 -2120
rect -10288 -2520 -8288 -2480
rect -10288 -4440 -10248 -2520
rect -8328 -4440 -8288 -2520
rect -10288 -4480 -8288 -4440
rect -7676 -2520 -5676 -2480
rect -7676 -4440 -7636 -2520
rect -5716 -4440 -5676 -2520
rect -7676 -4480 -5676 -4440
rect -5064 -2520 -3064 -2480
rect -5064 -4440 -5024 -2520
rect -3104 -4440 -3064 -2520
rect -5064 -4480 -3064 -4440
rect -2452 -2520 -452 -2480
rect -2452 -4440 -2412 -2520
rect -492 -4440 -452 -2520
rect -2452 -4480 -452 -4440
rect 160 -2520 2160 -2480
rect 160 -4440 200 -2520
rect 2120 -4440 2160 -2520
rect 160 -4480 2160 -4440
rect 2772 -2520 4772 -2480
rect 2772 -4440 2812 -2520
rect 4732 -4440 4772 -2520
rect 2772 -4480 4772 -4440
rect 5384 -2520 7384 -2480
rect 5384 -4440 5424 -2520
rect 7344 -4440 7384 -2520
rect 5384 -4480 7384 -4440
rect 7996 -2520 9996 -2480
rect 7996 -4440 8036 -2520
rect 9956 -4440 9996 -2520
rect 7996 -4480 9996 -4440
<< mimcapcontact >>
rect -10248 2520 -8328 4440
rect -7636 2520 -5716 4440
rect -5024 2520 -3104 4440
rect -2412 2520 -492 4440
rect 200 2520 2120 4440
rect 2812 2520 4732 4440
rect 5424 2520 7344 4440
rect 8036 2520 9956 4440
rect -10248 200 -8328 2120
rect -7636 200 -5716 2120
rect -5024 200 -3104 2120
rect -2412 200 -492 2120
rect 200 200 2120 2120
rect 2812 200 4732 2120
rect 5424 200 7344 2120
rect 8036 200 9956 2120
rect -10248 -2120 -8328 -200
rect -7636 -2120 -5716 -200
rect -5024 -2120 -3104 -200
rect -2412 -2120 -492 -200
rect 200 -2120 2120 -200
rect 2812 -2120 4732 -200
rect 5424 -2120 7344 -200
rect 8036 -2120 9956 -200
rect -10248 -4440 -8328 -2520
rect -7636 -4440 -5716 -2520
rect -5024 -4440 -3104 -2520
rect -2412 -4440 -492 -2520
rect 200 -4440 2120 -2520
rect 2812 -4440 4732 -2520
rect 5424 -4440 7344 -2520
rect 8036 -4440 9956 -2520
<< metal4 >>
rect -9340 4441 -9236 4640
rect -8060 4492 -7956 4640
rect -10249 4440 -8327 4441
rect -10249 2520 -10248 4440
rect -8328 2520 -8327 4440
rect -10249 2519 -8327 2520
rect -9340 2121 -9236 2519
rect -8060 2468 -8040 4492
rect -7976 2468 -7956 4492
rect -6728 4441 -6624 4640
rect -5448 4492 -5344 4640
rect -7637 4440 -5715 4441
rect -7637 2520 -7636 4440
rect -5716 2520 -5715 4440
rect -7637 2519 -5715 2520
rect -8060 2172 -7956 2468
rect -10249 2120 -8327 2121
rect -10249 200 -10248 2120
rect -8328 200 -8327 2120
rect -10249 199 -8327 200
rect -9340 -199 -9236 199
rect -8060 148 -8040 2172
rect -7976 148 -7956 2172
rect -6728 2121 -6624 2519
rect -5448 2468 -5428 4492
rect -5364 2468 -5344 4492
rect -4116 4441 -4012 4640
rect -2836 4492 -2732 4640
rect -5025 4440 -3103 4441
rect -5025 2520 -5024 4440
rect -3104 2520 -3103 4440
rect -5025 2519 -3103 2520
rect -5448 2172 -5344 2468
rect -7637 2120 -5715 2121
rect -7637 200 -7636 2120
rect -5716 200 -5715 2120
rect -7637 199 -5715 200
rect -8060 -148 -7956 148
rect -10249 -200 -8327 -199
rect -10249 -2120 -10248 -200
rect -8328 -2120 -8327 -200
rect -10249 -2121 -8327 -2120
rect -9340 -2519 -9236 -2121
rect -8060 -2172 -8040 -148
rect -7976 -2172 -7956 -148
rect -6728 -199 -6624 199
rect -5448 148 -5428 2172
rect -5364 148 -5344 2172
rect -4116 2121 -4012 2519
rect -2836 2468 -2816 4492
rect -2752 2468 -2732 4492
rect -1504 4441 -1400 4640
rect -224 4492 -120 4640
rect -2413 4440 -491 4441
rect -2413 2520 -2412 4440
rect -492 2520 -491 4440
rect -2413 2519 -491 2520
rect -2836 2172 -2732 2468
rect -5025 2120 -3103 2121
rect -5025 200 -5024 2120
rect -3104 200 -3103 2120
rect -5025 199 -3103 200
rect -5448 -148 -5344 148
rect -7637 -200 -5715 -199
rect -7637 -2120 -7636 -200
rect -5716 -2120 -5715 -200
rect -7637 -2121 -5715 -2120
rect -8060 -2468 -7956 -2172
rect -10249 -2520 -8327 -2519
rect -10249 -4440 -10248 -2520
rect -8328 -4440 -8327 -2520
rect -10249 -4441 -8327 -4440
rect -9340 -4640 -9236 -4441
rect -8060 -4492 -8040 -2468
rect -7976 -4492 -7956 -2468
rect -6728 -2519 -6624 -2121
rect -5448 -2172 -5428 -148
rect -5364 -2172 -5344 -148
rect -4116 -199 -4012 199
rect -2836 148 -2816 2172
rect -2752 148 -2732 2172
rect -1504 2121 -1400 2519
rect -224 2468 -204 4492
rect -140 2468 -120 4492
rect 1108 4441 1212 4640
rect 2388 4492 2492 4640
rect 199 4440 2121 4441
rect 199 2520 200 4440
rect 2120 2520 2121 4440
rect 199 2519 2121 2520
rect -224 2172 -120 2468
rect -2413 2120 -491 2121
rect -2413 200 -2412 2120
rect -492 200 -491 2120
rect -2413 199 -491 200
rect -2836 -148 -2732 148
rect -5025 -200 -3103 -199
rect -5025 -2120 -5024 -200
rect -3104 -2120 -3103 -200
rect -5025 -2121 -3103 -2120
rect -5448 -2468 -5344 -2172
rect -7637 -2520 -5715 -2519
rect -7637 -4440 -7636 -2520
rect -5716 -4440 -5715 -2520
rect -7637 -4441 -5715 -4440
rect -8060 -4640 -7956 -4492
rect -6728 -4640 -6624 -4441
rect -5448 -4492 -5428 -2468
rect -5364 -4492 -5344 -2468
rect -4116 -2519 -4012 -2121
rect -2836 -2172 -2816 -148
rect -2752 -2172 -2732 -148
rect -1504 -199 -1400 199
rect -224 148 -204 2172
rect -140 148 -120 2172
rect 1108 2121 1212 2519
rect 2388 2468 2408 4492
rect 2472 2468 2492 4492
rect 3720 4441 3824 4640
rect 5000 4492 5104 4640
rect 2811 4440 4733 4441
rect 2811 2520 2812 4440
rect 4732 2520 4733 4440
rect 2811 2519 4733 2520
rect 2388 2172 2492 2468
rect 199 2120 2121 2121
rect 199 200 200 2120
rect 2120 200 2121 2120
rect 199 199 2121 200
rect -224 -148 -120 148
rect -2413 -200 -491 -199
rect -2413 -2120 -2412 -200
rect -492 -2120 -491 -200
rect -2413 -2121 -491 -2120
rect -2836 -2468 -2732 -2172
rect -5025 -2520 -3103 -2519
rect -5025 -4440 -5024 -2520
rect -3104 -4440 -3103 -2520
rect -5025 -4441 -3103 -4440
rect -5448 -4640 -5344 -4492
rect -4116 -4640 -4012 -4441
rect -2836 -4492 -2816 -2468
rect -2752 -4492 -2732 -2468
rect -1504 -2519 -1400 -2121
rect -224 -2172 -204 -148
rect -140 -2172 -120 -148
rect 1108 -199 1212 199
rect 2388 148 2408 2172
rect 2472 148 2492 2172
rect 3720 2121 3824 2519
rect 5000 2468 5020 4492
rect 5084 2468 5104 4492
rect 6332 4441 6436 4640
rect 7612 4492 7716 4640
rect 5423 4440 7345 4441
rect 5423 2520 5424 4440
rect 7344 2520 7345 4440
rect 5423 2519 7345 2520
rect 5000 2172 5104 2468
rect 2811 2120 4733 2121
rect 2811 200 2812 2120
rect 4732 200 4733 2120
rect 2811 199 4733 200
rect 2388 -148 2492 148
rect 199 -200 2121 -199
rect 199 -2120 200 -200
rect 2120 -2120 2121 -200
rect 199 -2121 2121 -2120
rect -224 -2468 -120 -2172
rect -2413 -2520 -491 -2519
rect -2413 -4440 -2412 -2520
rect -492 -4440 -491 -2520
rect -2413 -4441 -491 -4440
rect -2836 -4640 -2732 -4492
rect -1504 -4640 -1400 -4441
rect -224 -4492 -204 -2468
rect -140 -4492 -120 -2468
rect 1108 -2519 1212 -2121
rect 2388 -2172 2408 -148
rect 2472 -2172 2492 -148
rect 3720 -199 3824 199
rect 5000 148 5020 2172
rect 5084 148 5104 2172
rect 6332 2121 6436 2519
rect 7612 2468 7632 4492
rect 7696 2468 7716 4492
rect 8944 4441 9048 4640
rect 10224 4492 10328 4640
rect 8035 4440 9957 4441
rect 8035 2520 8036 4440
rect 9956 2520 9957 4440
rect 8035 2519 9957 2520
rect 7612 2172 7716 2468
rect 5423 2120 7345 2121
rect 5423 200 5424 2120
rect 7344 200 7345 2120
rect 5423 199 7345 200
rect 5000 -148 5104 148
rect 2811 -200 4733 -199
rect 2811 -2120 2812 -200
rect 4732 -2120 4733 -200
rect 2811 -2121 4733 -2120
rect 2388 -2468 2492 -2172
rect 199 -2520 2121 -2519
rect 199 -4440 200 -2520
rect 2120 -4440 2121 -2520
rect 199 -4441 2121 -4440
rect -224 -4640 -120 -4492
rect 1108 -4640 1212 -4441
rect 2388 -4492 2408 -2468
rect 2472 -4492 2492 -2468
rect 3720 -2519 3824 -2121
rect 5000 -2172 5020 -148
rect 5084 -2172 5104 -148
rect 6332 -199 6436 199
rect 7612 148 7632 2172
rect 7696 148 7716 2172
rect 8944 2121 9048 2519
rect 10224 2468 10244 4492
rect 10308 2468 10328 4492
rect 10224 2172 10328 2468
rect 8035 2120 9957 2121
rect 8035 200 8036 2120
rect 9956 200 9957 2120
rect 8035 199 9957 200
rect 7612 -148 7716 148
rect 5423 -200 7345 -199
rect 5423 -2120 5424 -200
rect 7344 -2120 7345 -200
rect 5423 -2121 7345 -2120
rect 5000 -2468 5104 -2172
rect 2811 -2520 4733 -2519
rect 2811 -4440 2812 -2520
rect 4732 -4440 4733 -2520
rect 2811 -4441 4733 -4440
rect 2388 -4640 2492 -4492
rect 3720 -4640 3824 -4441
rect 5000 -4492 5020 -2468
rect 5084 -4492 5104 -2468
rect 6332 -2519 6436 -2121
rect 7612 -2172 7632 -148
rect 7696 -2172 7716 -148
rect 8944 -199 9048 199
rect 10224 148 10244 2172
rect 10308 148 10328 2172
rect 10224 -148 10328 148
rect 8035 -200 9957 -199
rect 8035 -2120 8036 -200
rect 9956 -2120 9957 -200
rect 8035 -2121 9957 -2120
rect 7612 -2468 7716 -2172
rect 5423 -2520 7345 -2519
rect 5423 -4440 5424 -2520
rect 7344 -4440 7345 -2520
rect 5423 -4441 7345 -4440
rect 5000 -4640 5104 -4492
rect 6332 -4640 6436 -4441
rect 7612 -4492 7632 -2468
rect 7696 -4492 7716 -2468
rect 8944 -2519 9048 -2121
rect 10224 -2172 10244 -148
rect 10308 -2172 10328 -148
rect 10224 -2468 10328 -2172
rect 8035 -2520 9957 -2519
rect 8035 -4440 8036 -2520
rect 9956 -4440 9957 -2520
rect 8035 -4441 9957 -4440
rect 7612 -4640 7716 -4492
rect 8944 -4640 9048 -4441
rect 10224 -4492 10244 -2468
rect 10308 -4492 10328 -2468
rect 10224 -4640 10328 -4492
<< properties >>
string FIXED_BBOX 7956 2440 10036 4520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 8 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
