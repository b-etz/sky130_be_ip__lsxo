magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< nwell >>
rect -246 -5281 246 5281
<< pmos >>
rect -50 4262 50 5062
rect -50 3226 50 4026
rect -50 2190 50 2990
rect -50 1154 50 1954
rect -50 118 50 918
rect -50 -918 50 -118
rect -50 -1954 50 -1154
rect -50 -2990 50 -2190
rect -50 -4026 50 -3226
rect -50 -5062 50 -4262
<< pdiff >>
rect -108 5050 -50 5062
rect -108 4274 -96 5050
rect -62 4274 -50 5050
rect -108 4262 -50 4274
rect 50 5050 108 5062
rect 50 4274 62 5050
rect 96 4274 108 5050
rect 50 4262 108 4274
rect -108 4014 -50 4026
rect -108 3238 -96 4014
rect -62 3238 -50 4014
rect -108 3226 -50 3238
rect 50 4014 108 4026
rect 50 3238 62 4014
rect 96 3238 108 4014
rect 50 3226 108 3238
rect -108 2978 -50 2990
rect -108 2202 -96 2978
rect -62 2202 -50 2978
rect -108 2190 -50 2202
rect 50 2978 108 2990
rect 50 2202 62 2978
rect 96 2202 108 2978
rect 50 2190 108 2202
rect -108 1942 -50 1954
rect -108 1166 -96 1942
rect -62 1166 -50 1942
rect -108 1154 -50 1166
rect 50 1942 108 1954
rect 50 1166 62 1942
rect 96 1166 108 1942
rect 50 1154 108 1166
rect -108 906 -50 918
rect -108 130 -96 906
rect -62 130 -50 906
rect -108 118 -50 130
rect 50 906 108 918
rect 50 130 62 906
rect 96 130 108 906
rect 50 118 108 130
rect -108 -130 -50 -118
rect -108 -906 -96 -130
rect -62 -906 -50 -130
rect -108 -918 -50 -906
rect 50 -130 108 -118
rect 50 -906 62 -130
rect 96 -906 108 -130
rect 50 -918 108 -906
rect -108 -1166 -50 -1154
rect -108 -1942 -96 -1166
rect -62 -1942 -50 -1166
rect -108 -1954 -50 -1942
rect 50 -1166 108 -1154
rect 50 -1942 62 -1166
rect 96 -1942 108 -1166
rect 50 -1954 108 -1942
rect -108 -2202 -50 -2190
rect -108 -2978 -96 -2202
rect -62 -2978 -50 -2202
rect -108 -2990 -50 -2978
rect 50 -2202 108 -2190
rect 50 -2978 62 -2202
rect 96 -2978 108 -2202
rect 50 -2990 108 -2978
rect -108 -3238 -50 -3226
rect -108 -4014 -96 -3238
rect -62 -4014 -50 -3238
rect -108 -4026 -50 -4014
rect 50 -3238 108 -3226
rect 50 -4014 62 -3238
rect 96 -4014 108 -3238
rect 50 -4026 108 -4014
rect -108 -4274 -50 -4262
rect -108 -5050 -96 -4274
rect -62 -5050 -50 -4274
rect -108 -5062 -50 -5050
rect 50 -4274 108 -4262
rect 50 -5050 62 -4274
rect 96 -5050 108 -4274
rect 50 -5062 108 -5050
<< pdiffc >>
rect -96 4274 -62 5050
rect 62 4274 96 5050
rect -96 3238 -62 4014
rect 62 3238 96 4014
rect -96 2202 -62 2978
rect 62 2202 96 2978
rect -96 1166 -62 1942
rect 62 1166 96 1942
rect -96 130 -62 906
rect 62 130 96 906
rect -96 -906 -62 -130
rect 62 -906 96 -130
rect -96 -1942 -62 -1166
rect 62 -1942 96 -1166
rect -96 -2978 -62 -2202
rect 62 -2978 96 -2202
rect -96 -4014 -62 -3238
rect 62 -4014 96 -3238
rect -96 -5050 -62 -4274
rect 62 -5050 96 -4274
<< nsubdiff >>
rect -210 5211 -114 5245
rect 114 5211 210 5245
rect -210 5149 -176 5211
rect 176 5149 210 5211
rect -210 -5211 -176 -5149
rect 176 -5211 210 -5149
rect -210 -5245 -114 -5211
rect 114 -5245 210 -5211
<< nsubdiffcont >>
rect -114 5211 114 5245
rect -210 -5149 -176 5149
rect 176 -5149 210 5149
rect -114 -5245 114 -5211
<< poly >>
rect -50 5143 50 5159
rect -50 5109 -34 5143
rect 34 5109 50 5143
rect -50 5062 50 5109
rect -50 4215 50 4262
rect -50 4181 -34 4215
rect 34 4181 50 4215
rect -50 4165 50 4181
rect -50 4107 50 4123
rect -50 4073 -34 4107
rect 34 4073 50 4107
rect -50 4026 50 4073
rect -50 3179 50 3226
rect -50 3145 -34 3179
rect 34 3145 50 3179
rect -50 3129 50 3145
rect -50 3071 50 3087
rect -50 3037 -34 3071
rect 34 3037 50 3071
rect -50 2990 50 3037
rect -50 2143 50 2190
rect -50 2109 -34 2143
rect 34 2109 50 2143
rect -50 2093 50 2109
rect -50 2035 50 2051
rect -50 2001 -34 2035
rect 34 2001 50 2035
rect -50 1954 50 2001
rect -50 1107 50 1154
rect -50 1073 -34 1107
rect 34 1073 50 1107
rect -50 1057 50 1073
rect -50 999 50 1015
rect -50 965 -34 999
rect 34 965 50 999
rect -50 918 50 965
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect -50 -965 50 -918
rect -50 -999 -34 -965
rect 34 -999 50 -965
rect -50 -1015 50 -999
rect -50 -1073 50 -1057
rect -50 -1107 -34 -1073
rect 34 -1107 50 -1073
rect -50 -1154 50 -1107
rect -50 -2001 50 -1954
rect -50 -2035 -34 -2001
rect 34 -2035 50 -2001
rect -50 -2051 50 -2035
rect -50 -2109 50 -2093
rect -50 -2143 -34 -2109
rect 34 -2143 50 -2109
rect -50 -2190 50 -2143
rect -50 -3037 50 -2990
rect -50 -3071 -34 -3037
rect 34 -3071 50 -3037
rect -50 -3087 50 -3071
rect -50 -3145 50 -3129
rect -50 -3179 -34 -3145
rect 34 -3179 50 -3145
rect -50 -3226 50 -3179
rect -50 -4073 50 -4026
rect -50 -4107 -34 -4073
rect 34 -4107 50 -4073
rect -50 -4123 50 -4107
rect -50 -4181 50 -4165
rect -50 -4215 -34 -4181
rect 34 -4215 50 -4181
rect -50 -4262 50 -4215
rect -50 -5109 50 -5062
rect -50 -5143 -34 -5109
rect 34 -5143 50 -5109
rect -50 -5159 50 -5143
<< polycont >>
rect -34 5109 34 5143
rect -34 4181 34 4215
rect -34 4073 34 4107
rect -34 3145 34 3179
rect -34 3037 34 3071
rect -34 2109 34 2143
rect -34 2001 34 2035
rect -34 1073 34 1107
rect -34 965 34 999
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -999 34 -965
rect -34 -1107 34 -1073
rect -34 -2035 34 -2001
rect -34 -2143 34 -2109
rect -34 -3071 34 -3037
rect -34 -3179 34 -3145
rect -34 -4107 34 -4073
rect -34 -4215 34 -4181
rect -34 -5143 34 -5109
<< locali >>
rect -210 5211 -114 5245
rect 114 5211 210 5245
rect -210 5149 -176 5211
rect 176 5149 210 5211
rect -50 5109 -34 5143
rect 34 5109 50 5143
rect -96 5050 -62 5066
rect -96 4258 -62 4274
rect 62 5050 96 5066
rect 62 4258 96 4274
rect -50 4181 -34 4215
rect 34 4181 50 4215
rect -50 4073 -34 4107
rect 34 4073 50 4107
rect -96 4014 -62 4030
rect -96 3222 -62 3238
rect 62 4014 96 4030
rect 62 3222 96 3238
rect -50 3145 -34 3179
rect 34 3145 50 3179
rect -50 3037 -34 3071
rect 34 3037 50 3071
rect -96 2978 -62 2994
rect -96 2186 -62 2202
rect 62 2978 96 2994
rect 62 2186 96 2202
rect -50 2109 -34 2143
rect 34 2109 50 2143
rect -50 2001 -34 2035
rect 34 2001 50 2035
rect -96 1942 -62 1958
rect -96 1150 -62 1166
rect 62 1942 96 1958
rect 62 1150 96 1166
rect -50 1073 -34 1107
rect 34 1073 50 1107
rect -50 965 -34 999
rect 34 965 50 999
rect -96 906 -62 922
rect -96 114 -62 130
rect 62 906 96 922
rect 62 114 96 130
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -130 -62 -114
rect -96 -922 -62 -906
rect 62 -130 96 -114
rect 62 -922 96 -906
rect -50 -999 -34 -965
rect 34 -999 50 -965
rect -50 -1107 -34 -1073
rect 34 -1107 50 -1073
rect -96 -1166 -62 -1150
rect -96 -1958 -62 -1942
rect 62 -1166 96 -1150
rect 62 -1958 96 -1942
rect -50 -2035 -34 -2001
rect 34 -2035 50 -2001
rect -50 -2143 -34 -2109
rect 34 -2143 50 -2109
rect -96 -2202 -62 -2186
rect -96 -2994 -62 -2978
rect 62 -2202 96 -2186
rect 62 -2994 96 -2978
rect -50 -3071 -34 -3037
rect 34 -3071 50 -3037
rect -50 -3179 -34 -3145
rect 34 -3179 50 -3145
rect -96 -3238 -62 -3222
rect -96 -4030 -62 -4014
rect 62 -3238 96 -3222
rect 62 -4030 96 -4014
rect -50 -4107 -34 -4073
rect 34 -4107 50 -4073
rect -50 -4215 -34 -4181
rect 34 -4215 50 -4181
rect -96 -4274 -62 -4258
rect -96 -5066 -62 -5050
rect 62 -4274 96 -4258
rect 62 -5066 96 -5050
rect -50 -5143 -34 -5109
rect 34 -5143 50 -5109
rect -210 -5211 -176 -5149
rect 176 -5211 210 -5149
rect -210 -5245 -114 -5211
rect 114 -5245 210 -5211
<< viali >>
rect -34 5109 34 5143
rect -96 4274 -62 5050
rect 62 4274 96 5050
rect -34 4181 34 4215
rect -34 4073 34 4107
rect -96 3238 -62 4014
rect 62 3238 96 4014
rect -34 3145 34 3179
rect -34 3037 34 3071
rect -96 2202 -62 2978
rect 62 2202 96 2978
rect -34 2109 34 2143
rect -34 2001 34 2035
rect -96 1166 -62 1942
rect 62 1166 96 1942
rect -34 1073 34 1107
rect -34 965 34 999
rect -96 130 -62 906
rect 62 130 96 906
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -906 -62 -130
rect 62 -906 96 -130
rect -34 -999 34 -965
rect -34 -1107 34 -1073
rect -96 -1942 -62 -1166
rect 62 -1942 96 -1166
rect -34 -2035 34 -2001
rect -34 -2143 34 -2109
rect -96 -2978 -62 -2202
rect 62 -2978 96 -2202
rect -34 -3071 34 -3037
rect -34 -3179 34 -3145
rect -96 -4014 -62 -3238
rect 62 -4014 96 -3238
rect -34 -4107 34 -4073
rect -34 -4215 34 -4181
rect -96 -5050 -62 -4274
rect 62 -5050 96 -4274
rect -34 -5143 34 -5109
<< metal1 >>
rect -46 5143 46 5149
rect -46 5109 -34 5143
rect 34 5109 46 5143
rect -46 5103 46 5109
rect -102 5050 -56 5062
rect -102 4274 -96 5050
rect -62 4274 -56 5050
rect -102 4262 -56 4274
rect 56 5050 102 5062
rect 56 4274 62 5050
rect 96 4274 102 5050
rect 56 4262 102 4274
rect -46 4215 46 4221
rect -46 4181 -34 4215
rect 34 4181 46 4215
rect -46 4175 46 4181
rect -46 4107 46 4113
rect -46 4073 -34 4107
rect 34 4073 46 4107
rect -46 4067 46 4073
rect -102 4014 -56 4026
rect -102 3238 -96 4014
rect -62 3238 -56 4014
rect -102 3226 -56 3238
rect 56 4014 102 4026
rect 56 3238 62 4014
rect 96 3238 102 4014
rect 56 3226 102 3238
rect -46 3179 46 3185
rect -46 3145 -34 3179
rect 34 3145 46 3179
rect -46 3139 46 3145
rect -46 3071 46 3077
rect -46 3037 -34 3071
rect 34 3037 46 3071
rect -46 3031 46 3037
rect -102 2978 -56 2990
rect -102 2202 -96 2978
rect -62 2202 -56 2978
rect -102 2190 -56 2202
rect 56 2978 102 2990
rect 56 2202 62 2978
rect 96 2202 102 2978
rect 56 2190 102 2202
rect -46 2143 46 2149
rect -46 2109 -34 2143
rect 34 2109 46 2143
rect -46 2103 46 2109
rect -46 2035 46 2041
rect -46 2001 -34 2035
rect 34 2001 46 2035
rect -46 1995 46 2001
rect -102 1942 -56 1954
rect -102 1166 -96 1942
rect -62 1166 -56 1942
rect -102 1154 -56 1166
rect 56 1942 102 1954
rect 56 1166 62 1942
rect 96 1166 102 1942
rect 56 1154 102 1166
rect -46 1107 46 1113
rect -46 1073 -34 1107
rect 34 1073 46 1107
rect -46 1067 46 1073
rect -46 999 46 1005
rect -46 965 -34 999
rect 34 965 46 999
rect -46 959 46 965
rect -102 906 -56 918
rect -102 130 -96 906
rect -62 130 -56 906
rect -102 118 -56 130
rect 56 906 102 918
rect 56 130 62 906
rect 96 130 102 906
rect 56 118 102 130
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -130 -56 -118
rect -102 -906 -96 -130
rect -62 -906 -56 -130
rect -102 -918 -56 -906
rect 56 -130 102 -118
rect 56 -906 62 -130
rect 96 -906 102 -130
rect 56 -918 102 -906
rect -46 -965 46 -959
rect -46 -999 -34 -965
rect 34 -999 46 -965
rect -46 -1005 46 -999
rect -46 -1073 46 -1067
rect -46 -1107 -34 -1073
rect 34 -1107 46 -1073
rect -46 -1113 46 -1107
rect -102 -1166 -56 -1154
rect -102 -1942 -96 -1166
rect -62 -1942 -56 -1166
rect -102 -1954 -56 -1942
rect 56 -1166 102 -1154
rect 56 -1942 62 -1166
rect 96 -1942 102 -1166
rect 56 -1954 102 -1942
rect -46 -2001 46 -1995
rect -46 -2035 -34 -2001
rect 34 -2035 46 -2001
rect -46 -2041 46 -2035
rect -46 -2109 46 -2103
rect -46 -2143 -34 -2109
rect 34 -2143 46 -2109
rect -46 -2149 46 -2143
rect -102 -2202 -56 -2190
rect -102 -2978 -96 -2202
rect -62 -2978 -56 -2202
rect -102 -2990 -56 -2978
rect 56 -2202 102 -2190
rect 56 -2978 62 -2202
rect 96 -2978 102 -2202
rect 56 -2990 102 -2978
rect -46 -3037 46 -3031
rect -46 -3071 -34 -3037
rect 34 -3071 46 -3037
rect -46 -3077 46 -3071
rect -46 -3145 46 -3139
rect -46 -3179 -34 -3145
rect 34 -3179 46 -3145
rect -46 -3185 46 -3179
rect -102 -3238 -56 -3226
rect -102 -4014 -96 -3238
rect -62 -4014 -56 -3238
rect -102 -4026 -56 -4014
rect 56 -3238 102 -3226
rect 56 -4014 62 -3238
rect 96 -4014 102 -3238
rect 56 -4026 102 -4014
rect -46 -4073 46 -4067
rect -46 -4107 -34 -4073
rect 34 -4107 46 -4073
rect -46 -4113 46 -4107
rect -46 -4181 46 -4175
rect -46 -4215 -34 -4181
rect 34 -4215 46 -4181
rect -46 -4221 46 -4215
rect -102 -4274 -56 -4262
rect -102 -5050 -96 -4274
rect -62 -5050 -56 -4274
rect -102 -5062 -56 -5050
rect 56 -4274 102 -4262
rect 56 -5050 62 -4274
rect 96 -5050 102 -4274
rect 56 -5062 102 -5050
rect -46 -5109 46 -5103
rect -46 -5143 -34 -5109
rect 34 -5143 46 -5109
rect -46 -5149 46 -5143
<< properties >>
string FIXED_BBOX -193 -5228 193 5228
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.0 l 0.5 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
