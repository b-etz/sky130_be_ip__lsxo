magic
tech sky130A
magscale 1 2
timestamp 1712437813
<< pwell >>
rect -2193 -11102 2193 11102
<< psubdiff >>
rect -2157 11032 -2061 11066
rect 2061 11032 2157 11066
rect -2157 10970 -2123 11032
rect 2123 10970 2157 11032
rect -2157 -11032 -2123 -10970
rect 2123 -11032 2157 -10970
rect -2157 -11066 -2061 -11032
rect 2061 -11066 2157 -11032
<< psubdiffcont >>
rect -2061 11032 2061 11066
rect -2157 -10970 -2123 10970
rect 2123 -10970 2157 10970
rect -2061 -11066 2061 -11032
<< xpolycontact >>
rect 1957 10504 2027 10936
rect -2027 -10936 -1957 -10504
<< xpolyres >>
rect -2027 10330 -1791 10400
rect -2027 -10504 -1957 10330
rect -1861 -10330 -1791 10330
rect -1695 10330 -1459 10400
rect -1695 -10330 -1625 10330
rect -1861 -10400 -1625 -10330
rect -1529 -10330 -1459 10330
rect -1363 10330 -1127 10400
rect -1363 -10330 -1293 10330
rect -1529 -10400 -1293 -10330
rect -1197 -10330 -1127 10330
rect -1031 10330 -795 10400
rect -1031 -10330 -961 10330
rect -1197 -10400 -961 -10330
rect -865 -10330 -795 10330
rect -699 10330 -463 10400
rect -699 -10330 -629 10330
rect -865 -10400 -629 -10330
rect -533 -10330 -463 10330
rect -367 10330 -131 10400
rect -367 -10330 -297 10330
rect -533 -10400 -297 -10330
rect -201 -10330 -131 10330
rect -35 10330 201 10400
rect -35 -10330 35 10330
rect -201 -10400 35 -10330
rect 131 -10330 201 10330
rect 297 10330 533 10400
rect 297 -10330 367 10330
rect 131 -10400 367 -10330
rect 463 -10330 533 10330
rect 629 10330 865 10400
rect 629 -10330 699 10330
rect 463 -10400 699 -10330
rect 795 -10330 865 10330
rect 961 10330 1197 10400
rect 961 -10330 1031 10330
rect 795 -10400 1031 -10330
rect 1127 -10330 1197 10330
rect 1293 10330 1529 10400
rect 1293 -10330 1363 10330
rect 1127 -10400 1363 -10330
rect 1459 -10330 1529 10330
rect 1625 10330 1861 10400
rect 1625 -10330 1695 10330
rect 1459 -10400 1695 -10330
rect 1791 -10330 1861 10330
rect 1957 -10330 2027 10504
rect 1791 -10400 2027 -10330
<< locali >>
rect -2157 11032 -2061 11066
rect 2061 11032 2157 11066
rect -2157 10970 -2123 11032
rect 2123 10970 2157 11032
rect -2157 -11032 -2123 -10970
rect 2123 -11032 2157 -10970
rect -2157 -11066 -2061 -11032
rect 2061 -11066 2157 -11032
<< properties >>
string FIXED_BBOX -2140 -11049 2140 11049
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 104.0 m 1 nx 25 wmin 0.350 lmin 0.50 rho 2000 val 14.906meg dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
