magic
tech sky130A
magscale 1 2
timestamp 1713225924
<< metal3 >>
rect -1892 120 -394 1600
rect -150 130 1336 1610
rect -1892 -1600 -394 -120
rect -150 -1590 1336 -110
<< mimcap >>
rect -1852 1520 -452 1560
rect -1852 200 -1812 1520
rect -492 200 -452 1520
rect -1852 160 -452 200
rect -110 1530 1290 1570
rect -110 210 -70 1530
rect 1250 210 1290 1530
rect -110 170 1290 210
rect -1852 -200 -452 -160
rect -1852 -1520 -1812 -200
rect -492 -1520 -452 -200
rect -1852 -1560 -452 -1520
rect -110 -190 1290 -150
rect -110 -1510 -70 -190
rect 1250 -1510 1290 -190
rect -110 -1550 1290 -1510
<< mimcapcontact >>
rect -1812 200 -492 1520
rect -70 210 1250 1530
rect -1812 -1520 -492 -200
rect -70 -1510 1250 -190
<< metal4 >>
rect -1204 1521 -1100 1614
rect 538 1531 642 1624
rect -71 1530 1251 1531
rect -1813 1520 -491 1521
rect -1813 200 -1812 1520
rect -492 200 -491 1520
rect -71 210 -70 1530
rect 1250 210 1251 1530
rect -71 209 1251 210
rect -1813 199 -491 200
rect -1204 -199 -1100 199
rect 538 -189 642 209
rect -71 -190 1251 -189
rect -1813 -200 -491 -199
rect -1813 -1520 -1812 -200
rect -492 -1520 -491 -200
rect -71 -1510 -70 -190
rect 1250 -1510 1251 -190
rect -71 -1511 1251 -1510
rect -1813 -1521 -491 -1520
rect -1204 -1614 -1100 -1521
rect 538 -1604 642 -1511
<< properties >>
string FIXED_BBOX 120 120 1600 1600
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 6.999 l 6.999 val 103.318 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
