* NGSPICE file created from sky130_be_ip__lsxo.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p35_WHP78W a_131_6584# a_n367_6584# a_n1031_n7016#
+ a_961_n7016# a_n201_n7016# a_n699_n7016# a_n865_6584# a_463_n7016# a_463_6584# a_n699_6584#
+ a_n1197_6584# a_297_6584# a_1127_n7016# a_n533_n7016# a_961_6584# a_n35_n7016# a_795_n7016#
+ a_795_6584# a_n201_6584# a_629_6584# a_297_n7016# a_629_n7016# a_n35_6584# a_n865_n7016#
+ a_n1197_n7016# a_n367_n7016# a_n533_6584# a_n1327_n7146# a_131_n7016# a_n1031_6584#
+ a_1127_6584#
X0 a_n699_6584# a_n699_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X1 a_131_6584# a_131_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X2 a_n1197_6584# a_n1197_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X3 a_n533_6584# a_n533_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X4 a_1127_6584# a_1127_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X5 a_463_6584# a_463_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X6 a_629_6584# a_629_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X7 a_n1031_6584# a_n1031_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X8 a_n35_6584# a_n35_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X9 a_961_6584# a_961_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X10 a_n367_6584# a_n367_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X11 a_297_6584# a_297_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X12 a_n865_6584# a_n865_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X13 a_795_6584# a_795_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X14 a_n201_6584# a_n201_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
C0 a_131_6584# a_n35_6584# 0.296258f
C1 a_n1197_6584# a_n1031_6584# 0.296258f
C2 a_n699_n7016# a_n533_n7016# 0.296258f
C3 a_1127_n7016# a_961_n7016# 0.296258f
C4 a_961_n7016# a_795_n7016# 0.296258f
C5 a_n865_n7016# a_n1031_n7016# 0.296258f
C6 a_n201_n7016# a_n367_n7016# 0.296258f
C7 a_n1197_n7016# a_n1031_n7016# 0.296258f
C8 a_795_6584# a_961_6584# 0.296258f
C9 a_463_n7016# a_297_n7016# 0.296258f
C10 a_629_n7016# a_795_n7016# 0.296258f
C11 a_n865_n7016# a_n699_n7016# 0.296258f
C12 a_n367_6584# a_n533_6584# 0.296258f
C13 a_795_6584# a_629_6584# 0.296258f
C14 a_n1031_6584# a_n865_6584# 0.296258f
C15 a_629_6584# a_463_6584# 0.296258f
C16 a_n367_n7016# a_n533_n7016# 0.296258f
C17 a_n201_6584# a_n367_6584# 0.296258f
C18 a_297_6584# a_463_6584# 0.296258f
C19 a_n699_6584# a_n533_6584# 0.296258f
C20 a_n35_n7016# a_n201_n7016# 0.296258f
C21 a_n699_6584# a_n865_6584# 0.296258f
C22 a_1127_6584# a_961_6584# 0.296258f
C23 a_629_n7016# a_463_n7016# 0.296258f
C24 a_297_6584# a_131_6584# 0.296258f
C25 a_n35_6584# a_n201_6584# 0.296258f
C26 a_297_n7016# a_131_n7016# 0.296258f
C27 a_n35_n7016# a_131_n7016# 0.296258f
C28 a_1127_n7016# a_n1327_n7146# 0.387223f
C29 a_1127_6584# a_n1327_n7146# 0.387223f
C30 a_961_n7016# a_n1327_n7146# 0.17691f
C31 a_961_6584# a_n1327_n7146# 0.17691f
C32 a_795_n7016# a_n1327_n7146# 0.17691f
C33 a_795_6584# a_n1327_n7146# 0.17691f
C34 a_629_n7016# a_n1327_n7146# 0.17691f
C35 a_629_6584# a_n1327_n7146# 0.17691f
C36 a_463_n7016# a_n1327_n7146# 0.17691f
C37 a_463_6584# a_n1327_n7146# 0.17691f
C38 a_297_n7016# a_n1327_n7146# 0.17691f
C39 a_297_6584# a_n1327_n7146# 0.17691f
C40 a_131_n7016# a_n1327_n7146# 0.17691f
C41 a_131_6584# a_n1327_n7146# 0.17691f
C42 a_n35_n7016# a_n1327_n7146# 0.17691f
C43 a_n35_6584# a_n1327_n7146# 0.17691f
C44 a_n201_n7016# a_n1327_n7146# 0.17691f
C45 a_n201_6584# a_n1327_n7146# 0.17691f
C46 a_n367_n7016# a_n1327_n7146# 0.17691f
C47 a_n367_6584# a_n1327_n7146# 0.17691f
C48 a_n533_n7016# a_n1327_n7146# 0.17691f
C49 a_n533_6584# a_n1327_n7146# 0.17691f
C50 a_n699_n7016# a_n1327_n7146# 0.17691f
C51 a_n699_6584# a_n1327_n7146# 0.17691f
C52 a_n865_n7016# a_n1327_n7146# 0.17691f
C53 a_n865_6584# a_n1327_n7146# 0.17691f
C54 a_n1031_n7016# a_n1327_n7146# 0.17691f
C55 a_n1031_6584# a_n1327_n7146# 0.17691f
C56 a_n1197_n7016# a_n1327_n7146# 0.387223f
C57 a_n1197_6584# a_n1327_n7146# 0.387223f
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_M35ED8 a_1210_n8616# a_546_8184# a_878_n8616#
+ a_n118_n8616# a_1210_8184# a_n450_8184# a_n1944_8184# a_n1778_n8616# a_1044_8184#
+ a_n284_8184# a_n948_n8616# a_n1778_8184# a_878_8184# a_380_n8616# a_1542_n8616#
+ a_712_n8616# a_2040_8184# a_n1280_n8616# a_2040_n8616# a_1542_8184# a_n118_8184#
+ a_n1612_n8616# a_n450_n8616# a_1044_n8616# a_214_n8616# a_n782_8184# a_1376_8184#
+ a_n1280_8184# a_n2110_n8616# a_380_8184# a_n1114_n8616# a_n616_8184# a_1874_n8616#
+ a_n1114_8184# a_48_n8616# a_214_8184# a_1874_8184# a_n1944_n8616# a_1376_n8616#
+ a_n782_n8616# a_546_n8616# a_n2110_8184# a_1708_n8616# a_1708_8184# a_48_8184# a_n1612_8184#
+ a_n1446_n8616# a_n2240_n8746# a_712_8184# a_n284_n8616# a_n948_8184# a_n616_n8616#
+ a_n1446_8184#
X0 a_n616_8184# a_n616_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X1 a_1044_8184# a_1044_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X2 a_546_8184# a_546_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X3 a_380_8184# a_380_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X4 a_n1114_8184# a_n1114_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X5 a_1708_8184# a_1708_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X6 a_1542_8184# a_1542_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X7 a_2040_8184# a_2040_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X8 a_n450_8184# a_n450_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X9 a_n1612_8184# a_n1612_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X10 a_n284_8184# a_n284_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X11 a_48_8184# a_48_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X12 a_n948_8184# a_n948_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X13 a_n782_8184# a_n782_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X14 a_1376_8184# a_1376_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X15 a_878_8184# a_878_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X16 a_n1446_8184# a_n1446_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X17 a_n2110_8184# a_n2110_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X18 a_1874_8184# a_1874_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X19 a_n1944_8184# a_n1944_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X20 a_214_8184# a_214_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X21 a_n1280_8184# a_n1280_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X22 a_1210_8184# a_1210_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X23 a_712_8184# a_712_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X24 a_n118_8184# a_n118_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X25 a_n1778_8184# a_n1778_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
C0 a_1210_n8616# a_1376_n8616# 0.296258f
C1 a_n450_8184# a_n616_8184# 0.296258f
C2 a_1542_8184# a_1708_8184# 0.296258f
C3 a_878_8184# a_1044_8184# 0.296258f
C4 a_1874_n8616# a_1708_n8616# 0.296258f
C5 a_2040_n8616# a_1874_n8616# 0.296258f
C6 a_n1944_8184# a_n1778_8184# 0.296258f
C7 a_n1944_n8616# a_n2110_n8616# 0.296258f
C8 a_n1944_n8616# a_n1778_n8616# 0.296258f
C9 a_n118_n8616# a_n284_n8616# 0.296258f
C10 a_n948_8184# a_n782_8184# 0.296258f
C11 a_n616_n8616# a_n782_n8616# 0.296258f
C12 a_n118_n8616# a_48_n8616# 0.296258f
C13 a_n450_n8616# a_n616_n8616# 0.296258f
C14 a_214_8184# a_380_8184# 0.296258f
C15 a_1210_8184# a_1376_8184# 0.296258f
C16 a_n1280_n8616# a_n1446_n8616# 0.296258f
C17 a_1542_8184# a_1376_8184# 0.296258f
C18 a_1044_n8616# a_1210_n8616# 0.296258f
C19 a_712_8184# a_546_8184# 0.296258f
C20 a_n948_8184# a_n1114_8184# 0.296258f
C21 a_214_n8616# a_48_n8616# 0.296258f
C22 a_2040_8184# a_1874_8184# 0.296258f
C23 a_878_n8616# a_1044_n8616# 0.296258f
C24 a_214_n8616# a_380_n8616# 0.296258f
C25 a_n118_8184# a_n284_8184# 0.296258f
C26 a_n450_n8616# a_n284_n8616# 0.296258f
C27 a_n1114_n8616# a_n948_n8616# 0.296258f
C28 a_380_8184# a_546_8184# 0.296258f
C29 a_n782_n8616# a_n948_n8616# 0.296258f
C30 a_878_8184# a_712_8184# 0.296258f
C31 a_n616_8184# a_n782_8184# 0.296258f
C32 a_1542_n8616# a_1376_n8616# 0.296258f
C33 a_n1446_8184# a_n1280_8184# 0.296258f
C34 a_1210_8184# a_1044_8184# 0.296258f
C35 a_n1612_n8616# a_n1446_n8616# 0.296258f
C36 a_214_8184# a_48_8184# 0.296258f
C37 a_n1944_8184# a_n2110_8184# 0.296258f
C38 a_n1446_8184# a_n1612_8184# 0.296258f
C39 a_n1114_n8616# a_n1280_n8616# 0.296258f
C40 a_n1612_n8616# a_n1778_n8616# 0.296258f
C41 a_n450_8184# a_n284_8184# 0.296258f
C42 a_n1280_8184# a_n1114_8184# 0.296258f
C43 a_n1778_8184# a_n1612_8184# 0.296258f
C44 a_n118_8184# a_48_8184# 0.296258f
C45 a_712_n8616# a_546_n8616# 0.296258f
C46 a_878_n8616# a_712_n8616# 0.296258f
C47 a_1708_8184# a_1874_8184# 0.296258f
C48 a_1542_n8616# a_1708_n8616# 0.296258f
C49 a_380_n8616# a_546_n8616# 0.296258f
C50 a_2040_n8616# a_n2240_n8746# 0.387223f
C51 a_2040_8184# a_n2240_n8746# 0.387223f
C52 a_1874_n8616# a_n2240_n8746# 0.17691f
C53 a_1874_8184# a_n2240_n8746# 0.17691f
C54 a_1708_n8616# a_n2240_n8746# 0.17691f
C55 a_1708_8184# a_n2240_n8746# 0.17691f
C56 a_1542_n8616# a_n2240_n8746# 0.17691f
C57 a_1542_8184# a_n2240_n8746# 0.17691f
C58 a_1376_n8616# a_n2240_n8746# 0.17691f
C59 a_1376_8184# a_n2240_n8746# 0.17691f
C60 a_1210_n8616# a_n2240_n8746# 0.17691f
C61 a_1210_8184# a_n2240_n8746# 0.17691f
C62 a_1044_n8616# a_n2240_n8746# 0.17691f
C63 a_1044_8184# a_n2240_n8746# 0.17691f
C64 a_878_n8616# a_n2240_n8746# 0.17691f
C65 a_878_8184# a_n2240_n8746# 0.17691f
C66 a_712_n8616# a_n2240_n8746# 0.17691f
C67 a_712_8184# a_n2240_n8746# 0.17691f
C68 a_546_n8616# a_n2240_n8746# 0.17691f
C69 a_546_8184# a_n2240_n8746# 0.17691f
C70 a_380_n8616# a_n2240_n8746# 0.17691f
C71 a_380_8184# a_n2240_n8746# 0.17691f
C72 a_214_n8616# a_n2240_n8746# 0.17691f
C73 a_214_8184# a_n2240_n8746# 0.17691f
C74 a_48_n8616# a_n2240_n8746# 0.17691f
C75 a_48_8184# a_n2240_n8746# 0.17691f
C76 a_n118_n8616# a_n2240_n8746# 0.17691f
C77 a_n118_8184# a_n2240_n8746# 0.17691f
C78 a_n284_n8616# a_n2240_n8746# 0.17691f
C79 a_n284_8184# a_n2240_n8746# 0.17691f
C80 a_n450_n8616# a_n2240_n8746# 0.17691f
C81 a_n450_8184# a_n2240_n8746# 0.17691f
C82 a_n616_n8616# a_n2240_n8746# 0.17691f
C83 a_n616_8184# a_n2240_n8746# 0.17691f
C84 a_n782_n8616# a_n2240_n8746# 0.17691f
C85 a_n782_8184# a_n2240_n8746# 0.17691f
C86 a_n948_n8616# a_n2240_n8746# 0.17691f
C87 a_n948_8184# a_n2240_n8746# 0.17691f
C88 a_n1114_n8616# a_n2240_n8746# 0.17691f
C89 a_n1114_8184# a_n2240_n8746# 0.17691f
C90 a_n1280_n8616# a_n2240_n8746# 0.17691f
C91 a_n1280_8184# a_n2240_n8746# 0.17691f
C92 a_n1446_n8616# a_n2240_n8746# 0.17691f
C93 a_n1446_8184# a_n2240_n8746# 0.17691f
C94 a_n1612_n8616# a_n2240_n8746# 0.17691f
C95 a_n1612_8184# a_n2240_n8746# 0.17691f
C96 a_n1778_n8616# a_n2240_n8746# 0.17691f
C97 a_n1778_8184# a_n2240_n8746# 0.17691f
C98 a_n1944_n8616# a_n2240_n8746# 0.17691f
C99 a_n1944_8184# a_n2240_n8746# 0.17691f
C100 a_n2110_n8616# a_n2240_n8746# 0.387223f
C101 a_n2110_8184# a_n2240_n8746# 0.387223f
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
C0 A a_27_47# 0.181449f
C1 VPWR a_27_47# 0.135101f
C2 X a_27_47# 0.107446f
C3 VGND a_27_47# 0.104759f
C4 VGND VNB 0.207322f
C5 VPWR VNB 0.175402f
C6 A VNB 0.164055f
C7 VPB VNB 0.338976f
C8 a_27_47# VNB 0.207781f
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_VTNT3C a_n118_7484# a_214_n7916# a_48_n7916#
+ a_214_7484# a_n414_n8046# a_48_7484# a_n284_n7916# a_n118_n7916# a_n284_7484#
X0 a_n284_7484# a_n284_n7916# a_n414_n8046# sky130_fd_pr__res_xhigh_po_0p35 l=75
X1 a_48_7484# a_48_n7916# a_n414_n8046# sky130_fd_pr__res_xhigh_po_0p35 l=75
X2 a_214_7484# a_214_n7916# a_n414_n8046# sky130_fd_pr__res_xhigh_po_0p35 l=75
X3 a_n118_7484# a_n118_n7916# a_n414_n8046# sky130_fd_pr__res_xhigh_po_0p35 l=75
C0 a_n118_n7916# a_n284_n7916# 0.296258f
C1 a_214_n7916# a_48_n7916# 0.296258f
C2 a_n118_7484# a_n284_7484# 0.296258f
C3 a_48_7484# a_n118_7484# 0.296258f
C4 a_48_7484# a_214_7484# 0.296258f
C5 a_n118_n7916# a_48_n7916# 0.296258f
C6 a_214_n7916# a_n414_n8046# 0.387223f
C7 a_214_7484# a_n414_n8046# 0.387223f
C8 a_48_n7916# a_n414_n8046# 0.17691f
C9 a_48_7484# a_n414_n8046# 0.17691f
C10 a_n118_n7916# a_n414_n8046# 0.17691f
C11 a_n118_7484# a_n414_n8046# 0.17691f
C12 a_n284_n7916# a_n414_n8046# 0.387223f
C13 a_n284_7484# a_n414_n8046# 0.387223f
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RJ a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
C0 a_n45_n45# a_n147_n147# 0.169345f
.ends

.subckt sky130_fd_pr__nfet_01v8_LHQHT5 a_n29_n400# a_887_n400# a_429_n400# a_n887_n488#
+ a_n1047_n574# a_n429_n488# a_487_n488# a_n945_n400# a_29_n488# a_n487_n400#
X0 a_n487_n400# a_n887_n488# a_n945_n400# a_n1047_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=2
X1 a_n29_n400# a_n429_n488# a_n487_n400# a_n1047_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X2 a_429_n400# a_29_n488# a_n29_n400# a_n1047_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X3 a_887_n400# a_487_n488# a_429_n400# a_n1047_n574# sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=2
C0 a_887_n400# a_n1047_n574# 0.336596f
C1 a_429_n400# a_n1047_n574# 0.216749f
C2 a_n29_n400# a_n1047_n574# 0.216749f
C3 a_n487_n400# a_n1047_n574# 0.216749f
C4 a_n945_n400# a_n1047_n574# 0.336596f
C5 a_487_n488# a_n1047_n574# 1.23765f
C6 a_29_n488# a_n1047_n574# 1.17381f
C7 a_n429_n488# a_n1047_n574# 1.17381f
C8 a_n887_n488# a_n1047_n574# 1.23765f
.ends

.subckt sky130_fd_pr__nfet_01v8_69TQ3K a_n260_n274# a_100_n100# a_n158_n100# a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n260_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_100_n100# a_n260_n274# 0.146358f
C1 a_n158_n100# a_n260_n274# 0.146358f
C2 a_n100_n188# a_n260_n274# 0.724275f
.ends

.subckt sky130_fd_pr__pfet_01v8_3HMWVM 0. w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 w_n296_n319# a_n100_n197# 0.434431f
C1 a_n100_n197# 0. 0.310981f
C2 w_n296_n319# 0. 1.64714f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B a_29_n388# a_n129_n388# a_n321_n522# a_n29_n300#
+ a_n187_n300# a_129_n300#
X0 a_129_n300# a_29_n388# a_n29_n300# a_n321_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X1 a_n29_n300# a_n129_n388# a_n187_n300# a_n321_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
C0 a_n129_n388# a_29_n388# 0.104496f
C1 a_n29_n300# a_129_n300# 0.268329f
C2 a_n29_n300# a_n187_n300# 0.268329f
C3 a_129_n300# a_n321_n522# 0.329514f
C4 a_n187_n300# a_n321_n522# 0.329514f
C5 a_29_n388# a_n321_n522# 0.368192f
C6 a_n129_n388# a_n321_n522# 0.368192f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_VHBZVD 0. a_n400_n197# a_400_n100# w_n658_n397#
+ a_n458_n100#
X0 a_400_n100# a_n400_n197# a_n458_n100# w_n658_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
C0 w_n658_n397# a_n400_n197# 1.31949f
C1 a_n400_n197# 0. 1.01545f
C2 w_n658_n397# 0. 4.01834f
.ends

.subckt level_shift dvdd 0. in in_b out_b out dw_2668_n1758# avss avdd
XXM1 0. in_b 0. in sky130_fd_pr__nfet_01v8_69TQ3K
XXM2 0. dvdd in dvdd in_b sky130_fd_pr__pfet_01v8_3HMWVM
XXM3 in in avss out_b avss avss sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B
XXM4 in_b in_b avss out avss avss sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B
XXM5 0. out avdd avdd out_b sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
XXM6 0. out_b out avdd avdd sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
C0 out_b out 0.606335f
C1 out_b avdd 2.455349f
C2 out in_b 0.852906f
C3 avdd out 2.447048f
C4 avss in 1.40922f
C5 avss out_b 0.796108f
C6 avss in_b 1.423692f
C7 avss dw_2668_n1758# 4.93164f
C8 avss out 0.85934f
C9 avss avdd 0.861367f
C10 out_b in 0.84957f
C11 in dvdd 0.370698f
C12 in in_b 0.605523f
C13 avss 0. 1.518337f
C14 dw_2668_n1758# 0. 4.93164f
C15 avdd 0. 8.316299f
C16 out 0. 1.155064f
C17 in_b 0. 1.345128f
C18 out_b 0. 1.23154f
C19 in 0. 2.261764f
C20 dvdd 0. 2.21807f
.ends

.subckt sky130_fd_pr__nfet_01v8_6G4XAN a_n29_n155# a_29_n243# a_n287_n155# a_n389_n329#
+ a_n229_n243# a_229_55# a_229_n155# a_n287_55# a_n29_55#
X0 a_n29_n155# a_n229_n243# a_n287_n155# a_n389_n329# sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X1 a_229_n155# a_29_n243# a_n29_n155# a_n389_n329# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X2 a_229_55# a_29_n243# a_n29_55# a_n389_n329# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X3 a_n29_55# a_n229_n243# a_n287_55# a_n389_n329# sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
C0 a_29_n243# a_n229_n243# 0.155031f
C1 a_29_n243# a_n389_n329# 0.884838f
C2 a_n229_n243# a_n389_n329# 0.884838f
.ends

.subckt sky130_fd_sc_hd__and2_0 A B VGND VNB VPB VPWR X
X0 VPWR B a_40_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_40_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X2 VGND B a_123_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_40_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X4 a_123_47# A a_40_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 a_40_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
C0 A B 0.117044f
C1 VPWR X 0.111278f
C2 B a_40_47# 0.206108f
C3 VGND X 0.105358f
C4 VPWR a_40_47# 0.141098f
C5 X a_40_47# 0.11426f
C6 A a_40_47# 0.12536f
C7 VGND a_40_47# 0.138964f
C8 VGND VNB 0.300193f
C9 X VNB 0.10272f
C10 VPWR VNB 0.262881f
C11 B VNB 0.121465f
C12 A VNB 0.194569f
C13 VPB VNB 0.516168f
C14 a_40_47# VNB 0.230074f
.ends

.subckt sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N a_1847_47#
+ a_193_47# a_27_47#
X0 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2 VPWR a_1283_21# a_1847_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 Q_N a_1847_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND a_1283_21# a_1847_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X13 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X17 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X18 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X19 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X20 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X26 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X27 Q_N a_1847_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X28 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X29 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
C0 VPWR a_1847_47# 0.153243f
C1 D VPB 0.137565f
C2 a_27_47# RESET_B 0.296336f
C3 a_1283_21# RESET_B 0.278608f
C4 a_27_47# a_543_47# 0.115353f
C5 VPWR VPB 0.235545f
C6 D a_27_47# 0.132849f
C7 a_27_47# VPWR 0.152297f
C8 VPWR a_1283_21# 0.161911f
C9 a_1108_47# RESET_B 0.236601f
C10 VPWR a_1108_47# 0.171246f
C11 VGND RESET_B 0.288101f
C12 a_761_289# RESET_B 0.166114f
C13 VGND a_543_47# 0.122935f
C14 a_761_289# a_543_47# 0.209641f
C15 a_761_289# VPWR 0.10497f
C16 a_193_47# VPB 0.170766f
C17 a_27_47# a_193_47# 0.906454f
C18 a_543_47# RESET_B 0.153272f
C19 a_1108_47# a_193_47# 0.125324f
C20 VPWR a_543_47# 0.100285f
C21 a_761_289# a_193_47# 0.186387f
C22 a_651_413# VPWR 0.12856f
C23 a_1847_47# a_1283_21# 0.106826f
C24 a_27_47# VPB 0.261876f
C25 a_1283_21# VPB 0.246515f
C26 a_543_47# a_193_47# 0.229804f
C27 D a_193_47# 0.217945f
C28 VPWR a_193_47# 0.396049f
C29 a_1108_47# VPB 0.112685f
C30 a_27_47# a_1108_47# 0.102355f
C31 a_1108_47# a_1283_21# 0.251137f
C32 a_27_47# CLK 0.233602f
C33 a_27_47# VGND 0.253982f
C34 Q a_1847_47# 0.161495f
C35 VGND a_1283_21# 0.266204f
C36 Q a_1283_21# 0.119961f
C37 VGND a_1108_47# 0.148194f
C38 D a_448_47# 0.155634f
C39 VPB RESET_B 0.138482f
C40 VGND VNB 1.17272f
C41 VPWR VNB 0.959088f
C42 RESET_B VNB 0.260061f
C43 D VNB 0.159894f
C44 CLK VNB 0.195254f
C45 VPB VNB 2.1109f
C46 a_1847_47# VNB 0.132899f
C47 a_1108_47# VNB 0.126214f
C48 a_1283_21# VNB 0.478567f
C49 a_543_47# VNB 0.157869f
C50 a_761_289# VNB 0.120848f
C51 a_193_47# VNB 0.272684f
C52 a_27_47# VNB 0.495665f
.ends

.subckt ripple_dly_4 clkin doneb x2/a_27_47# Qb2 x3/a_27_47# ena x2/a_193_47# x4/a_27_47#
+ 0. Qb1 dvdd
Xx1 clkin doneb 0. 0. dvdd dvdd x1/X sky130_fd_sc_hd__and2_0
Xx3 Qb1 Qb2 ena 0. 0. dvdd dvdd x3/Q Qb2 x3/a_1847_47# x3/a_193_47# x3/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xx2 x1/X Qb1 ena 0. 0. dvdd dvdd x2/Q Qb1 x2/a_1847_47# x2/a_193_47# x2/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xx4 Qb2 doneb ena 0. 0. dvdd dvdd x4/Q doneb x4/a_1847_47# x4/a_193_47# x4/a_27_47#
+ sky130_fd_sc_hd__dfrbp_1
C0 ena x4/a_27_47# 0.317074f
C1 x3/a_27_47# x3/a_193_47# -0.298091f
C2 ena x3/a_27_47# 0.317225f
C3 doneb x2/a_193_47# 0.202238f
C4 x2/a_27_47# Qb1 0.497822f
C5 dvdd x1/X 0.143961f
C6 x2/a_27_47# 0. -0.108344f
C7 doneb Qb2 0.141763f
C8 ena Qb1 0.34662f
C9 x4/a_27_47# 0. -0.10834f
C10 doneb x4/a_193_47# 0.74189f
C11 ena 0. 2.192297f
C12 doneb x4/a_1847_47# 0.11114f
C13 x3/a_27_47# 0. -0.10834f
C14 x2/a_27_47# x2/a_193_47# -0.298092f
C15 ena clkin 0.125078f
C16 Qb1 dvdd 0.364399f
C17 doneb x3/a_193_47# 0.199885f
C18 doneb x4/a_27_47# 0.542089f
C19 0. dvdd -0.376178f
C20 ena doneb 0.328336f
C21 Qb2 x3/a_193_47# 0.538587f
C22 ena Qb2 0.346581f
C23 x4/a_27_47# x4/a_193_47# -0.298091f
C24 x3/a_27_47# Qb2 0.497823f
C25 clkin dvdd 0.183034f
C26 doneb x4/a_1283_21# 0.107576f
C27 x2/a_193_47# Qb1 0.538585f
C28 doneb Qb1 0.142549f
C29 doneb 0. 0.217949f
C30 doneb dvdd 2.074138f
C31 ena x2/a_27_47# 0.31541f
C32 Qb2 dvdd 0.364487f
C33 x4/a_1847_47# 0 0.132899f
C34 x4/a_1108_47# 0 0.126214f $ **FLOATING
C35 x4/a_1283_21# 0 0.478567f $ **FLOATING
C36 x4/a_543_47# 0 0.157869f $ **FLOATING
C37 x4/a_761_289# 0 0.120848f $ **FLOATING
C38 x4/a_193_47# 0 0.272684f
C39 x4/a_27_47# 0 0.495665f
C40 0. 0 3.076656f
C41 dvdd 0 9.8956f
C42 ena 0 0.978923f
C43 Qb1 0 0.335308f
C44 x1/X 0 0.180099f
C45 x2/a_1847_47# 0 0.132899f
C46 x2/a_1108_47# 0 0.126214f $ **FLOATING
C47 x2/a_1283_21# 0 0.478567f $ **FLOATING
C48 x2/a_543_47# 0 0.157869f $ **FLOATING
C49 x2/a_761_289# 0 0.120848f $ **FLOATING
C50 x2/a_193_47# 0 0.272684f
C51 x2/a_27_47# 0 0.495665f
C52 Qb2 0 0.335611f
C53 x3/a_1847_47# 0 0.132899f
C54 x3/a_1108_47# 0 0.126214f $ **FLOATING
C55 x3/a_1283_21# 0 0.478567f $ **FLOATING
C56 x3/a_543_47# 0 0.157869f $ **FLOATING
C57 x3/a_761_289# 0 0.120848f $ **FLOATING
C58 x3/a_193_47# 0 0.272684f
C59 x3/a_27_47# 0 0.495665f
C60 doneb 0 1.588155f
C61 clkin 0 0.301494f
C62 x1/a_40_47# 0 0.230074f $ **FLOATING
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
C0 a_193_297# a_27_47# 0.143754f
C1 a_193_297# VPWR 0.169243f
C2 a_27_47# VGND 0.395423f
C3 a_27_47# A2 0.152957f
C4 a_109_297# VPWR 0.150131f
C5 B1 a_27_47# 0.11237f
C6 VGND VNB 0.437277f
C7 VPWR VNB 0.363959f
C8 A1 VNB 0.105908f
C9 B1 VNB 0.108471f
C10 C1 VNB 0.139233f
C11 VPB VNB 0.781956f
C12 a_27_47# VNB 0.216317f
.ends

.subckt sky130_fd_sc_hd__einvn_0 A TE_B VGND VNB VPB VPWR Z a_30_47#
X0 VGND TE_B a_30_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07665 pd=0.785 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 Z A a_215_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0672 ps=0.85 w=0.64 l=0.15
X2 a_215_369# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.10855 ps=1.005 w=0.64 l=0.15
X3 a_215_47# a_30_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.07665 ps=0.785 w=0.42 l=0.15
X4 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR TE_B a_30_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.005 as=0.1092 ps=1.36 w=0.42 l=0.15
C0 Z A 0.188537f
C1 a_30_47# VPWR 0.116195f
C2 a_30_47# VGND 0.124215f
C3 TE_B VPB 0.136539f
C4 a_30_47# Z 0.133869f
C5 a_30_47# TE_B 0.265521f
C6 VGND VNB 0.251746f
C7 VPWR VNB 0.213824f
C8 A VNB 0.206932f
C9 TE_B VNB 0.220088f
C10 VPB VNB 0.427572f
C11 a_30_47# VNB 0.145562f
.ends

.subckt sky130_fd_pr__nfet_01v8_AHZR5K a_n458_n50# a_n400_n138# a_n560_n224# a_400_n50#
X0 a_400_n50# a_n400_n138# a_n458_n50# a_n560_n224# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
C0 a_n400_n138# a_n560_n224# 2.37082f
.ends

.subckt ripl_dly_clk_buf clkin stby x1/x2/a_27_47# x2/x2/a_27_47# x1/x3/a_27_47# x2/x3/a_27_47#
+ x2/Qb1 x1/Qb1 x1/x4/a_27_47# x2/x4/a_27_47# x2/Qb2 ena_done_b stby_done_b clk_disable
+ clkout ena x1/Qb2 dvss x5/VPB stby_b x1/x2/a_193_47#
Xx1 clkin ena_done_b x1/x2/a_27_47# x1/Qb2 x1/x3/a_27_47# ena x1/x2/a_193_47# x1/x4/a_27_47#
+ dvss x1/Qb1 x5/VPB ripple_dly_4
Xx2 clkin stby_done_b x2/x2/a_27_47# x2/Qb2 x2/x3/a_27_47# stby_b x2/x2/a_193_47#
+ x2/x4/a_27_47# dvss x2/Qb1 x5/VPB ripple_dly_4
Xx3 stby_b stby_done_b ena ena_done_b stby dvss dvss x5/VPB x5/VPB clk_disable sky130_fd_sc_hd__a221o_1
Xx5 clkin clk_disable dvss dvss x5/VPB x5/VPB clkout x5/a_30_47# sky130_fd_sc_hd__einvn_0
XXM3 clkout clk_disable dvss dvss sky130_fd_pr__nfet_01v8_AHZR5K
C0 stby_done_b clkout 0.187099f
C1 stby_b ena 0.664996f
C2 clk_disable clkin 0.106197f
C3 stby_done_b x5/VPB 0.451845f
C4 dvss stby 0.278618f
C5 clk_disable x5/a_30_47# 0.15444f
C6 dvss stby_b 0.136205f
C7 ena ena_done_b 0.394686f
C8 dvss clk_disable 0.410059f
C9 stby_done_b stby_b 0.449182f
C10 clk_disable clkout 0.458364f
C11 stby_b x5/VPB 0.337201f
C12 stby_done_b clk_disable 0.72273f
C13 clk_disable x5/VPB 0.111141f
C14 dvss ena 0.146489f
C15 clkin clkout 0.624163f
C16 dvss ena_done_b 0.353487f
C17 x5/VPB clkin 0.550211f
C18 x5/VPB ena 0.173428f
C19 stby_done_b ena_done_b 1.608666f
C20 x5/VPB ena_done_b 0.713195f
C21 stby_done_b dvss 0.277332f
C22 dvss x5/VPB 1.081624f
C23 stby_b clkin 0.188961f
C24 clkout 0 0.628268f
C25 clk_disable 0 2.783535f
C26 x5/a_30_47# 0 0.145562f
C27 stby 0 0.668001f
C28 x3/a_27_47# 0 0.216317f $ **FLOATING
C29 x2/x4/a_1847_47# 0 0.132899f
C30 x2/x4/a_1108_47# 0 0.126214f $ **FLOATING
C31 x2/x4/a_1283_21# 0 0.478567f $ **FLOATING
C32 x2/x4/a_543_47# 0 0.157869f $ **FLOATING
C33 x2/x4/a_761_289# 0 0.120848f $ **FLOATING
C34 x2/x4/a_193_47# 0 0.272684f
C35 x2/x4/a_27_47# 0 0.495665f
C36 x5/VPB 0 14.113154f
C37 stby_b 0 1.158189f
C38 x2/Qb1 0 0.335308f
C39 x2/x1/X 0 0.180099f
C40 x2/x2/a_1847_47# 0 0.132899f
C41 x2/x2/a_1108_47# 0 0.126214f $ **FLOATING
C42 x2/x2/a_1283_21# 0 0.478567f $ **FLOATING
C43 x2/x2/a_543_47# 0 0.157869f $ **FLOATING
C44 x2/x2/a_761_289# 0 0.120848f $ **FLOATING
C45 x2/x2/a_193_47# 0 0.272684f
C46 x2/x2/a_27_47# 0 0.495665f
C47 x2/Qb2 0 0.335611f
C48 x2/x3/a_1847_47# 0 0.132899f
C49 x2/x3/a_1108_47# 0 0.126214f $ **FLOATING
C50 x2/x3/a_1283_21# 0 0.478567f $ **FLOATING
C51 x2/x3/a_543_47# 0 0.157869f $ **FLOATING
C52 x2/x3/a_761_289# 0 0.120848f $ **FLOATING
C53 x2/x3/a_193_47# 0 0.272684f
C54 x2/x3/a_27_47# 0 0.495665f
C55 stby_done_b 0 1.263094f
C56 clkin 0 1.465572f
C57 x2/x1/a_40_47# 0 0.230074f $ **FLOATING
C58 x1/x4/a_1847_47# 0 0.132899f
C59 x1/x4/a_1108_47# 0 0.126214f $ **FLOATING
C60 x1/x4/a_1283_21# 0 0.478567f $ **FLOATING
C61 x1/x4/a_543_47# 0 0.157869f $ **FLOATING
C62 x1/x4/a_761_289# 0 0.120848f $ **FLOATING
C63 x1/x4/a_193_47# 0 0.272684f
C64 x1/x4/a_27_47# 0 0.495665f
C65 dvss 0 7.210984f
C66 ena 0 1.117279f
C67 x1/Qb1 0 0.335308f
C68 x1/x1/X 0 0.180099f
C69 x1/x2/a_1847_47# 0 0.132899f
C70 x1/x2/a_1108_47# 0 0.126214f $ **FLOATING
C71 x1/x2/a_1283_21# 0 0.478567f $ **FLOATING
C72 x1/x2/a_543_47# 0 0.157869f $ **FLOATING
C73 x1/x2/a_761_289# 0 0.120848f $ **FLOATING
C74 x1/x2/a_193_47# 0 0.272684f
C75 x1/x2/a_27_47# 0 0.495665f
C76 x1/Qb2 0 0.335611f
C77 x1/x3/a_1847_47# 0 0.132899f
C78 x1/x3/a_1108_47# 0 0.126214f $ **FLOATING
C79 x1/x3/a_1283_21# 0 0.478567f $ **FLOATING
C80 x1/x3/a_543_47# 0 0.157869f $ **FLOATING
C81 x1/x3/a_761_289# 0 0.120848f $ **FLOATING
C82 x1/x3/a_193_47# 0 0.272684f
C83 x1/x3/a_27_47# 0 0.495665f
C84 ena_done_b 0 1.398332f
C85 x1/x1/a_40_47# 0 0.230074f $ **FLOATING
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z a_100_n100# a_n292_n322# a_n158_n100#
+ a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n292_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_100_n100# a_n292_n322# 0.137447f
C1 a_n158_n100# a_n292_n322# 0.137447f
C2 a_n100_n188# a_n292_n322# 0.688242f
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_68VL2P a_961_n11416# a_463_10984# a_n35_n11416#
+ a_1625_10984# a_n201_n11416# a_n1197_n11416# a_n1363_10984# a_1625_n11416# a_629_n11416#
+ a_1127_10984# a_131_n11416# a_n533_10984# a_n35_10984# a_n533_n11416# a_1957_n11416#
+ a_795_10984# a_n2157_n11546# a_463_n11416# a_1957_10984# a_n865_n11416# a_n1861_n11416#
+ a_n1695_10984# a_1791_n11416# a_1127_n11416# a_795_n11416# a_297_10984# a_1459_10984#
+ a_n865_10984# a_629_10984# a_n1529_n11416# a_n1031_n11416# a_n1197_10984# a_1459_n11416#
+ a_n1529_10984# a_n367_10984# a_n367_n11416# a_131_10984# a_n1363_n11416# a_n2027_10984#
+ a_297_n11416# a_1293_n11416# a_n699_n11416# a_n1031_10984# a_1791_10984# a_n1695_n11416#
+ a_961_10984# a_n201_10984# a_n2027_n11416# a_n699_10984# a_n1861_10984# a_1293_10984#
X0 a_1957_10984# a_1957_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X1 a_n1861_10984# a_n1861_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X2 a_463_10984# a_463_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X3 a_1791_10984# a_1791_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X4 a_n35_10984# a_n35_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X5 a_795_10984# a_795_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X6 a_n2027_10984# a_n2027_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X7 a_961_10984# a_961_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X8 a_n1197_10984# a_n1197_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X9 a_n1031_10984# a_n1031_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X10 a_1127_10984# a_1127_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X11 a_n1529_10984# a_n1529_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X12 a_n367_10984# a_n367_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X13 a_n201_10984# a_n201_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X14 a_1459_10984# a_1459_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X15 a_n1363_10984# a_n1363_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X16 a_n699_10984# a_n699_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X17 a_n533_10984# a_n533_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X18 a_1293_10984# a_1293_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X19 a_n1695_10984# a_n1695_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X20 a_297_10984# a_297_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X21 a_1625_10984# a_1625_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X22 a_n865_10984# a_n865_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X23 a_131_10984# a_131_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X24 a_629_10984# a_629_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
C0 a_n699_n11416# a_n533_n11416# 0.296258f
C1 a_1791_n11416# a_1957_n11416# 0.296258f
C2 a_1791_10984# a_1957_10984# 0.296258f
C3 a_629_n11416# a_463_n11416# 0.296258f
C4 a_297_n11416# a_131_n11416# 0.296258f
C5 a_n367_10984# a_n533_10984# 0.296258f
C6 a_n367_10984# a_n201_10984# 0.296258f
C7 a_n1363_10984# a_n1529_10984# 0.296258f
C8 a_n1363_n11416# a_n1197_n11416# 0.296258f
C9 a_n865_n11416# a_n699_n11416# 0.296258f
C10 a_n1861_10984# a_n2027_10984# 0.296258f
C11 a_1459_n11416# a_1293_n11416# 0.296258f
C12 a_1127_n11416# a_1293_n11416# 0.296258f
C13 a_795_10984# a_629_10984# 0.296258f
C14 a_297_10984# a_131_10984# 0.296258f
C15 a_795_n11416# a_629_n11416# 0.296258f
C16 a_n1031_n11416# a_n865_n11416# 0.296258f
C17 a_n35_n11416# a_n201_n11416# 0.296258f
C18 a_1459_n11416# a_1625_n11416# 0.296258f
C19 a_961_n11416# a_1127_n11416# 0.296258f
C20 a_1791_n11416# a_1625_n11416# 0.296258f
C21 a_n533_10984# a_n699_10984# 0.296258f
C22 a_1625_10984# a_1459_10984# 0.296258f
C23 a_795_10984# a_961_10984# 0.296258f
C24 a_1127_10984# a_1293_10984# 0.296258f
C25 a_n35_10984# a_131_10984# 0.296258f
C26 a_n367_n11416# a_n201_n11416# 0.296258f
C27 a_n1695_10984# a_n1529_10984# 0.296258f
C28 a_n865_10984# a_n699_10984# 0.296258f
C29 a_1127_10984# a_961_10984# 0.296258f
C30 a_961_n11416# a_795_n11416# 0.296258f
C31 a_n1695_n11416# a_n1861_n11416# 0.296258f
C32 a_n1031_n11416# a_n1197_n11416# 0.296258f
C33 a_n2027_n11416# a_n1861_n11416# 0.296258f
C34 a_131_n11416# a_n35_n11416# 0.296258f
C35 a_n1197_10984# a_n1031_10984# 0.296258f
C36 a_1625_10984# a_1791_10984# 0.296258f
C37 a_463_10984# a_629_10984# 0.296258f
C38 a_n1861_10984# a_n1695_10984# 0.296258f
C39 a_1293_10984# a_1459_10984# 0.296258f
C40 a_n865_10984# a_n1031_10984# 0.296258f
C41 a_n35_10984# a_n201_10984# 0.296258f
C42 a_n1197_10984# a_n1363_10984# 0.296258f
C43 a_463_10984# a_297_10984# 0.296258f
C44 a_n1529_n11416# a_n1363_n11416# 0.296258f
C45 a_n367_n11416# a_n533_n11416# 0.296258f
C46 a_n1695_n11416# a_n1529_n11416# 0.296258f
C47 a_297_n11416# a_463_n11416# 0.296258f
C48 a_1957_n11416# a_n2157_n11546# 0.387223f
C49 a_1957_10984# a_n2157_n11546# 0.387223f
C50 a_1791_n11416# a_n2157_n11546# 0.17691f
C51 a_1791_10984# a_n2157_n11546# 0.17691f
C52 a_1625_n11416# a_n2157_n11546# 0.17691f
C53 a_1625_10984# a_n2157_n11546# 0.17691f
C54 a_1459_n11416# a_n2157_n11546# 0.17691f
C55 a_1459_10984# a_n2157_n11546# 0.17691f
C56 a_1293_n11416# a_n2157_n11546# 0.17691f
C57 a_1293_10984# a_n2157_n11546# 0.17691f
C58 a_1127_n11416# a_n2157_n11546# 0.17691f
C59 a_1127_10984# a_n2157_n11546# 0.17691f
C60 a_961_n11416# a_n2157_n11546# 0.17691f
C61 a_961_10984# a_n2157_n11546# 0.17691f
C62 a_795_n11416# a_n2157_n11546# 0.17691f
C63 a_795_10984# a_n2157_n11546# 0.17691f
C64 a_629_n11416# a_n2157_n11546# 0.17691f
C65 a_629_10984# a_n2157_n11546# 0.17691f
C66 a_463_n11416# a_n2157_n11546# 0.17691f
C67 a_463_10984# a_n2157_n11546# 0.17691f
C68 a_297_n11416# a_n2157_n11546# 0.17691f
C69 a_297_10984# a_n2157_n11546# 0.17691f
C70 a_131_n11416# a_n2157_n11546# 0.17691f
C71 a_131_10984# a_n2157_n11546# 0.17691f
C72 a_n35_n11416# a_n2157_n11546# 0.17691f
C73 a_n35_10984# a_n2157_n11546# 0.17691f
C74 a_n201_n11416# a_n2157_n11546# 0.17691f
C75 a_n201_10984# a_n2157_n11546# 0.17691f
C76 a_n367_n11416# a_n2157_n11546# 0.17691f
C77 a_n367_10984# a_n2157_n11546# 0.17691f
C78 a_n533_n11416# a_n2157_n11546# 0.17691f
C79 a_n533_10984# a_n2157_n11546# 0.17691f
C80 a_n699_n11416# a_n2157_n11546# 0.17691f
C81 a_n699_10984# a_n2157_n11546# 0.17691f
C82 a_n865_n11416# a_n2157_n11546# 0.17691f
C83 a_n865_10984# a_n2157_n11546# 0.17691f
C84 a_n1031_n11416# a_n2157_n11546# 0.17691f
C85 a_n1031_10984# a_n2157_n11546# 0.17691f
C86 a_n1197_n11416# a_n2157_n11546# 0.17691f
C87 a_n1197_10984# a_n2157_n11546# 0.17691f
C88 a_n1363_n11416# a_n2157_n11546# 0.17691f
C89 a_n1363_10984# a_n2157_n11546# 0.17691f
C90 a_n1529_n11416# a_n2157_n11546# 0.17691f
C91 a_n1529_10984# a_n2157_n11546# 0.17691f
C92 a_n1695_n11416# a_n2157_n11546# 0.17691f
C93 a_n1695_10984# a_n2157_n11546# 0.17691f
C94 a_n1861_n11416# a_n2157_n11546# 0.17691f
C95 a_n1861_10984# a_n2157_n11546# 0.17691f
C96 a_n2027_n11416# a_n2157_n11546# 0.387223f
C97 a_n2027_10984# a_n2157_n11546# 0.387223f
.ends

.subckt sky130_fd_pr__nfet_01v8_UY343Z a_n800_n138# a_n960_n224# a_n858_n50# a_800_n50#
X0 a_800_n50# a_n800_n138# a_n858_n50# a_n960_n224# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
C0 a_800_n50# a_n960_n224# 0.104672f
C1 a_n858_n50# a_n960_n224# 0.104672f
C2 a_n800_n138# a_n960_n224# 4.5759f
.ends

.subckt sky130_fd_pr__pfet_01v8_EDYT7U w_n996_n269# a_n858_n50# a_n800_n147# a_800_n50#
X0 a_800_n50# a_n800_n147# a_n858_n50# w_n996_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
C0 a_n800_n147# w_n996_n269# 2.59374f
C1 a_n800_n147# 0. 2.08416f
C2 w_n996_n269# 0. 4.35498f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_YG6WAD a_n287_n488# a_761_n400# a_819_n488# a_345_n488#
+ a_n1111_n622# a_n29_n400# a_n919_n488# a_n187_n400# a_n445_n488# a_503_n488# a_n819_n400#
+ a_n345_n400# a_n603_n488# a_661_n488# a_n977_n400# a_n761_n488# a_129_n400# a_n503_n400#
+ a_287_n400# a_n661_n400# a_919_n400# a_445_n400# a_29_n488# a_n129_n488# a_603_n400#
+ a_187_n488#
X0 a_n503_n400# a_n603_n488# a_n661_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X1 a_n29_n400# a_n129_n488# a_n187_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 a_603_n400# a_503_n488# a_445_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n819_n400# a_n919_n488# a_n977_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X4 a_n661_n400# a_n761_n488# a_n819_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X5 a_919_n400# a_819_n488# a_761_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X6 a_n187_n400# a_n287_n488# a_n345_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X7 a_761_n400# a_661_n488# a_603_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X8 a_287_n400# a_187_n488# a_129_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X9 a_n345_n400# a_n445_n488# a_n503_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X10 a_129_n400# a_29_n488# a_n29_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X11 a_445_n400# a_345_n488# a_287_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
C0 a_661_n488# a_819_n488# 0.104496f
C1 a_445_n400# a_287_n400# 0.135867f
C2 a_n761_n488# a_n919_n488# 0.104496f
C3 a_n761_n488# a_n603_n488# 0.104496f
C4 a_919_n400# a_761_n400# 0.135867f
C5 a_n187_n400# a_n29_n400# 0.135867f
C6 a_n445_n488# a_n603_n488# 0.104496f
C7 a_345_n488# a_503_n488# 0.104496f
C8 a_129_n400# a_287_n400# 0.135867f
C9 a_603_n400# a_761_n400# 0.135867f
C10 a_n819_n400# a_n661_n400# 0.135867f
C11 a_187_n488# a_29_n488# 0.104496f
C12 a_29_n488# a_n129_n488# 0.104496f
C13 a_445_n400# a_603_n400# 0.135867f
C14 a_n819_n400# a_n977_n400# 0.135867f
C15 a_n503_n400# a_n345_n400# 0.135867f
C16 a_187_n488# a_345_n488# 0.104496f
C17 a_n187_n400# a_n345_n400# 0.135867f
C18 a_n661_n400# a_n503_n400# 0.135867f
C19 a_n287_n488# a_n129_n488# 0.104496f
C20 a_129_n400# a_n29_n400# 0.135867f
C21 a_n287_n488# a_n445_n488# 0.104496f
C22 a_503_n488# a_661_n488# 0.104496f
C23 a_919_n400# a_n1111_n622# 0.255186f
C24 a_761_n400# a_n1111_n622# 0.100572f
C25 a_603_n400# a_n1111_n622# 0.100572f
C26 a_445_n400# a_n1111_n622# 0.100572f
C27 a_287_n400# a_n1111_n622# 0.100572f
C28 a_129_n400# a_n1111_n622# 0.100572f
C29 a_n29_n400# a_n1111_n622# 0.100572f
C30 a_n187_n400# a_n1111_n622# 0.100572f
C31 a_n345_n400# a_n1111_n622# 0.100572f
C32 a_n503_n400# a_n1111_n622# 0.100572f
C33 a_n661_n400# a_n1111_n622# 0.100572f
C34 a_n819_n400# a_n1111_n622# 0.100572f
C35 a_n977_n400# a_n1111_n622# 0.255186f
C36 a_819_n488# a_n1111_n622# 0.37002f
C37 a_661_n488# a_n1111_n622# 0.307217f
C38 a_503_n488# a_n1111_n622# 0.307217f
C39 a_345_n488# a_n1111_n622# 0.307217f
C40 a_187_n488# a_n1111_n622# 0.307217f
C41 a_29_n488# a_n1111_n622# 0.307217f
C42 a_n129_n488# a_n1111_n622# 0.307217f
C43 a_n287_n488# a_n1111_n622# 0.307217f
C44 a_n445_n488# a_n1111_n622# 0.307217f
C45 a_n603_n488# a_n1111_n622# 0.307217f
C46 a_n761_n488# a_n1111_n622# 0.307217f
C47 a_n919_n488# a_n1111_n622# 0.37002f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_VMUSDZ m3_n2386_n11680# m3_n2386_2480# c1_n2346_n11640#
+ m3_n2386_n6960# m3_n2386_n2240# m3_n2386_7200#
X0 c1_n2346_n11640# m3_n2386_n11680# sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X1 c1_n2346_n11640# m3_n2386_7200# sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X2 c1_n2346_n11640# m3_n2386_n2240# sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X3 c1_n2346_n11640# m3_n2386_2480# sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X4 c1_n2346_n11640# m3_n2386_n6960# sky130_fd_pr__cap_mim_m3_1 l=22 w=22
C0 c1_n2346_n11640# m3_n2386_n6960# 41.7747f
C1 m3_n2386_2480# c1_n2346_n11640# 41.7747f
C2 c1_n2346_n11640# m3_n2386_n11680# 41.6938f
C3 m3_n2386_n2240# m3_n2386_n6960# 1.03554f
C4 m3_n2386_2480# m3_n2386_n2240# 1.03554f
C5 m3_n2386_2480# m3_n2386_7200# 1.03554f
C6 c1_n2346_n11640# m3_n2386_n2240# 41.7747f
C7 c1_n2346_n11640# m3_n2386_7200# 41.696503f
C8 m3_n2386_n11680# m3_n2386_n6960# 1.03554f
C9 c1_n2346_n11640# 0. 10.3799f
C10 m3_n2386_n11680# 0. 9.126731f
C11 m3_n2386_n6960# 0. 8.37757f
C12 m3_n2386_n2240# 0. 8.37757f
C13 m3_n2386_2480# 0. 8.37757f
C14 m3_n2386_7200# 0. 9.126731f
.ends

.subckt sky130_fd_pr__nfet_01v8_HZ6WG7 a_100_n75# a_n260_n249# a_n100_n163# a_n158_n75#
X0 a_100_n75# a_n100_n163# a_n158_n75# a_n260_n249# sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=1
C0 a_100_n75# a_n260_n249# 0.118508f
C1 a_n158_n75# a_n260_n249# 0.118508f
C2 a_n100_n163# a_n260_n249# 0.720332f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_67RTNB m3_n3798_n4520# c1_n3758_n4480#
X0 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X1 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X2 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X3 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X4 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X5 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X6 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X7 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X8 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X9 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X10 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X11 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
C0 c1_n3758_n4480# m3_n3798_n4520# 0.112041p
C1 c1_n3758_n4480# 0. 10.105801f
C2 m3_n3798_n4520# 0. 29.130802f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WXTTNJ c1_n2146_n2000# m3_n2186_n2040#
X0 c1_n2146_n2000# m3_n2186_n2040# sky130_fd_pr__cap_mim_m3_1 l=20 w=20
C0 c1_n2146_n2000# m3_n2186_n2040# 34.313103f
C1 c1_n2146_n2000# 0. 2.76013f
C2 m3_n2186_n2040# 0. 8.47262f
.ends

.subckt sky130_fd_pr__diode_pd2nw_05v5_K4SERG a_n45_n45# w_n183_n183# a_n285_n285#
X0 a_n45_n45# w_n183_n183# sky130_fd_pr__diode_pd2nw_05v5 perim=1.8e+06 area=2.025e+11
C0 a_n45_n45# w_n183_n183# 0.112783f
C1 w_n183_n183# a_n285_n285# 0.690324f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_GZN5JV a_208_n400# a_366_n400# a_n558_n622# a_108_n488#
+ a_50_n400# a_n208_n488# a_266_n488# a_n366_n488# a_n108_n400# a_n266_n400# a_n50_n488#
+ a_n424_n400#
X0 a_n266_n400# a_n366_n488# a_n424_n400# a_n558_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_366_n400# a_266_n488# a_208_n400# a_n558_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2 a_50_n400# a_n50_n488# a_n108_n400# a_n558_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n108_n400# a_n208_n488# a_n266_n400# a_n558_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X4 a_208_n400# a_108_n488# a_50_n400# a_n558_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
C0 a_n424_n400# a_n266_n400# 0.135867f
C1 a_50_n400# a_n108_n400# 0.135867f
C2 a_n108_n400# a_n266_n400# 0.135867f
C3 a_208_n400# a_366_n400# 0.135867f
C4 a_50_n400# a_208_n400# 0.135867f
C5 a_366_n400# a_n558_n622# 0.255186f
C6 a_208_n400# a_n558_n622# 0.100572f
C7 a_50_n400# a_n558_n622# 0.100572f
C8 a_n108_n400# a_n558_n622# 0.100572f
C9 a_n266_n400# a_n558_n622# 0.100572f
C10 a_n424_n400# a_n558_n622# 0.255186f
C11 a_266_n488# a_n558_n622# 0.313219f
C12 a_108_n488# a_n558_n622# 0.267823f
C13 a_n50_n488# a_n558_n622# 0.267823f
C14 a_n208_n488# a_n558_n622# 0.267823f
C15 a_n366_n488# a_n558_n622# 0.313219f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_F5PPB9 c1_n1946_n7680# m3_n1986_n3800# m3_n1986_4040#
+ m3_n1986_120# m3_n1986_n7720#
X0 c1_n1946_n7680# m3_n1986_n7720# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X1 c1_n1946_n7680# m3_n1986_120# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X2 c1_n1946_n7680# m3_n1986_4040# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X3 c1_n1946_n7680# m3_n1986_n3800# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
C0 c1_n1946_n7680# m3_n1986_n3800# 28.1857f
C1 c1_n1946_n7680# m3_n1986_120# 28.1857f
C2 m3_n1986_120# m3_n1986_n3800# 0.852388f
C3 m3_n1986_4040# c1_n1946_n7680# 28.1195f
C4 m3_n1986_n7720# c1_n1946_n7680# 28.119198f
C5 m3_n1986_n7720# m3_n1986_n3800# 0.852388f
C6 m3_n1986_4040# m3_n1986_120# 0.852388f
C7 c1_n1946_n7680# 0. 7.02526f
C8 m3_n1986_n7720# 0. 6.59748f
C9 m3_n1986_n3800# 0. 5.98082f
C10 m3_n1986_120# 0. 5.98082f
C11 m3_n1986_4040# 0. 6.59748f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_E4RF2H a_2054_64# a_n2112_64# a_n1934_n961# a_898_n864#
+ a_n258_n864# a_778_n864# a_n1356_n961# a_898_64# a_n200_n961# a_n378_64# a_n956_64#
+ a_n1992_n864# a_2512_n864# a_2512_64# a_1534_n961# a_n2570_64# a_n1534_n864# a_2054_n864#
+ a_320_64# a_n1414_n864# a_956_n961# w_n2770_n1161# a_n778_n961# a_1476_64# a_778_64#
+ a_n1534_64# a_n2512_n961# a_n258_64# a_n836_64# a_378_n961# a_320_n864# a_n956_n864#
+ a_1934_n864# a_200_64# a_200_n864# a_n2570_n864# a_1476_n864# a_n836_n864# a_1934_64#
+ a_1356_64# a_n1414_64# a_2112_n961# a_n378_n864# a_n1992_64# a_1356_n864# a_n2112_n864#
X0 a_n2112_64# a_n2512_n961# a_n2570_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X1 a_n2112_n864# a_n2512_n961# a_n2570_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X2 a_n1534_n864# a_n1934_n961# a_n1992_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X3 a_200_n864# a_n200_n961# a_n258_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X4 a_1356_n864# a_956_n961# a_898_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X5 a_778_64# a_378_n961# a_320_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X6 a_n956_64# a_n1356_n961# a_n1414_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X7 a_n956_n864# a_n1356_n961# a_n1414_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X8 a_1356_64# a_956_n961# a_898_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X9 a_1934_64# a_1534_n961# a_1476_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X10 a_778_n864# a_378_n961# a_320_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X11 a_n1534_64# a_n1934_n961# a_n1992_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X12 a_200_64# a_n200_n961# a_n258_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X13 a_n378_n864# a_n778_n961# a_n836_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X14 a_2512_n864# a_2112_n961# a_2054_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X15 a_n378_64# a_n778_n961# a_n836_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X16 a_1934_n864# a_1534_n961# a_1476_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X17 a_2512_64# a_2112_n961# a_2054_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
C0 w_n2770_n1161# a_n1356_n961# 0.872004f
C1 w_n2770_n1161# a_n2570_n864# 0.171295f
C2 w_n2770_n1161# a_1534_n961# 0.872004f
C3 a_n200_n961# w_n2770_n1161# 0.872004f
C4 w_n2770_n1161# a_378_n961# 0.872004f
C5 a_n836_n864# a_n956_n864# 0.181112f
C6 a_n378_n864# a_n258_n864# 0.181112f
C7 a_1476_64# a_1356_64# 0.181112f
C8 a_n1992_64# a_n2112_64# 0.181112f
C9 w_n2770_n1161# a_n778_n961# 0.872004f
C10 w_n2770_n1161# a_2512_64# 0.171295f
C11 a_n1992_n864# a_n2112_n864# 0.181112f
C12 w_n2770_n1161# a_n1934_n961# 0.872004f
C13 a_778_64# a_898_64# 0.181112f
C14 w_n2770_n1161# a_2112_n961# 0.899231f
C15 a_n1414_n864# a_n1534_n864# 0.181112f
C16 a_778_n864# a_898_n864# 0.181112f
C17 a_n1414_64# a_n1534_64# 0.181112f
C18 a_n258_64# a_n378_64# 0.181112f
C19 w_n2770_n1161# a_n2512_n961# 0.899231f
C20 w_n2770_n1161# a_956_n961# 0.872004f
C21 w_n2770_n1161# a_n2570_64# 0.171295f
C22 a_n836_64# a_n956_64# 0.181112f
C23 a_2054_64# a_1934_64# 0.181112f
C24 a_200_64# a_320_64# 0.181112f
C25 a_1934_n864# a_2054_n864# 0.181112f
C26 w_n2770_n1161# a_2512_n864# 0.171295f
C27 a_320_n864# a_200_n864# 0.181112f
C28 a_1476_n864# a_1356_n864# 0.181112f
C29 a_2512_n864# 0. 0.136466f
C30 a_2054_n864# 0. 0.131812f
C31 a_1934_n864# 0. 0.131812f
C32 a_1476_n864# 0. 0.131812f
C33 a_1356_n864# 0. 0.131812f
C34 a_898_n864# 0. 0.131812f
C35 a_778_n864# 0. 0.131812f
C36 a_320_n864# 0. 0.131812f
C37 a_200_n864# 0. 0.131812f
C38 a_n258_n864# 0. 0.131812f
C39 a_n378_n864# 0. 0.131812f
C40 a_n836_n864# 0. 0.131812f
C41 a_n956_n864# 0. 0.131812f
C42 a_n1414_n864# 0. 0.131812f
C43 a_n1534_n864# 0. 0.131812f
C44 a_n1992_n864# 0. 0.131812f
C45 a_n2112_n864# 0. 0.131812f
C46 a_n2570_n864# 0. 0.136466f
C47 a_2512_64# 0. 0.136466f
C48 a_2054_64# 0. 0.131812f
C49 a_1934_64# 0. 0.131812f
C50 a_1476_64# 0. 0.131812f
C51 a_1356_64# 0. 0.131812f
C52 a_898_64# 0. 0.131812f
C53 a_778_64# 0. 0.131812f
C54 a_320_64# 0. 0.131812f
C55 a_200_64# 0. 0.131812f
C56 a_n258_64# 0. 0.131812f
C57 a_n378_64# 0. 0.131812f
C58 a_n836_64# 0. 0.131812f
C59 a_n956_64# 0. 0.131812f
C60 a_n1414_64# 0. 0.131812f
C61 a_n1534_64# 0. 0.131812f
C62 a_n1992_64# 0. 0.131812f
C63 a_n2112_64# 0. 0.131812f
C64 a_n2570_64# 0. 0.136466f
C65 a_2112_n961# 0. 0.879173f
C66 a_1534_n961# 0. 0.843044f
C67 a_956_n961# 0. 0.843044f
C68 a_378_n961# 0. 0.843044f
C69 a_n200_n961# 0. 0.843044f
C70 a_n778_n961# 0. 0.843044f
C71 a_n1356_n961# 0. 0.843044f
C72 a_n1934_n961# 0. 0.843044f
C73 a_n2512_n961# 0. 0.879173f
C74 w_n2770_n1161# 0. 42.723698f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_74GBJT a_n208_n497# a_266_n497# a_208_n400# a_n366_n497#
+ a_366_n400# a_n50_n497# a_50_n400# a_n108_n400# a_n266_n400# w_n624_n697# a_n424_n400#
+ a_108_n497#
X0 a_n266_n400# a_n366_n497# a_n424_n400# w_n624_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_366_n400# a_266_n497# a_208_n400# w_n624_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2 a_50_n400# a_n50_n497# a_n108_n400# w_n624_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n108_n400# a_n208_n497# a_n266_n400# w_n624_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X4 a_208_n400# a_108_n497# a_50_n400# w_n624_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
C0 a_208_n400# a_366_n400# 0.135867f
C1 a_n424_n400# w_n624_n697# 0.176254f
C2 a_208_n400# a_50_n400# 0.135867f
C3 a_n366_n497# w_n624_n697# 0.213438f
C4 a_366_n400# w_n624_n697# 0.176254f
C5 a_n266_n400# a_n108_n400# 0.135867f
C6 a_50_n400# a_n108_n400# 0.135867f
C7 a_n424_n400# a_n266_n400# 0.135867f
C8 a_n208_n497# w_n624_n697# 0.176568f
C9 a_n50_n497# w_n624_n697# 0.176568f
C10 w_n624_n697# a_266_n497# 0.213438f
C11 w_n624_n697# a_108_n497# 0.176568f
C12 a_266_n497# 0. 0.111687f
C13 a_n366_n497# 0. 0.111687f
C14 w_n624_n697# 0. 6.40384f
.ends

.subckt sky130_fd_pr__pfet_01v8_3H68VM w_n296_n619# a_n100_n497# a_100_n400# a_n158_n400#
X0 a_100_n400# a_n100_n497# a_n158_n400# w_n296_n619# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
C0 a_n158_n400# a_100_n400# 0.219309f
C1 a_100_n400# w_n296_n619# 0.268146f
C2 a_n158_n400# w_n296_n619# 0.268146f
C3 a_n100_n497# w_n296_n619# 0.434431f
C4 a_100_n400# 0. 0.211982f
C5 a_n158_n400# 0. 0.211982f
C6 a_n100_n497# 0. 0.333234f
C7 w_n296_n619# 0. 3.00565f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6RLJVT 0. a_n50_n497# a_50_n400# w_n308_n697#
+ a_n108_n400#
X0 a_50_n400# a_n50_n497# a_n108_n400# w_n308_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
C0 a_n108_n400# a_50_n400# 0.135867f
C1 a_50_n400# w_n308_n697# 0.176254f
C2 a_n108_n400# w_n308_n697# 0.176254f
C3 a_n50_n497# w_n308_n697# 0.280349f
C4 a_n50_n497# 0. 0.168405f
C5 w_n308_n697# 0. 3.39795f
.ends

.subckt sky130_fd_pr__pfet_01v8_MTZJAC 0. a_761_n400# a_n29_n400# a_n187_n400# a_n819_n400#
+ a_n345_n400# a_29_n497# a_n129_n497# a_187_n497# a_129_n400# a_n503_n400# a_n287_n497#
+ a_287_n400# a_n661_n400# a_345_n497# a_n445_n497# a_445_n400# a_503_n497# a_n603_n497#
+ a_661_n497# w_n957_n619# a_603_n400# a_n761_n497#
X0 a_n661_n400# a_n761_n497# a_n819_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_n187_n400# a_n287_n497# a_n345_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 a_761_n400# a_661_n497# a_603_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X3 a_287_n400# a_187_n497# a_129_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X4 a_n345_n400# a_n445_n497# a_n503_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X5 a_129_n400# a_29_n497# a_n29_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X6 a_445_n400# a_345_n497# a_287_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X7 a_n503_n400# a_n603_n497# a_n661_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X8 a_n29_n400# a_n129_n497# a_n187_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X9 a_603_n400# a_503_n497# a_445_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
C0 a_n819_n400# a_n661_n400# 0.135867f
C1 a_287_n400# a_129_n400# 0.135867f
C2 a_n661_n400# a_n503_n400# 0.135867f
C3 a_187_n497# w_n957_n619# 0.183383f
C4 a_n29_n400# a_n187_n400# 0.135867f
C5 a_603_n400# a_445_n400# 0.135867f
C6 a_n445_n497# w_n957_n619# 0.183435f
C7 w_n957_n619# a_761_n400# 0.206529f
C8 a_n29_n400# a_129_n400# 0.135867f
C9 a_n603_n497# w_n957_n619# 0.183581f
C10 a_n761_n497# w_n957_n619# 0.218643f
C11 a_n345_n400# a_n187_n400# 0.135867f
C12 a_29_n497# w_n957_n619# 0.183364f
C13 a_n287_n497# w_n957_n619# 0.183383f
C14 a_n129_n497# w_n957_n619# 0.183364f
C15 a_603_n400# a_761_n400# 0.135867f
C16 a_503_n497# w_n957_n619# 0.183581f
C17 a_661_n497# w_n957_n619# 0.218643f
C18 a_345_n497# w_n957_n619# 0.183435f
C19 a_n819_n400# w_n957_n619# 0.206529f
C20 a_n345_n400# a_n503_n400# 0.135867f
C21 a_287_n400# a_445_n400# 0.135867f
C22 a_661_n497# 0. 0.120549f
C23 a_503_n497# 0. 0.105254f
C24 a_345_n497# 0. 0.105254f
C25 a_187_n497# 0. 0.105254f
C26 a_29_n497# 0. 0.105254f
C27 a_n129_n497# 0. 0.105254f
C28 a_n287_n497# 0. 0.105254f
C29 a_n445_n497# 0. 0.105254f
C30 a_n603_n497# 0. 0.105254f
C31 a_n761_n497# 0. 0.120549f
C32 w_n957_n619# 0. 8.63602f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_Z6W9J4 a_2223_n200# a_n1703_n200# a_1245_n288#
+ a_n1245_n200# a_n1125_n200# a_667_n288# a_n489_n288# a_n2223_n288# a_1765_n200#
+ a_n667_n200# a_89_n288# a_1645_n200# a_31_n200# a_n2281_n200# a_1187_n200# a_n547_n200#
+ a_1067_n200# a_n89_n200# a_n1645_n288# a_609_n200# a_489_n200# a_1823_n288# a_n1067_n288#
+ a_n1823_n200# a_n2415_n422#
X0 a_n89_n200# a_n489_n288# a_n547_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X1 a_1645_n200# a_1245_n288# a_1187_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X2 a_n1823_n200# a_n2223_n288# a_n2281_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X3 a_n1245_n200# a_n1645_n288# a_n1703_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X4 a_489_n200# a_89_n288# a_31_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X5 a_1067_n200# a_667_n288# a_609_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X6 a_n667_n200# a_n1067_n288# a_n1125_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X7 a_2223_n200# a_1823_n288# a_1765_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
C0 a_2223_n200# a_n2415_n422# 0.162747f
C1 a_n2281_n200# a_n2415_n422# 0.162747f
C2 a_1823_n288# a_n2415_n422# 1.20369f
C3 a_1245_n288# a_n2415_n422# 1.16396f
C4 a_667_n288# a_n2415_n422# 1.16396f
C5 a_89_n288# a_n2415_n422# 1.16396f
C6 a_n489_n288# a_n2415_n422# 1.16396f
C7 a_n1067_n288# a_n2415_n422# 1.16396f
C8 a_n1645_n288# a_n2415_n422# 1.16396f
C9 a_n2223_n288# a_n2415_n422# 1.20369f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_8CDM6Z a_n887_n497# a_n29_n400# w_n1145_n697#
+ a_887_n400# a_n429_n497# a_487_n497# a_429_n400# a_29_n497# a_n945_n400# a_n487_n400#
X0 a_n487_n400# a_n887_n497# a_n945_n400# w_n1145_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=2
X1 a_n29_n400# a_n429_n497# a_n487_n400# w_n1145_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X2 a_429_n400# a_29_n497# a_n29_n400# w_n1145_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X3 a_887_n400# a_487_n497# a_429_n400# w_n1145_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=2
C0 w_n1145_n697# a_n429_n497# 0.574033f
C1 w_n1145_n697# a_487_n497# 0.610903f
C2 w_n1145_n697# a_887_n400# 0.176229f
C3 w_n1145_n697# a_n887_n497# 0.610903f
C4 w_n1145_n697# a_n945_n400# 0.176229f
C5 a_29_n497# w_n1145_n697# 0.574033f
C6 a_887_n400# 0. 0.136466f
C7 a_429_n400# 0. 0.201699f
C8 a_n29_n400# 0. 0.201699f
C9 a_n487_n400# 0. 0.201699f
C10 a_n945_n400# 0. 0.136466f
C11 a_487_n497# 0. 0.451792f
C12 a_29_n497# 0. 0.439839f
C13 a_n429_n497# 0. 0.439839f
C14 a_n887_n497# 0. 0.451792f
C15 w_n1145_n697# 0. 11.293f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_UYSCL3 c1_n1852_n1560# m3_n1892_120# m3_n150_130#
+ c1_n110_n1550# m3_n150_n1590# m3_n1892_n1600#
X0 c1_n110_n1550# m3_n150_n1590# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1 c1_n1852_n1560# m3_n1892_120# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X2 c1_n1852_n1560# m3_n1892_n1600# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X3 c1_n110_n1550# m3_n150_130# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
C0 c1_n110_n1550# m3_n150_n1590# 4.5192f
C1 c1_n110_n1550# m3_n150_130# 4.5192f
C2 m3_n150_130# m3_n150_n1590# 0.343637f
C3 c1_n110_n1550# c1_n1852_n1560# 0.465192f
C4 m3_n1892_n1600# m3_n150_n1590# 0.335741f
C5 m3_n150_130# m3_n1892_120# 0.335741f
C6 c1_n1852_n1560# m3_n1892_120# 4.53819f
C7 m3_n1892_n1600# m3_n1892_120# 0.346413f
C8 m3_n1892_n1600# c1_n1852_n1560# 4.53819f
C9 c1_n110_n1550# 0. 1.21594f
C10 c1_n1852_n1560# 0. 1.21725f
C11 m3_n150_n1590# 0. 1.40223f
C12 m3_n1892_n1600# 0. 1.41064f
C13 m3_n150_130# 0. 1.40223f
C14 m3_n1892_120# 0. 1.41064f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_43FTN9 m3_n3546_n7996# c1_n3506_n7956#
X0 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X1 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X2 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X3 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X4 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X5 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X6 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X7 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X8 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X9 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X10 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X11 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X12 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X13 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X14 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X15 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X16 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X17 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X18 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X19 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X20 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
C0 c1_n3506_n7956# m3_n3546_n7996# 0.19948p
C1 c1_n3506_n7956# 0. 14.9827f
C2 m3_n3546_n7996# 0. 48.056602f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_3DMTNZ m3_n2492_120# m3_n134_n2252# m3_n136_122#
+ c1_n2452_160# m3_n2490_n2254#
X0 c1_n2452_160# m3_n2492_120# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X1 c1_n2452_160# m3_n2490_n2254# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X2 c1_n2452_160# m3_n134_n2252# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X3 c1_n2452_160# m3_n136_122# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
C0 m3_n136_122# m3_n134_n2252# 0.411947f
C1 c1_n2452_160# m3_n134_n2252# 9.11198f
C2 m3_n2490_n2254# m3_n134_n2252# 0.431944f
C3 m3_n136_122# m3_n2492_120# 0.431944f
C4 c1_n2452_160# m3_n2492_120# 9.09961f
C5 m3_n2490_n2254# m3_n2492_120# 0.411155f
C6 c1_n2452_160# m3_n136_122# 9.10957f
C7 m3_n2490_n2254# c1_n2452_160# 9.102059f
C8 c1_n2452_160# 0. 3.76699f
C9 m3_n134_n2252# 0. 2.37869f
C10 m3_n2490_n2254# 0. 2.37512f
C11 m3_n136_122# 0. 2.37869f
C12 m3_n2492_120# 0. 2.37512f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_4HHTN9 0. m3_n1186_n4520# c1_n1146_n4480#
X0 c1_n1146_n4480# m3_n1186_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X1 c1_n1146_n4480# m3_n1186_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X2 c1_n1146_n4480# m3_n1186_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X3 c1_n1146_n4480# m3_n1186_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
C0 c1_n1146_n4480# m3_n1186_n4520# 36.4513f
C1 c1_n1146_n4480# 0. 4.0756f
C2 m3_n1186_n4520# 0. 10.3653f
.ends

.subckt sky130_fd_pr__pfet_01v8_M6QFHF a_229_n164# a_229_64# a_n287_64# a_n29_64#
+ a_29_n261# a_n29_n164# a_n229_n261# w_n425_n383# a_n287_n164#
X0 a_n29_64# a_n229_n261# a_n287_64# w_n425_n383# sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X1 a_n29_n164# a_n229_n261# a_n287_n164# w_n425_n383# sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X2 a_229_n164# a_29_n261# a_n29_n164# w_n425_n383# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X3 a_229_64# a_29_n261# a_n29_64# w_n425_n383# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
C0 a_n229_n261# w_n425_n383# 0.508421f
C1 a_29_n261# w_n425_n383# 0.508421f
C2 a_29_n261# a_n229_n261# 0.164962f
C3 a_29_n261# 0. 0.412709f
C4 a_n229_n261# 0. 0.412709f
C5 w_n425_n383# 0. 2.68504f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_H6M2KM a_n2516_n42# a_2458_n42# a_800_n42# a_858_n130#
+ a_n2650_n264# a_n800_n130# a_n2458_n130#
X0 a_800_n42# a_n800_n130# a_n858_n42# a_n2650_n264# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X1 a_n858_n42# a_n2458_n130# a_n2516_n42# a_n2650_n264# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X2 a_2458_n42# a_858_n130# a_800_n42# a_n2650_n264# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
C0 a_n800_n130# a_858_n130# 0.104496f
C1 a_n800_n130# a_n2458_n130# 0.104496f
C2 a_858_n130# a_n2650_n264# 4.24097f
C3 a_n800_n130# a_n2650_n264# 4.17816f
C4 a_n2458_n130# a_n2650_n264# 4.24097f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_BKL7UB a_n1414_n855# a_n1548_n1077# a_778_55#
+ a_n836_55# a_n258_55# a_n1356_n943# a_n200_n943# a_320_n855# a_n956_n855# a_200_55#
+ a_200_n855# a_n836_n855# a_n1414_55# a_1356_55# a_n378_n855# a_1356_n855# a_956_n943#
+ a_n778_n943# a_898_n855# a_n258_n855# a_778_n855# a_378_n943# a_898_55# a_n956_55#
+ a_n378_55# a_320_55#
X0 a_n956_55# a_n1356_n943# a_n1414_55# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X1 a_n956_n855# a_n1356_n943# a_n1414_n855# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X2 a_1356_55# a_956_n943# a_898_55# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X3 a_778_n855# a_378_n943# a_320_n855# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X4 a_200_55# a_n200_n943# a_n258_55# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X5 a_n378_n855# a_n778_n943# a_n836_n855# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X6 a_n378_55# a_n778_n943# a_n836_55# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X7 a_200_n855# a_n200_n943# a_n258_n855# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X8 a_1356_n855# a_956_n943# a_898_n855# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X9 a_778_55# a_378_n943# a_320_55# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
C0 a_n836_55# a_n956_55# 0.181112f
C1 a_n258_55# a_n378_55# 0.181112f
C2 a_320_n855# a_200_n855# 0.181112f
C3 a_320_55# a_200_55# 0.181112f
C4 a_n378_n855# a_n258_n855# 0.181112f
C5 a_n836_n855# a_n956_n855# 0.181112f
C6 a_898_n855# a_778_n855# 0.181112f
C7 a_778_55# a_898_55# 0.181112f
C8 a_1356_n855# a_n1548_n1077# 0.307524f
C9 a_898_n855# a_n1548_n1077# 0.141567f
C10 a_778_n855# a_n1548_n1077# 0.141567f
C11 a_320_n855# a_n1548_n1077# 0.141567f
C12 a_200_n855# a_n1548_n1077# 0.141567f
C13 a_n258_n855# a_n1548_n1077# 0.141567f
C14 a_n378_n855# a_n1548_n1077# 0.141567f
C15 a_n836_n855# a_n1548_n1077# 0.141567f
C16 a_n956_n855# a_n1548_n1077# 0.141567f
C17 a_n1414_n855# a_n1548_n1077# 0.307524f
C18 a_1356_55# a_n1548_n1077# 0.307524f
C19 a_898_55# a_n1548_n1077# 0.141567f
C20 a_778_55# a_n1548_n1077# 0.141567f
C21 a_320_55# a_n1548_n1077# 0.141567f
C22 a_200_55# a_n1548_n1077# 0.141567f
C23 a_n258_55# a_n1548_n1077# 0.141567f
C24 a_n378_55# a_n1548_n1077# 0.141567f
C25 a_n836_55# a_n1548_n1077# 0.141567f
C26 a_n956_55# a_n1548_n1077# 0.141567f
C27 a_n1414_55# a_n1548_n1077# 0.307524f
C28 a_956_n943# a_n1548_n1077# 1.72027f
C29 a_378_n943# a_n1548_n1077# 1.66049f
C30 a_n200_n943# a_n1548_n1077# 1.66049f
C31 a_n778_n943# a_n1548_n1077# 1.66049f
C32 a_n1356_n943# a_n1548_n1077# 1.72027f
.ends

.subckt sky130_fd_pr__nfet_01v8_Y7GPAW a_n287_n488# a_761_n400# a_345_n488# a_n29_n400#
+ a_n187_n400# a_n445_n488# a_503_n488# a_n819_n400# a_n345_n400# a_n603_n488# a_661_n488#
+ a_n761_n488# a_129_n400# a_n503_n400# a_287_n400# a_n661_n400# a_n921_n574# a_445_n400#
+ a_29_n488# a_n129_n488# a_603_n400# a_187_n488#
X0 a_n503_n400# a_n603_n488# a_n661_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X1 a_n29_n400# a_n129_n488# a_n187_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 a_603_n400# a_503_n488# a_445_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n661_n400# a_n761_n488# a_n819_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X4 a_n187_n400# a_n287_n488# a_n345_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X5 a_761_n400# a_661_n488# a_603_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X6 a_287_n400# a_187_n488# a_129_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X7 a_n345_n400# a_n445_n488# a_n503_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X8 a_129_n400# a_29_n488# a_n29_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X9 a_445_n400# a_345_n488# a_287_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
C0 a_n345_n400# a_n187_n400# 0.135867f
C1 a_445_n400# a_603_n400# 0.135867f
C2 a_129_n400# a_287_n400# 0.135867f
C3 a_n29_n400# a_n187_n400# 0.135867f
C4 a_n503_n400# a_n345_n400# 0.135867f
C5 a_445_n400# a_287_n400# 0.135867f
C6 a_n661_n400# a_n503_n400# 0.135867f
C7 a_129_n400# a_n29_n400# 0.135867f
C8 a_n819_n400# a_n661_n400# 0.135867f
C9 a_603_n400# a_761_n400# 0.135867f
C10 a_761_n400# a_n921_n574# 0.279003f
C11 a_603_n400# a_n921_n574# 0.101564f
C12 a_445_n400# a_n921_n574# 0.101564f
C13 a_287_n400# a_n921_n574# 0.101564f
C14 a_129_n400# a_n921_n574# 0.101564f
C15 a_n29_n400# a_n921_n574# 0.101564f
C16 a_n187_n400# a_n921_n574# 0.101564f
C17 a_n345_n400# a_n921_n574# 0.101564f
C18 a_n503_n400# a_n921_n574# 0.101564f
C19 a_n661_n400# a_n921_n574# 0.101564f
C20 a_n819_n400# a_n921_n574# 0.279003f
C21 a_661_n488# a_n921_n574# 0.32743f
C22 a_503_n488# a_n921_n574# 0.280464f
C23 a_345_n488# a_n921_n574# 0.280318f
C24 a_187_n488# a_n921_n574# 0.280266f
C25 a_29_n488# a_n921_n574# 0.280247f
C26 a_n129_n488# a_n921_n574# 0.280247f
C27 a_n287_n488# a_n921_n574# 0.280266f
C28 a_n445_n488# a_n921_n574# 0.280318f
C29 a_n603_n488# a_n921_n574# 0.280464f
C30 a_n761_n488# a_n921_n574# 0.32743f
.ends

.subckt sky130_fd_pr__pfet_01v8_LL48TN a_n1802_n464# a_86_n561# a_2202_n464# a_1744_64#
+ a_n1802_64# a_486_64# a_n544_n464# a_n1116_n464# a_n544_64# a_658_n561# a_600_n464#
+ a_1172_64# a_n86_64# a_n1230_64# a_1630_n464# a_n1688_n464# a_28_64# a_1172_n464#
+ a_n86_n464# a_n2202_n561# a_n1688_64# a_1058_64# a_n1116_64# a_n658_n464# a_1744_n464#
+ a_486_n464# a_n1630_n561# w_n2398_n683# a_1630_64# a_1058_n464# a_n2260_n464# a_28_n464#
+ a_n658_64# a_1230_n561# a_n1230_n464# a_n1058_n561# a_n486_n561# a_600_64# a_2202_64#
+ a_1802_n561# a_n2260_64#
X0 a_1058_64# a_658_n561# a_600_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X1 a_2202_64# a_1802_n561# a_1744_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X2 a_n1802_n464# a_n2202_n561# a_n2260_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X3 a_486_n464# a_86_n561# a_28_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X4 a_1630_64# a_1230_n561# a_1172_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X5 a_486_64# a_86_n561# a_28_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X6 a_n1802_64# a_n2202_n561# a_n2260_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X7 a_1058_n464# a_658_n561# a_600_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X8 a_2202_n464# a_1802_n561# a_1744_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X9 a_n1230_n464# a_n1630_n561# a_n1688_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X10 a_1630_n464# a_1230_n561# a_1172_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X11 a_n86_64# a_n486_n561# a_n544_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X12 a_n658_n464# a_n1058_n561# a_n1116_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X13 a_n86_n464# a_n486_n561# a_n544_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X14 a_n1230_64# a_n1630_n561# a_n1688_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X15 a_n658_64# a_n1058_n561# a_n1116_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
C0 w_n2398_n683# a_n1630_n561# 0.893055f
C1 w_n2398_n683# a_1230_n561# 0.893055f
C2 w_n2398_n683# a_2202_n464# 0.106719f
C3 w_n2398_n683# a_2202_64# 0.106719f
C4 w_n2398_n683# a_n2202_n561# 0.917079f
C5 w_n2398_n683# a_n2260_n464# 0.106719f
C6 w_n2398_n683# a_1802_n561# 0.917079f
C7 w_n2398_n683# a_658_n561# 0.892931f
C8 w_n2398_n683# a_n486_n561# 0.892875f
C9 w_n2398_n683# a_n1058_n561# 0.892931f
C10 w_n2398_n683# a_n2260_64# 0.106719f
C11 w_n2398_n683# a_86_n561# 0.892875f
C12 a_1802_n561# 0. 0.875166f
C13 a_1230_n561# 0. 0.831559f
C14 a_658_n561# 0. 0.831559f
C15 a_86_n561# 0. 0.831559f
C16 a_n486_n561# 0. 0.831559f
C17 a_n1058_n561# 0. 0.831559f
C18 a_n1630_n561# 0. 0.831559f
C19 a_n2202_n561# 0. 0.875166f
C20 w_n2398_n683# 0. 22.788599f
.ends

.subckt sky130_be_ip__lsxo avdd avss dvdd dvss ibias ena standby dout xout xin
Xamp_XR1 m1_24220_n8834# m1_24220_n8502# m1_10618_n7674# m1_10620_n9664# m1_10620_n8670#
+ m1_10620_n8006# m1_24220_n7840# m1_10620_n9334# m1_24220_n9166# m1_24220_n8172#
+ inv_in m1_24220_n9166# li_9150_n9268# m1_10620_n8338# m1_24220_n9832# m1_10620_n8670#
+ m1_10620_n9664# m1_24220_n9500# m1_24220_n8502# m1_24220_n9500# m1_10620_n9002#
+ m1_10620_n9334# m1_24220_n8834# m1_10620_n8006# m1_10618_n7674# m1_10620_n8338#
+ m1_24220_n8172# dvss_ip m1_10620_n9002# m1_24220_n7840# m1_24220_n9832# sky130_fd_pr__res_xhigh_po_0p35_WHP78W
Xbias_XR2 m1_2130_n17240# m1_18932_n16742# m1_2130_n16908# m1_2132_n15912# m1_18932_n17406#
+ m1_18932_n15746# vg2 m1_2132_n14254# m1_18932_n17074# m1_18932_n15746# m1_2132_n15248#
+ m1_18932_n14418# m1_18932_n17074# m1_2132_n16576# m1_2132_n17570# m1_2130_n16908#
+ avss_ip m1_2132_n14916# avss_ip m1_18932_n17738# m1_18932_n16078# m1_2134_n14584#
+ m1_2130_n15578# m1_2130_n17240# m1_2132_n16242# m1_18932_n15414# m1_18932_n17406#
+ m1_18932_n14750# avss_ip m1_18932_n16410# m1_2132_n14916# m1_18932_n15414# m1_2132_n17904#
+ m1_18932_n15082# m1_2132_n16242# m1_18932_n16410# vg1 m1_2132_n14254# m1_2132_n17570#
+ m1_2132_n15248# m1_2132_n16576# avss_ip m1_2132_n17904# m1_18932_n17738# m1_18932_n16078#
+ m1_18932_n14418# m1_2134_n14584# avss_ip m1_18932_n16742# m1_2132_n15912# m1_18932_n15082#
+ m1_2130_n15578# m1_18932_n14750# sky130_fd_pr__res_xhigh_po_0p35_M35ED8
Xx1 ena dvss dvss dvdd dvdd ena_ip sky130_fd_sc_hd__buf_1
Xbias_XR3 avss_ip avss_ip m1_3134_n13314# avss_ip avss_ip vrb avss_ip m1_3134_n13314#
+ avss_ip sky130_fd_pr__res_xhigh_po_0p35_VTNT3C
Xesd_n_xout avss_ip xout sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
Xant_diode_standby dvss standby sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
Xx2 standby dvss dvss dvdd dvdd standby_ip sky130_fd_sc_hd__buf_1
Xamp_XM4_18 dvss_ip xin_buf xin_buf vn dvss_ip vn vn vn vn vn sky130_fd_pr__nfet_01v8_LHQHT5
Xx3 dvdd dvss ena_ip x3/in_b x3/out_b x3/out avdd avss avdd level_shift
Xx4 dvdd dvss standby_ip standby_b x4/out_b standby_33 avdd avss avdd level_shift
Xesd_n_xin avss_ip xin sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
Xamp_XM11_13 dvss_ip inv_m2 inv_m2 dvss_ip inv_m1 dout_ip dout_ip dvss_ip dvss_ip
+ sky130_fd_pr__nfet_01v8_6G4XAN
Xx7 dout_ip standby_ip x7/x1/x2/a_27_47# x7/x2/x2/a_27_47# x7/x1/x3/a_27_47# x7/x2/x3/a_27_47#
+ x7/x2/Qb1 x7/x1/Qb1 x7/x1/x4/a_27_47# x7/x2/x4/a_27_47# x7/x2/Qb2 x7/ena_done_b
+ x7/stby_done_b x7/clk_disable dout_filt ena_ip x7/x1/Qb2 dvss dvdd standby_b x7/x1/x2/a_193_47#
+ ripl_dly_clk_buf
Xbias_XM5 icnode avss_ip avss_ip vg2 sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXR2 m1_2130_n21506# m1_24530_n21008# m1_2130_n20510# m1_24528_n22338# m1_2130_n20510#
+ m1_2130_n19514# m1_24530_n19348# m1_2128_n22170# m1_2128_n21174# m1_24530_n21672#
+ m1_2130_n20842# m1_24530_n20012# m1_24530_n20676# m1_2130_n20180# avss_ip m1_24528_n21342#
+ avss_ip m1_2128_n21174# avss_ip m1_2130_n19846# m1_2130_n18850# m1_24530_n19016#
+ xin m1_2130_n21838# m1_2130_n21506# m1_24530_n21008# m1_24528_n22004# m1_24530_n19680#
+ m1_24528_n21342# m1_2130_n19184# m1_2130_n19514# m1_24530_n19348# m1_2128_n22170#
+ m1_24530_n19016# m1_24530_n20344# m1_2130_n20180# m1_24530_n20676# m1_2130_n19184#
+ avss_ip m1_2130_n20842# m1_2130_n21838# m1_2130_n19846# m1_24530_n19680# m1_24528_n22338#
+ m1_2130_n18850# m1_24530_n21672# m1_24530_n20344# avss_ip m1_24530_n20012# xout
+ m1_24528_n22004# sky130_fd_pr__res_xhigh_po_0p35_68VL2P
Xamp_XM7 inv_in dvss_ip inv_m1 dvss_ip sky130_fd_pr__nfet_01v8_UY343Z
Xamp_XM6 dvdd_ip inv_m1 inv_in dvdd_ip sky130_fd_pr__pfet_01v8_EDYT7U
Xamp_XM8 dvdd_ip dvdd_ip li_9150_n9268# li_9150_n9268# sky130_fd_pr__pfet_01v8_EDYT7U
XXM1 xin avss_ip xin xin avss_ip xout xin avss_ip xin xin avss_ip xout xin xin avss_ip
+ xin avss_ip avss_ip xout xout avss_ip avss_ip xin xin xout xin sky130_fd_pr__nfet_g5v0d10v5_YG6WAD
Xamp_XM9 li_9150_n9268# dvss_ip li_9150_n9268# dvss_ip sky130_fd_pr__nfet_01v8_UY343Z
XXM3 dvss standby_ip dvss dout_ip sky130_fd_pr__nfet_01v8_AHZR5K
Xbias_XC1 xin xin vg1 xin xin xin sky130_fd_pr__cap_mim_m3_1_VMUSDZ
XXM4 dout dvss_ip dout_filt dvss_ip sky130_fd_pr__nfet_01v8_HZ6WG7
Xamp_XC1 xin_buf inv_in sky130_fd_pr__cap_mim_m3_1_67RTNB
Xbias_XC2 avdd_ip icnode sky130_fd_pr__cap_mim_m3_1_WXTTNJ
Xesd_p_xout xout avdd_ip avss_ip sky130_fd_pr__diode_pd2nw_05v5_K4SERG
XXM5 avss_ip avss avss x3/out avss x3/out x3/out x3/out avss_ip avss x3/out avss_ip
+ sky130_fd_pr__nfet_g5v0d10v5_GZN5JV
Xbias_XC3 avss_ip vg2 vg2 vg2 vg2 sky130_fd_pr__cap_mim_m3_1_F5PPB9
XXM2_bias_XM3_4 avdd_ip avdd_ip vbreg avdd_ip li_22598_n15512# avdd_ip vbreg avdd_ip
+ vbreg xout avdd_ip avdd_ip avdd_ip avdd_ip vbreg avdd_ip xout avdd_ip xout xout
+ vbreg avdd_ip vbreg xout avdd_ip xout vbreg xout avdd_ip vbreg vbreg avdd_ip avdd_ip
+ xout li_22598_n15512# avdd_ip xout avdd_ip avdd_ip xout xout vbreg vg1 avdd_ip xout
+ avdd_ip sky130_fd_pr__pfet_g5v0d10v5_E4RF2H
Xant_diode_ena dvss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
XXM6 x3/out_b x3/out_b avdd_ip x3/out_b avdd x3/out_b avdd avdd_ip avdd avdd avdd_ip
+ x3/out_b sky130_fd_pr__pfet_g5v0d10v5_74GBJT
XXM7 dvdd_ip dout_filt dout dvdd_ip sky130_fd_pr__pfet_01v8_3H68VM
XXM9 dvss standby_33 ibias ibias ibias_ip sky130_fd_pr__pfet_g5v0d10v5_6RLJVT
XXM8 dvss dvdd dvdd_ip dvdd dvdd dvdd_ip standby_ip standby_ip standby_ip dvdd dvdd
+ standby_ip dvdd_ip dvdd_ip standby_ip standby_ip dvdd standby_ip standby_ip standby_ip
+ dvdd dvdd_ip standby_ip sky130_fd_pr__pfet_01v8_MTZJAC
Xamp_XM1_2 dvss_ip dvss_ip ibias_ip ibias_ip ibias_ip ibias_ip ibias_ip ibias_ip dvss_ip
+ dvss_ip ibias_ip dvss_ip vbp dvss_ip ibias_ip dvss_ip ibias_ip ibias_ip ibias_ip
+ dvss_ip dvss_ip ibias_ip ibias_ip dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5_Z6W9J4
Xamp_XM3_5 xin tail dvdd_ip xin_buf xin xout xin_buf xout vn vn sky130_fd_pr__pfet_g5v0d10v5_8CDM6Z
Xesd_p_xin xin avdd_ip avss_ip sky130_fd_pr__diode_pd2nw_05v5_K4SERG
XXC1 avdd_ip avss_ip avss_ip avdd_ip avss_ip avss_ip sky130_fd_pr__cap_mim_m3_1_UYSCL3
XXC2 dvss_ip dvdd_ip sky130_fd_pr__cap_mim_m3_1_43FTN9
XXC3 avdd avdd avdd avss avdd sky130_fd_pr__cap_mim_m3_1_3DMTNZ
XXC4 dvss dvss dvdd sky130_fd_pr__cap_mim_m3_1_4HHTN9
Xamp_XM10_12 dout_ip dout_ip inv_m2 dvdd_ip inv_m2 dvdd_ip inv_m1 dvdd_ip dvdd_ip
+ sky130_fd_pr__pfet_01v8_M6QFHF
Xbias_XM6_7_8 vbreg avss_ip li_8336_n12442# li_8336_n12442# avss_ip icnode icnode
+ sky130_fd_pr__nfet_g5v0d10v5_H6M2KM
Xbias_XM1_2 avss_ip avss_ip vrb vrb avss_ip avss_ip vg1 vbreg avss_ip vg1 vbreg vrb
+ avss_ip avss_ip vbreg avss_ip avss_ip vg2 avss_ip vbreg vrb vg2 avss_ip avss_ip
+ vbreg vbreg sky130_fd_pr__nfet_g5v0d10v5_BKL7UB
XXM11 standby_b dvss standby_b dvss_ip dvss standby_b standby_b dvss dvss_ip standby_b
+ standby_b standby_b dvss dvss dvss_ip dvss_ip dvss dvss standby_b standby_b dvss_ip
+ standby_b sky130_fd_pr__nfet_01v8_Y7GPAW
Xamp_XM16_17 dvdd_ip vbp dvdd_ip dvdd_ip dvdd_ip dvdd_ip dvdd_ip tail dvdd_ip vbp
+ dvdd_ip tail dvdd_ip tail dvdd_ip dvdd_ip vbp tail tail vbp dvdd_ip tail tail dvdd_ip
+ dvdd_ip dvdd_ip vbp dvdd_ip dvdd_ip tail dvdd_ip tail dvdd_ip vbp tail vbp vbp dvdd_ip
+ dvdd_ip vbp dvdd_ip sky130_fd_pr__pfet_01v8_LL48TN
C0 xin_buf m1_10620_n8670# 0.16582f
C1 inv_in vbp 0.265485f
C2 dvdd_ip dvss 5.10936f
C3 m1_2130_n18850# avss_ip 0.215196f
C4 vg1 xout 0.631204f
C5 dvss_ip li_9150_n9268# 6.801351f
C6 dvss_ip m1_10620_n9664# 0.148031f
C7 dvdd_ip dvss_ip 0.303008p
C8 avss_ip m1_18932_n14418# 0.105925f
C9 standby_33 dvss 0.577404f
C10 m1_2132_n15912# avss_ip 0.185425f
C11 vrb dvdd_ip 0.182588f
C12 xin_buf dout_ip 0.1539f
C13 avdd_ip x3/out_b 2.337762f
C14 dvss_ip standby_33 3.432307f
C15 avss_ip m1_24528_n22004# 0.141047f
C16 dvss_ip m1_24220_n8172# 0.366376f
C17 inv_in m1_24220_n7840# 0.127215f
C18 dvdd dout_filt 1.583258f
C19 dvdd x7/x2/Qb1 0.384866f
C20 vg2 m1_2130_n15578# 0.156683f
C21 ena_ip dvss 4.924581f
C22 dvss_ip m1_18932_n14418# 0.117297f
C23 m1_10618_n7674# dvdd_ip 0.100908f
C24 dvdd_ip vg2 0.10449f
C25 xin_buf li_9150_n9268# 1.093907f
C26 ena dvss 0.278448f
C27 xin_buf m1_10620_n9664# 0.140848f
C28 xin_buf dvdd_ip 19.03397f
C29 avdd_ip dvdd_ip 3.929127f
C30 m1_24530_n21672# avss_ip 0.148711f
C31 dvdd_ip tail 2.861027f
C32 m1_24530_n19680# xin 0.159253f
C33 dvss_ip avss_ip 24.136833f
C34 vn dvss_ip 5.211006f
C35 standby_b standby_33 0.114197f
C36 xin_buf standby_33 2.348183f
C37 x3/out_b x3/out 0.53847f
C38 m1_2130_n21838# avss_ip 0.188571f
C39 vrb avss_ip 5.123528f
C40 m1_18932_n14750# avss_ip 0.133139f
C41 dvss_ip dvss 16.725235f
C42 m1_24220_n9832# dvss_ip 0.48684f
C43 vg2 m1_18932_n14418# 0.272043f
C44 m1_2130_n20510# xin 0.164971f
C45 x3/out_b avss 0.468413f
C46 vg2 m1_2132_n15912# 0.154604f
C47 inv_in dvdd_ip 7.786261f
C48 ena_ip standby_b 3.082387f
C49 m1_18932_n15746# avss_ip 0.19127f
C50 vg2 avss_ip 42.440594f
C51 xin_buf avss_ip 10.849238f
C52 xin_buf vn 4.728283f
C53 vrb dvss_ip 1.203343f
C54 dvss_ip m1_18932_n14750# 0.144339f
C55 vbreg xin 0.157652f
C56 avdd_ip avss_ip 0.825243p
C57 m1_2130_n20180# xin 0.1652f
C58 m1_24530_n19016# avss_ip 0.141729f
C59 vn tail 0.624406f
C60 standby_b dvss 13.115542f
C61 xin_buf dvss 0.918436f
C62 vbreg li_22598_n15512# 2.192764f
C63 dvdd_ip vg1 0.707385f
C64 m1_10618_n7674# dvss_ip 0.16974f
C65 dvss_ip m1_18932_n15746# 0.124217f
C66 dvss_ip m1_10620_n8338# 0.157268f
C67 dvss_ip vg2 3.927598f
C68 avss_ip m1_18932_n16742# 0.406957f
C69 standby_b dvss_ip 3.570977f
C70 xin_buf dvss_ip 27.769085f
C71 dvss_ip m1_24220_n9500# 0.367115f
C72 standby_33 avss 0.151707f
C73 avdd_ip dvss_ip 20.912617f
C74 vrb vg2 4.613826f
C75 dvss_ip tail 0.416371f
C76 inv_in avss_ip 1.948904f
C77 vn inv_in 0.137437f
C78 icnode li_8336_n12442# 1.350289f
C79 avss_ip x3/out 2.407235f
C80 m1_2128_n22170# avss_ip 0.191378f
C81 inv_in dvss 0.100479f
C82 dvss_ip m1_18932_n16742# 0.11359f
C83 ena_ip avss 0.318302f
C84 avss_ip avss 6.445405f
C85 dvdd dout 0.550876f
C86 standby_ip ibias 0.288754f
C87 m1_10618_n7674# xin_buf 0.173169f
C88 xin_buf m1_10620_n8338# 0.166314f
C89 xin_buf vg2 3.568495f
C90 inv_in dvss_ip 13.663485f
C91 avdd_ip vg2 0.280688f
C92 xin_buf avdd_ip 9.058875f
C93 dvdd x7/x1/x4/a_27_47# 0.378977f
C94 vg1 avss_ip 20.391245f
C95 dvss avss 1.00273f
C96 m1_18932_n17406# avss_ip 0.518743f
C97 dvdd x7/x2/x2/a_27_47# 0.184908f
C98 xin_buf tail 4.362376f
C99 dvdd standby 0.312541f
C100 m1_18932_n15082# avss_ip 0.147881f
C101 dvdd x7/x2/x4/a_27_47# 0.378348f
C102 vg1 dvss_ip 6.367292f
C103 inv_in vg2 0.137694f
C104 xin_buf inv_in 1.533699f
C105 x7/clk_disable dout_filt 0.223819f
C106 avdd_ip inv_in 0.669037f
C107 vrb vg1 0.454276f
C108 inv_in tail 0.604094f
C109 dvss_ip m1_18932_n15082# 0.147461f
C110 m1_2128_n21174# xin 0.159603f
C111 standby_b avss 1.583655f
C112 m1_24530_n19348# avss_ip 0.147859f
C113 avdd_ip avss 0.573261f
C114 x3/out_b avdd 7.478639f
C115 vg1 m1_18932_n15746# 0.267005f
C116 vg1 vg2 1.229449f
C117 xin m1_2130_n19846# 0.165429f
C118 m1_2130_n21506# xin 0.167748f
C119 avdd_ip vg1 1.77908f
C120 m1_2130_n19514# xin 0.164972f
C121 dvdd dvdd_ip 12.609507f
C122 dvdd_ip avdd 0.116559f
C123 dvss_ip m1_24220_n8834# 0.375406f
C124 xout xin 12.304266f
C125 m1_24528_n21342# xin 0.166713f
C126 inv_in avss 0.144174f
C127 dvdd_ip inv_m1 2.234996f
C128 dvdd x7/x1/Qb1 0.459884f
C129 m1_24530_n20676# xin 0.159253f
C130 vbreg xout 16.469566f
C131 x3/out avss 4.193113f
C132 dvdd x7/x1/x2/a_27_47# 0.378403f
C133 dout_ip inv_m2 0.524614f
C134 m1_2130_n20842# xin 0.166057f
C135 avss_ip m1_2132_n17904# 0.186392f
C136 avdd standby_33 5.093125f
C137 m1_2130_n19184# xin 0.164971f
C138 x4/out_b avss 0.261089f
C139 dvdd ena_ip 6.010598f
C140 m1_24530_n20012# avss_ip 0.147858f
C141 dvdd_ip inv_m2 1.267868f
C142 dvdd ena 0.303504f
C143 ena_ip avdd 0.704795f
C144 m1_24530_n20344# xin 0.158905f
C145 icnode avss_ip 31.741272f
C146 avss_ip avdd 2.349381f
C147 dvdd dvss 66.30764f
C148 m1_24528_n22338# avss_ip 0.146396f
C149 m1_2134_n14584# avss_ip 0.746645f
C150 avdd dvss 4.046394f
C151 xin m1_24530_n21008# 0.159641f
C152 m1_18932_n17738# avss_ip 0.587814f
C153 dvdd dvss_ip 20.259176f
C154 m1_2132_n15248# avss_ip 0.200134f
C155 dvdd x7/x2/Qb2 0.448352f
C156 vg2 m1_2132_n17904# 0.154785f
C157 x3/in_b dvss 1.299144f
C158 dvss_ip inv_m1 2.861859f
C159 ibias ibias_ip 0.534567f
C160 m1_18932_n15414# avss_ip 0.17691f
C161 dout dout_filt 0.526935f
C162 dvdd standby_b 4.830365f
C163 icnode vg2 0.394667f
C164 icnode xin_buf 3.629111f
C165 dvss_ip m1_10620_n8006# 0.157361f
C166 standby_b avdd 0.802043f
C167 xin_buf avdd 0.176325f
C168 avss_ip m1_18932_n17074# 0.680482f
C169 icnode avdd_ip 9.185152f
C170 dvdd_ip xin 3.14062f
C171 avdd_ip avdd 8.450802f
C172 m1_2132_n14254# avss_ip 0.740949f
C173 dvss_ip inv_m2 1.434876f
C174 dvdd x7/x1/x3/a_27_47# 0.37895f
C175 standby_ip dvdd_ip 3.47259f
C176 dvss_ip m1_24220_n9166# 0.392413f
C177 dvdd_ip vbreg 0.81911f
C178 m1_2130_n16908# avss_ip 0.190797f
C179 vg2 m1_2132_n15248# 0.154162f
C180 dvdd x7/x2/x3/a_27_47# 0.378322f
C181 m1_24530_n19680# avss_ip 0.147859f
C182 dvdd inv_in 0.696511f
C183 icnode inv_in 0.110238f
C184 xin_buf m1_10620_n8006# 0.166951f
C185 x3/out avdd 5.358785f
C186 m1_2130_n20510# avss_ip 0.188318f
C187 inv_in inv_m1 0.186392f
C188 dvss_ip m1_10620_n9002# 0.146053f
C189 dout_ip dout_filt 2.833564f
C190 xin m1_24528_n22004# 0.166657f
C191 x7/stby_done_b dvss 1.497184f
C192 dvdd avss 0.142936f
C193 avss_ip xin 72.03212f
C194 vn xin 3.076653f
C195 standby_ip ena_ip 4.56584f
C196 avdd avss 62.68863f
C197 dvss_ip x7/stby_done_b 1.502074f
C198 vbreg avss_ip 13.52234f
C199 x7/ena_done_b dvss 1.179651f
C200 x4/out_b avdd 3.554538f
C201 m1_2130_n20180# avss_ip 0.188319f
C202 m1_24530_n21672# xin 0.159429f
C203 dvdd_ip dout_filt 2.111549f
C204 standby_ip dvss 6.437037f
C205 vg2 m1_2130_n16908# 0.156128f
C206 dvss_ip xin 1.630563f
C207 x7/ena_done_b dvss_ip 1.487094f
C208 x3/in_b avss 0.225595f
C209 ibias standby_33 0.82965f
C210 xin_buf m1_10620_n9002# 0.156922f
C211 vg1 m1_18932_n17738# 0.112041f
C212 m1_2130_n21838# xin 0.172287f
C213 dvss_ip vbreg 7.841845f
C214 dvss_ip li_22598_n15512# 0.147611f
C215 vbp ibias_ip 1.263543f
C216 x7/clk_disable dvss 1.678943f
C217 ena_ip ibias 0.172379f
C218 vg1 m1_18932_n15414# 0.560332f
C219 vg2 xin 6.287061f
C220 xin_buf xin 1.993682f
C221 avdd_ip xin 6.041913f
C222 standby_ip standby_b 0.851534f
C223 ibias dvss 1.970363f
C224 vg2 vbreg 4.264934f
C225 tail xin 1.606236f
C226 m1_24530_n19016# xin 0.126575f
C227 avdd_ip vbreg 31.015673f
C228 dout_filt dvss 2.748851f
C229 m1_2132_n17570# avss_ip 0.18406f
C230 dvss_ip dout_filt 7.257841f
C231 inv_in xin 0.302114f
C232 avss_ip m1_2132_n16576# 0.183822f
C233 dvdd_ip xout 3.620201f
C234 m1_2128_n22170# xin 0.284858f
C235 m1_2132_n16242# avss_ip 0.184971f
C236 dvdd x7/x1/x2/a_193_47# 0.105143f
C237 standby_b ibias 0.29964f
C238 m1_2132_n14916# avss_ip 0.607012f
C239 m1_3134_n13314# avss_ip 0.495081f
C240 standby_ip avss 1.62417f
C241 m1_2128_n21174# avss_ip 0.196826f
C242 vg1 xin 6.617878f
C243 avss_ip m1_2130_n17240# 0.190906f
C244 dvdd_ip vbp 18.736547f
C245 dvdd_ip dout 1.175677f
C246 dvdd_ip ibias_ip 1.470902f
C247 dvdd avdd 0.151932f
C248 avss_ip m1_2130_n19846# 0.188318f
C249 m1_2130_n21506# avss_ip 0.188488f
C250 vg1 vbreg 4.57073f
C251 icnode avdd 0.344893f
C252 m1_2130_n19514# avss_ip 0.188318f
C253 vg1 li_22598_n15512# 0.259059f
C254 dvdd x7/x1/Qb2 0.451701f
C255 vg2 m1_2132_n17570# 0.155259f
C256 standby_33 ibias_ip 0.618694f
C257 xout avss_ip 24.57516f
C258 m1_24528_n21342# avss_ip 0.141338f
C259 avss_ip li_8336_n12442# 2.749127f
C260 vg2 m1_2132_n16576# 0.154861f
C261 x3/in_b avdd 0.999306f
C262 dvss_ip m1_10620_n9334# 0.128841f
C263 m1_24530_n20676# avss_ip 0.147859f
C264 m1_2132_n16242# vg2 0.155116f
C265 m1_2130_n20842# avss_ip 0.188487f
C266 m1_24530_n19348# xin 0.159253f
C267 m1_2130_n19184# avss_ip 0.188319f
C268 dvss_ip xout 14.203502f
C269 vg2 m1_2130_n17240# 0.155881f
C270 dout_ip dvdd_ip 1.713335f
C271 inv_m2 inv_m1 0.595615f
C272 ibias_ip dvss 1.192912f
C273 dout dvss 0.170487f
C274 m1_18932_n16078# avss_ip 0.49845f
C275 xin_buf m1_10620_n9334# 0.138691f
C276 m1_24530_n20344# avss_ip 0.147654f
C277 dvss_ip vbp 1.256699f
C278 dvss_ip ibias_ip 18.52148f
C279 dvss_ip dout 6.565475f
C280 m1_18932_n16410# avss_ip 0.64459f
C281 vg2 xout 0.938911f
C282 m1_10620_n9664# li_9150_n9268# 0.106769f
C283 dvdd_ip li_9150_n9268# 0.603132f
C284 xin_buf xout 3.498235f
C285 avdd_ip xout 6.529395f
C286 standby dvss 0.267007f
C287 avss_ip m1_24530_n21008# 0.148183f
C288 xin_buf li_8336_n12442# 0.264063f
C289 xout tail 1.225035f
C290 dvdd x7/stby_done_b 2.392811f
C291 dvdd_ip standby_33 3.319999f
C292 dvss_ip m1_10620_n8670# 0.157269f
C293 xin_buf vbp 3.475593f
C294 dvss_ip m1_24220_n7840# 0.356811f
C295 xin_buf ibias_ip 1.728949f
C296 m1_24530_n20012# xin 0.159204f
C297 dvdd x7/ena_done_b 2.894243f
C298 vbp tail 10.071224f
C299 inv_in xout 1.165599f
C300 dout_ip dvss 2.669038f
C301 standby_ip dvdd 7.333838f
C302 dvss_ip m1_24220_n8502# 0.389794f
C303 avss_ip m1_2130_n15578# 0.196054f
C304 standby_ip avdd 0.683223f
C305 m1_24528_n22338# xin 0.168028f
C306 dvdd_ip avss_ip 2.34725f
C307 vn dvdd_ip 0.861771f
C308 dout_ip dvss_ip 6.656641f
C309 m1_24530_n19348# amp_XM16_17/0. 0.236835f
C310 m1_2130_n20842# amp_XM16_17/0. 0.251456f
C311 m1_2132_n17904# amp_XM16_17/0. 0.250246f
C312 m1_2132_n16576# amp_XM16_17/0. 0.250246f
C313 m1_2132_n15248# amp_XM16_17/0. 0.250246f
C314 m1_10620_n9664# amp_XM16_17/0. 0.232743f
C315 m1_24220_n8172# amp_XM16_17/0. 0.251507f
C316 vg1 amp_XM16_17/0. 9.89592f
C317 avss_ip amp_XM16_17/0. -26.136543f
C318 dvss_ip amp_XM16_17/0. 32.94271f
C319 tail amp_XM16_17/0. 0.375175f
C320 vbp amp_XM16_17/0. 3.494732f
C321 vrb amp_XM16_17/0. 0.162439f
C322 li_8336_n12442# amp_XM16_17/0. 1.864265f
C323 inv_m2 amp_XM16_17/0. 0.74678f
C324 inv_m1 amp_XM16_17/0. 0.894821f
C325 avdd_ip amp_XM16_17/0. 0.283987p
C326 xin_buf amp_XM16_17/0. 25.955637f
C327 vn amp_XM16_17/0. 2.283171f
C328 ibias_ip amp_XM16_17/0. 4.323137f
C329 standby_ip amp_XM16_17/0. 7.853122f
C330 ibias amp_XM16_17/0. 3.711352f
C331 x3/out_b amp_XM16_17/0. 1.159828f
C332 avdd amp_XM16_17/0. 85.680984f
C333 vbreg amp_XM16_17/0. 4.472168f
C334 vg2 amp_XM16_17/0. 10.895053f
C335 x3/out amp_XM16_17/0. 1.415974f
C336 xout amp_XM16_17/0. 3.165308f
C337 inv_in amp_XM16_17/0. 12.857133f
C338 dout amp_XM16_17/0. 0.19266f
C339 xin amp_XM16_17/0. 16.293684f
C340 dvdd_ip amp_XM16_17/0. 0.300975p
C341 m1_24528_n22338# amp_XM16_17/0. 0.24285f
C342 m1_2128_n22170# amp_XM16_17/0. 0.245373f
C343 m1_24528_n22004# amp_XM16_17/0. 0.24291f
C344 m1_2130_n21838# amp_XM16_17/0. 0.251475f
C345 m1_24530_n21672# amp_XM16_17/0. 0.236835f
C346 m1_2130_n21506# amp_XM16_17/0. 0.251455f
C347 m1_24528_n21342# amp_XM16_17/0. 0.243274f
C348 m1_2128_n21174# amp_XM16_17/0. 0.245478f
C349 m1_24530_n21008# amp_XM16_17/0. 0.236835f
C350 m1_24530_n20676# amp_XM16_17/0. 0.236835f
C351 m1_2130_n20510# amp_XM16_17/0. 0.251298f
C352 m1_24530_n20344# amp_XM16_17/0. 0.236676f
C353 m1_2130_n20180# amp_XM16_17/0. 0.251301f
C354 m1_24530_n20012# amp_XM16_17/0. 0.236739f
C355 m1_2130_n19846# amp_XM16_17/0. 0.251304f
C356 m1_24530_n19680# amp_XM16_17/0. 0.236835f
C357 m1_2130_n19514# amp_XM16_17/0. 0.251298f
C358 m1_2130_n19184# amp_XM16_17/0. 0.251301f
C359 m1_24530_n19016# amp_XM16_17/0. 0.236835f
C360 m1_2130_n18850# amp_XM16_17/0. 0.251304f
C361 icnode amp_XM16_17/0. 11.843518f
C362 dout_filt amp_XM16_17/0. 1.415894f
C363 x7/clk_disable amp_XM16_17/0. 2.783535f
C364 x7/x5/a_30_47# amp_XM16_17/0. 0.145562f
C365 x7/x3/a_27_47# amp_XM16_17/0. 0.216317f $ **FLOATING
C366 x7/x2/x4/a_1847_47# amp_XM16_17/0. 0.132899f
C367 x7/x2/x4/a_1108_47# amp_XM16_17/0. 0.126214f $ **FLOATING
C368 x7/x2/x4/a_1283_21# amp_XM16_17/0. 0.478567f $ **FLOATING
C369 x7/x2/x4/a_543_47# amp_XM16_17/0. 0.157869f $ **FLOATING
C370 x7/x2/x4/a_761_289# amp_XM16_17/0. 0.120848f $ **FLOATING
C371 x7/x2/x4/a_193_47# amp_XM16_17/0. 0.272684f
C372 x7/x2/x4/a_27_47# amp_XM16_17/0. 0.495665f
C373 dvdd amp_XM16_17/0. 31.67741f
C374 x7/x2/Qb1 amp_XM16_17/0. 0.335308f
C375 x7/x2/x1/X amp_XM16_17/0. 0.180099f
C376 x7/x2/x2/a_1847_47# amp_XM16_17/0. 0.132899f
C377 x7/x2/x2/a_1108_47# amp_XM16_17/0. 0.126214f $ **FLOATING
C378 x7/x2/x2/a_1283_21# amp_XM16_17/0. 0.478567f $ **FLOATING
C379 x7/x2/x2/a_543_47# amp_XM16_17/0. 0.157869f $ **FLOATING
C380 x7/x2/x2/a_761_289# amp_XM16_17/0. 0.120848f $ **FLOATING
C381 x7/x2/x2/a_193_47# amp_XM16_17/0. 0.272684f
C382 x7/x2/x2/a_27_47# amp_XM16_17/0. 0.495665f
C383 x7/x2/Qb2 amp_XM16_17/0. 0.335611f
C384 x7/x2/x3/a_1847_47# amp_XM16_17/0. 0.132899f
C385 x7/x2/x3/a_1108_47# amp_XM16_17/0. 0.126214f $ **FLOATING
C386 x7/x2/x3/a_1283_21# amp_XM16_17/0. 0.478567f $ **FLOATING
C387 x7/x2/x3/a_543_47# amp_XM16_17/0. 0.157869f $ **FLOATING
C388 x7/x2/x3/a_761_289# amp_XM16_17/0. 0.120848f $ **FLOATING
C389 x7/x2/x3/a_193_47# amp_XM16_17/0. 0.272684f
C390 x7/x2/x3/a_27_47# amp_XM16_17/0. 0.495665f
C391 x7/stby_done_b amp_XM16_17/0. 1.263094f
C392 dout_ip amp_XM16_17/0. 2.177488f
C393 x7/x2/x1/a_40_47# amp_XM16_17/0. 0.230074f $ **FLOATING
C394 x7/x1/x4/a_1847_47# amp_XM16_17/0. 0.132899f
C395 x7/x1/x4/a_1108_47# amp_XM16_17/0. 0.126214f $ **FLOATING
C396 x7/x1/x4/a_1283_21# amp_XM16_17/0. 0.478567f $ **FLOATING
C397 x7/x1/x4/a_543_47# amp_XM16_17/0. 0.157869f $ **FLOATING
C398 x7/x1/x4/a_761_289# amp_XM16_17/0. 0.120848f $ **FLOATING
C399 x7/x1/x4/a_193_47# amp_XM16_17/0. 0.272684f
C400 x7/x1/x4/a_27_47# amp_XM16_17/0. 0.495665f
C401 dvss amp_XM16_17/0. 30.006504f
C402 ena_ip amp_XM16_17/0. 3.095204f
C403 x7/x1/Qb1 amp_XM16_17/0. 0.335308f
C404 x7/x1/x1/X amp_XM16_17/0. 0.180099f
C405 x7/x1/x2/a_1847_47# amp_XM16_17/0. 0.132899f
C406 x7/x1/x2/a_1108_47# amp_XM16_17/0. 0.126214f $ **FLOATING
C407 x7/x1/x2/a_1283_21# amp_XM16_17/0. 0.478567f $ **FLOATING
C408 x7/x1/x2/a_543_47# amp_XM16_17/0. 0.157869f $ **FLOATING
C409 x7/x1/x2/a_761_289# amp_XM16_17/0. 0.120848f $ **FLOATING
C410 x7/x1/x2/a_193_47# amp_XM16_17/0. 0.272684f
C411 x7/x1/x2/a_27_47# amp_XM16_17/0. 0.495665f
C412 x7/x1/Qb2 amp_XM16_17/0. 0.335611f
C413 x7/x1/x3/a_1847_47# amp_XM16_17/0. 0.132899f
C414 x7/x1/x3/a_1108_47# amp_XM16_17/0. 0.126214f $ **FLOATING
C415 x7/x1/x3/a_1283_21# amp_XM16_17/0. 0.478567f $ **FLOATING
C416 x7/x1/x3/a_543_47# amp_XM16_17/0. 0.157869f $ **FLOATING
C417 x7/x1/x3/a_761_289# amp_XM16_17/0. 0.120848f $ **FLOATING
C418 x7/x1/x3/a_193_47# amp_XM16_17/0. 0.272684f
C419 x7/x1/x3/a_27_47# amp_XM16_17/0. 0.495665f
C420 x7/ena_done_b amp_XM16_17/0. 1.398332f
C421 x7/x1/x1/a_40_47# amp_XM16_17/0. 0.230074f $ **FLOATING
C422 standby_33 amp_XM16_17/0. 2.68323f
C423 standby_b amp_XM16_17/0. 6.77451f
C424 x4/out_b amp_XM16_17/0. 1.23154f
C425 avss amp_XM16_17/0. 3.020541f
C426 x3/in_b amp_XM16_17/0. 1.286801f
C427 standby amp_XM16_17/0. 1.021767f
C428 x2/a_27_47# amp_XM16_17/0. 0.207781f $ **FLOATING
C429 m1_3134_n13314# amp_XM16_17/0. 0.236373f
C430 ena amp_XM16_17/0. 1.000301f
C431 x1/a_27_47# amp_XM16_17/0. 0.207781f $ **FLOATING
C432 m1_18932_n17738# amp_XM16_17/0. 0.228879f
C433 m1_2132_n17570# amp_XM16_17/0. 0.250378f
C434 m1_18932_n17406# amp_XM16_17/0. 0.228879f
C435 m1_2130_n17240# amp_XM16_17/0. 0.245126f
C436 m1_18932_n17074# amp_XM16_17/0. 0.228879f
C437 m1_2130_n16908# amp_XM16_17/0. 0.245126f
C438 m1_18932_n16742# amp_XM16_17/0. 0.228879f
C439 m1_18932_n16410# amp_XM16_17/0. 0.228879f
C440 m1_2132_n16242# amp_XM16_17/0. 0.250378f
C441 m1_18932_n16078# amp_XM16_17/0. 0.228879f
C442 m1_2132_n15912# amp_XM16_17/0. 0.250246f
C443 m1_18932_n15746# amp_XM16_17/0. 0.228742f
C444 m1_2130_n15578# amp_XM16_17/0. 0.245259f
C445 m1_18932_n15414# amp_XM16_17/0. 0.227965f
C446 m1_18932_n15082# amp_XM16_17/0. 0.253441f
C447 m1_2132_n14916# amp_XM16_17/0. 0.250246f
C448 m1_18932_n14750# amp_XM16_17/0. 0.250246f
C449 m1_2134_n14584# amp_XM16_17/0. 0.250905f
C450 m1_18932_n14418# amp_XM16_17/0. 0.22541f
C451 m1_2132_n14254# amp_XM16_17/0. 0.250378f
C452 li_9150_n9268# amp_XM16_17/0. 3.463315f
C453 m1_24220_n9832# amp_XM16_17/0. 0.395618f
C454 m1_24220_n9500# amp_XM16_17/0. 0.251874f
C455 m1_10620_n9334# amp_XM16_17/0. 0.251414f
C456 m1_24220_n9166# amp_XM16_17/0. 0.232835f
C457 m1_10620_n9002# amp_XM16_17/0. 0.25178f
C458 m1_24220_n8834# amp_XM16_17/0. 0.232468f
C459 m1_10620_n8670# amp_XM16_17/0. 0.25178f
C460 m1_24220_n8502# amp_XM16_17/0. 0.232468f
C461 m1_10620_n8338# amp_XM16_17/0. 0.25178f
C462 m1_10620_n8006# amp_XM16_17/0. 0.25178f
C463 m1_24220_n7840# amp_XM16_17/0. 0.251874f
C464 m1_10618_n7674# amp_XM16_17/0. 0.389918f
.ends

