magic
tech sky130A
magscale 1 2
timestamp 1713142410
<< metal3 >>
rect -2492 120 -412 2200
rect -136 122 1948 2202
rect -2490 -2254 -410 -174
rect -134 -2252 1950 -172
<< mimcap >>
rect -2452 2120 -452 2160
rect -2452 200 -2412 2120
rect -492 200 -452 2120
rect -2452 160 -452 200
rect -96 2122 1904 2162
rect -96 202 -56 2122
rect 1864 202 1904 2122
rect -96 162 1904 202
rect -2450 -254 -450 -214
rect -2450 -2174 -2410 -254
rect -490 -2174 -450 -254
rect -2450 -2214 -450 -2174
rect -94 -252 1906 -212
rect -94 -2172 -54 -252
rect 1866 -2172 1906 -252
rect -94 -2212 1906 -2172
<< mimcapcontact >>
rect -2412 200 -492 2120
rect -56 202 1864 2122
rect -2410 -2174 -490 -254
rect -54 -2172 1866 -252
<< metal4 >>
rect -1504 2121 -1400 2220
rect 852 2123 956 2222
rect -57 2122 1865 2123
rect -2413 2120 -491 2121
rect -2413 200 -2412 2120
rect -492 1948 -491 2120
rect -57 1948 -56 2122
rect -492 1622 -56 1948
rect -492 200 -491 1622
rect -57 202 -56 1622
rect 1864 202 1865 2122
rect -57 201 1865 202
rect -2413 199 -491 200
rect -1630 -253 -1264 199
rect 714 -251 1080 201
rect -55 -252 1867 -251
rect -2411 -254 -489 -253
rect -2411 -2174 -2410 -254
rect -490 -1460 -489 -254
rect -55 -1460 -54 -252
rect -490 -1786 -54 -1460
rect -490 -2174 -489 -1786
rect -55 -2172 -54 -1786
rect 1866 -2172 1867 -252
rect -55 -2173 1867 -2172
rect -2411 -2175 -489 -2174
rect -1502 -2268 -1398 -2175
rect 854 -2266 958 -2173
<< properties >>
string FIXED_BBOX 120 120 2200 2200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
