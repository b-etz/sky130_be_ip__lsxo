magic
tech sky130A
magscale 1 2
timestamp 1712782684
<< nwell >>
rect -1374 -1215 1374 1215
<< mvpmos >>
rect -1116 118 -716 918
rect -658 118 -258 918
rect -200 118 200 918
rect 258 118 658 918
rect 716 118 1116 918
rect -1116 -918 -716 -118
rect -658 -918 -258 -118
rect -200 -918 200 -118
rect 258 -918 658 -118
rect 716 -918 1116 -118
<< mvpdiff >>
rect -1174 906 -1116 918
rect -1174 130 -1162 906
rect -1128 130 -1116 906
rect -1174 118 -1116 130
rect -716 906 -658 918
rect -716 130 -704 906
rect -670 130 -658 906
rect -716 118 -658 130
rect -258 906 -200 918
rect -258 130 -246 906
rect -212 130 -200 906
rect -258 118 -200 130
rect 200 906 258 918
rect 200 130 212 906
rect 246 130 258 906
rect 200 118 258 130
rect 658 906 716 918
rect 658 130 670 906
rect 704 130 716 906
rect 658 118 716 130
rect 1116 906 1174 918
rect 1116 130 1128 906
rect 1162 130 1174 906
rect 1116 118 1174 130
rect -1174 -130 -1116 -118
rect -1174 -906 -1162 -130
rect -1128 -906 -1116 -130
rect -1174 -918 -1116 -906
rect -716 -130 -658 -118
rect -716 -906 -704 -130
rect -670 -906 -658 -130
rect -716 -918 -658 -906
rect -258 -130 -200 -118
rect -258 -906 -246 -130
rect -212 -906 -200 -130
rect -258 -918 -200 -906
rect 200 -130 258 -118
rect 200 -906 212 -130
rect 246 -906 258 -130
rect 200 -918 258 -906
rect 658 -130 716 -118
rect 658 -906 670 -130
rect 704 -906 716 -130
rect 658 -918 716 -906
rect 1116 -130 1174 -118
rect 1116 -906 1128 -130
rect 1162 -906 1174 -130
rect 1116 -918 1174 -906
<< mvpdiffc >>
rect -1162 130 -1128 906
rect -704 130 -670 906
rect -246 130 -212 906
rect 212 130 246 906
rect 670 130 704 906
rect 1128 130 1162 906
rect -1162 -906 -1128 -130
rect -704 -906 -670 -130
rect -246 -906 -212 -130
rect 212 -906 246 -130
rect 670 -906 704 -130
rect 1128 -906 1162 -130
<< mvnsubdiff >>
rect -1308 1137 1308 1149
rect -1308 1103 -1200 1137
rect 1200 1103 1308 1137
rect -1308 1091 1308 1103
rect -1308 1041 -1250 1091
rect -1308 -1041 -1296 1041
rect -1262 -1041 -1250 1041
rect 1250 1041 1308 1091
rect -1308 -1091 -1250 -1041
rect 1250 -1041 1262 1041
rect 1296 -1041 1308 1041
rect 1250 -1091 1308 -1041
rect -1308 -1103 1308 -1091
rect -1308 -1137 -1200 -1103
rect 1200 -1137 1308 -1103
rect -1308 -1149 1308 -1137
<< mvnsubdiffcont >>
rect -1200 1103 1200 1137
rect -1296 -1041 -1262 1041
rect 1262 -1041 1296 1041
rect -1200 -1137 1200 -1103
<< poly >>
rect -1116 999 -716 1015
rect -1116 965 -1100 999
rect -732 965 -716 999
rect -1116 918 -716 965
rect -658 999 -258 1015
rect -658 965 -642 999
rect -274 965 -258 999
rect -658 918 -258 965
rect -200 999 200 1015
rect -200 965 -184 999
rect 184 965 200 999
rect -200 918 200 965
rect 258 999 658 1015
rect 258 965 274 999
rect 642 965 658 999
rect 258 918 658 965
rect 716 999 1116 1015
rect 716 965 732 999
rect 1100 965 1116 999
rect 716 918 1116 965
rect -1116 71 -716 118
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -1116 21 -716 37
rect -658 71 -258 118
rect -658 37 -642 71
rect -274 37 -258 71
rect -658 21 -258 37
rect -200 71 200 118
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect 258 71 658 118
rect 258 37 274 71
rect 642 37 658 71
rect 258 21 658 37
rect 716 71 1116 118
rect 716 37 732 71
rect 1100 37 1116 71
rect 716 21 1116 37
rect -1116 -37 -716 -21
rect -1116 -71 -1100 -37
rect -732 -71 -716 -37
rect -1116 -118 -716 -71
rect -658 -37 -258 -21
rect -658 -71 -642 -37
rect -274 -71 -258 -37
rect -658 -118 -258 -71
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -118 200 -71
rect 258 -37 658 -21
rect 258 -71 274 -37
rect 642 -71 658 -37
rect 258 -118 658 -71
rect 716 -37 1116 -21
rect 716 -71 732 -37
rect 1100 -71 1116 -37
rect 716 -118 1116 -71
rect -1116 -965 -716 -918
rect -1116 -999 -1100 -965
rect -732 -999 -716 -965
rect -1116 -1015 -716 -999
rect -658 -965 -258 -918
rect -658 -999 -642 -965
rect -274 -999 -258 -965
rect -658 -1015 -258 -999
rect -200 -965 200 -918
rect -200 -999 -184 -965
rect 184 -999 200 -965
rect -200 -1015 200 -999
rect 258 -965 658 -918
rect 258 -999 274 -965
rect 642 -999 658 -965
rect 258 -1015 658 -999
rect 716 -965 1116 -918
rect 716 -999 732 -965
rect 1100 -999 1116 -965
rect 716 -1015 1116 -999
<< polycont >>
rect -1100 965 -732 999
rect -642 965 -274 999
rect -184 965 184 999
rect 274 965 642 999
rect 732 965 1100 999
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect -1100 -71 -732 -37
rect -642 -71 -274 -37
rect -184 -71 184 -37
rect 274 -71 642 -37
rect 732 -71 1100 -37
rect -1100 -999 -732 -965
rect -642 -999 -274 -965
rect -184 -999 184 -965
rect 274 -999 642 -965
rect 732 -999 1100 -965
<< locali >>
rect -1296 1103 -1200 1137
rect 1200 1103 1296 1137
rect -1296 1041 -1262 1103
rect 1262 1041 1296 1103
rect -1116 965 -1100 999
rect -732 965 -716 999
rect -658 965 -642 999
rect -274 965 -258 999
rect -200 965 -184 999
rect 184 965 200 999
rect 258 965 274 999
rect 642 965 658 999
rect 716 965 732 999
rect 1100 965 1116 999
rect -1162 906 -1128 922
rect -1162 114 -1128 130
rect -704 906 -670 922
rect -704 114 -670 130
rect -246 906 -212 922
rect -246 114 -212 130
rect 212 906 246 922
rect 212 114 246 130
rect 670 906 704 922
rect 670 114 704 130
rect 1128 906 1162 922
rect 1128 114 1162 130
rect -1116 37 -1100 71
rect -732 37 -716 71
rect -658 37 -642 71
rect -274 37 -258 71
rect -200 37 -184 71
rect 184 37 200 71
rect 258 37 274 71
rect 642 37 658 71
rect 716 37 732 71
rect 1100 37 1116 71
rect -1116 -71 -1100 -37
rect -732 -71 -716 -37
rect -658 -71 -642 -37
rect -274 -71 -258 -37
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect 258 -71 274 -37
rect 642 -71 658 -37
rect 716 -71 732 -37
rect 1100 -71 1116 -37
rect -1162 -130 -1128 -114
rect -1162 -922 -1128 -906
rect -704 -130 -670 -114
rect -704 -922 -670 -906
rect -246 -130 -212 -114
rect -246 -922 -212 -906
rect 212 -130 246 -114
rect 212 -922 246 -906
rect 670 -130 704 -114
rect 670 -922 704 -906
rect 1128 -130 1162 -114
rect 1128 -922 1162 -906
rect -1116 -999 -1100 -965
rect -732 -999 -716 -965
rect -658 -999 -642 -965
rect -274 -999 -258 -965
rect -200 -999 -184 -965
rect 184 -999 200 -965
rect 258 -999 274 -965
rect 642 -999 658 -965
rect 716 -999 732 -965
rect 1100 -999 1116 -965
rect -1296 -1103 -1262 -1041
rect 1262 -1103 1296 -1041
rect -1296 -1137 -1200 -1103
rect 1200 -1137 1296 -1103
<< viali >>
rect -1100 965 -732 999
rect -642 965 -274 999
rect -184 965 184 999
rect 274 965 642 999
rect 732 965 1100 999
rect -1162 130 -1128 906
rect -704 130 -670 906
rect -246 130 -212 906
rect 212 130 246 906
rect 670 130 704 906
rect 1128 130 1162 906
rect -1100 37 -732 71
rect -642 37 -274 71
rect -184 37 184 71
rect 274 37 642 71
rect 732 37 1100 71
rect -1100 -71 -732 -37
rect -642 -71 -274 -37
rect -184 -71 184 -37
rect 274 -71 642 -37
rect 732 -71 1100 -37
rect -1162 -906 -1128 -130
rect -704 -906 -670 -130
rect -246 -906 -212 -130
rect 212 -906 246 -130
rect 670 -906 704 -130
rect 1128 -906 1162 -130
rect -1100 -999 -732 -965
rect -642 -999 -274 -965
rect -184 -999 184 -965
rect 274 -999 642 -965
rect 732 -999 1100 -965
<< metal1 >>
rect -1112 999 -720 1005
rect -1112 965 -1100 999
rect -732 965 -720 999
rect -1112 959 -720 965
rect -654 999 -262 1005
rect -654 965 -642 999
rect -274 965 -262 999
rect -654 959 -262 965
rect -196 999 196 1005
rect -196 965 -184 999
rect 184 965 196 999
rect -196 959 196 965
rect 262 999 654 1005
rect 262 965 274 999
rect 642 965 654 999
rect 262 959 654 965
rect 720 999 1112 1005
rect 720 965 732 999
rect 1100 965 1112 999
rect 720 959 1112 965
rect -1168 906 -1122 918
rect -1168 130 -1162 906
rect -1128 130 -1122 906
rect -1168 118 -1122 130
rect -710 906 -664 918
rect -710 130 -704 906
rect -670 130 -664 906
rect -710 118 -664 130
rect -252 906 -206 918
rect -252 130 -246 906
rect -212 130 -206 906
rect -252 118 -206 130
rect 206 906 252 918
rect 206 130 212 906
rect 246 130 252 906
rect 206 118 252 130
rect 664 906 710 918
rect 664 130 670 906
rect 704 130 710 906
rect 664 118 710 130
rect 1122 906 1168 918
rect 1122 130 1128 906
rect 1162 130 1168 906
rect 1122 118 1168 130
rect -1112 71 -720 77
rect -1112 37 -1100 71
rect -732 37 -720 71
rect -1112 31 -720 37
rect -654 71 -262 77
rect -654 37 -642 71
rect -274 37 -262 71
rect -654 31 -262 37
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect 262 71 654 77
rect 262 37 274 71
rect 642 37 654 71
rect 262 31 654 37
rect 720 71 1112 77
rect 720 37 732 71
rect 1100 37 1112 71
rect 720 31 1112 37
rect -1112 -37 -720 -31
rect -1112 -71 -1100 -37
rect -732 -71 -720 -37
rect -1112 -77 -720 -71
rect -654 -37 -262 -31
rect -654 -71 -642 -37
rect -274 -71 -262 -37
rect -654 -77 -262 -71
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect 262 -37 654 -31
rect 262 -71 274 -37
rect 642 -71 654 -37
rect 262 -77 654 -71
rect 720 -37 1112 -31
rect 720 -71 732 -37
rect 1100 -71 1112 -37
rect 720 -77 1112 -71
rect -1168 -130 -1122 -118
rect -1168 -906 -1162 -130
rect -1128 -906 -1122 -130
rect -1168 -918 -1122 -906
rect -710 -130 -664 -118
rect -710 -906 -704 -130
rect -670 -906 -664 -130
rect -710 -918 -664 -906
rect -252 -130 -206 -118
rect -252 -906 -246 -130
rect -212 -906 -206 -130
rect -252 -918 -206 -906
rect 206 -130 252 -118
rect 206 -906 212 -130
rect 246 -906 252 -130
rect 206 -918 252 -906
rect 664 -130 710 -118
rect 664 -906 670 -130
rect 704 -906 710 -130
rect 664 -918 710 -906
rect 1122 -130 1168 -118
rect 1122 -906 1128 -130
rect 1162 -906 1168 -130
rect 1122 -918 1168 -906
rect -1112 -965 -720 -959
rect -1112 -999 -1100 -965
rect -732 -999 -720 -965
rect -1112 -1005 -720 -999
rect -654 -965 -262 -959
rect -654 -999 -642 -965
rect -274 -999 -262 -965
rect -654 -1005 -262 -999
rect -196 -965 196 -959
rect -196 -999 -184 -965
rect 184 -999 196 -965
rect -196 -1005 196 -999
rect 262 -965 654 -959
rect 262 -999 274 -965
rect 642 -999 654 -965
rect 262 -1005 654 -999
rect 720 -965 1112 -959
rect 720 -999 732 -965
rect 1100 -999 1112 -965
rect 720 -1005 1112 -999
<< properties >>
string FIXED_BBOX -1279 -1120 1279 1120
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 2.0 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
