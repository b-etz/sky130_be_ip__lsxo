magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< nwell >>
rect -308 -2769 308 2769
<< mvpmos >>
rect -50 1672 50 2472
rect -50 636 50 1436
rect -50 -400 50 400
rect -50 -1436 50 -636
rect -50 -2472 50 -1672
<< mvpdiff >>
rect -108 2460 -50 2472
rect -108 1684 -96 2460
rect -62 1684 -50 2460
rect -108 1672 -50 1684
rect 50 2460 108 2472
rect 50 1684 62 2460
rect 96 1684 108 2460
rect 50 1672 108 1684
rect -108 1424 -50 1436
rect -108 648 -96 1424
rect -62 648 -50 1424
rect -108 636 -50 648
rect 50 1424 108 1436
rect 50 648 62 1424
rect 96 648 108 1424
rect 50 636 108 648
rect -108 388 -50 400
rect -108 -388 -96 388
rect -62 -388 -50 388
rect -108 -400 -50 -388
rect 50 388 108 400
rect 50 -388 62 388
rect 96 -388 108 388
rect 50 -400 108 -388
rect -108 -648 -50 -636
rect -108 -1424 -96 -648
rect -62 -1424 -50 -648
rect -108 -1436 -50 -1424
rect 50 -648 108 -636
rect 50 -1424 62 -648
rect 96 -1424 108 -648
rect 50 -1436 108 -1424
rect -108 -1684 -50 -1672
rect -108 -2460 -96 -1684
rect -62 -2460 -50 -1684
rect -108 -2472 -50 -2460
rect 50 -1684 108 -1672
rect 50 -2460 62 -1684
rect 96 -2460 108 -1684
rect 50 -2472 108 -2460
<< mvpdiffc >>
rect -96 1684 -62 2460
rect 62 1684 96 2460
rect -96 648 -62 1424
rect 62 648 96 1424
rect -96 -388 -62 388
rect 62 -388 96 388
rect -96 -1424 -62 -648
rect 62 -1424 96 -648
rect -96 -2460 -62 -1684
rect 62 -2460 96 -1684
<< mvnsubdiff >>
rect -242 2691 242 2703
rect -242 2657 -134 2691
rect 134 2657 242 2691
rect -242 2645 242 2657
rect -242 2595 -184 2645
rect -242 -2595 -230 2595
rect -196 -2595 -184 2595
rect 184 2595 242 2645
rect -242 -2645 -184 -2595
rect 184 -2595 196 2595
rect 230 -2595 242 2595
rect 184 -2645 242 -2595
rect -242 -2657 242 -2645
rect -242 -2691 -134 -2657
rect 134 -2691 242 -2657
rect -242 -2703 242 -2691
<< mvnsubdiffcont >>
rect -134 2657 134 2691
rect -230 -2595 -196 2595
rect 196 -2595 230 2595
rect -134 -2691 134 -2657
<< poly >>
rect -50 2553 50 2569
rect -50 2519 -34 2553
rect 34 2519 50 2553
rect -50 2472 50 2519
rect -50 1625 50 1672
rect -50 1591 -34 1625
rect 34 1591 50 1625
rect -50 1575 50 1591
rect -50 1517 50 1533
rect -50 1483 -34 1517
rect 34 1483 50 1517
rect -50 1436 50 1483
rect -50 589 50 636
rect -50 555 -34 589
rect 34 555 50 589
rect -50 539 50 555
rect -50 481 50 497
rect -50 447 -34 481
rect 34 447 50 481
rect -50 400 50 447
rect -50 -447 50 -400
rect -50 -481 -34 -447
rect 34 -481 50 -447
rect -50 -497 50 -481
rect -50 -555 50 -539
rect -50 -589 -34 -555
rect 34 -589 50 -555
rect -50 -636 50 -589
rect -50 -1483 50 -1436
rect -50 -1517 -34 -1483
rect 34 -1517 50 -1483
rect -50 -1533 50 -1517
rect -50 -1591 50 -1575
rect -50 -1625 -34 -1591
rect 34 -1625 50 -1591
rect -50 -1672 50 -1625
rect -50 -2519 50 -2472
rect -50 -2553 -34 -2519
rect 34 -2553 50 -2519
rect -50 -2569 50 -2553
<< polycont >>
rect -34 2519 34 2553
rect -34 1591 34 1625
rect -34 1483 34 1517
rect -34 555 34 589
rect -34 447 34 481
rect -34 -481 34 -447
rect -34 -589 34 -555
rect -34 -1517 34 -1483
rect -34 -1625 34 -1591
rect -34 -2553 34 -2519
<< locali >>
rect -230 2657 -134 2691
rect 134 2657 230 2691
rect -230 2595 -196 2657
rect 196 2595 230 2657
rect -50 2519 -34 2553
rect 34 2519 50 2553
rect -96 2460 -62 2476
rect -96 1668 -62 1684
rect 62 2460 96 2476
rect 62 1668 96 1684
rect -50 1591 -34 1625
rect 34 1591 50 1625
rect -50 1483 -34 1517
rect 34 1483 50 1517
rect -96 1424 -62 1440
rect -96 632 -62 648
rect 62 1424 96 1440
rect 62 632 96 648
rect -50 555 -34 589
rect 34 555 50 589
rect -50 447 -34 481
rect 34 447 50 481
rect -96 388 -62 404
rect -96 -404 -62 -388
rect 62 388 96 404
rect 62 -404 96 -388
rect -50 -481 -34 -447
rect 34 -481 50 -447
rect -50 -589 -34 -555
rect 34 -589 50 -555
rect -96 -648 -62 -632
rect -96 -1440 -62 -1424
rect 62 -648 96 -632
rect 62 -1440 96 -1424
rect -50 -1517 -34 -1483
rect 34 -1517 50 -1483
rect -50 -1625 -34 -1591
rect 34 -1625 50 -1591
rect -96 -1684 -62 -1668
rect -96 -2476 -62 -2460
rect 62 -1684 96 -1668
rect 62 -2476 96 -2460
rect -50 -2553 -34 -2519
rect 34 -2553 50 -2519
rect -230 -2657 -196 -2595
rect 196 -2657 230 -2595
rect -230 -2691 -134 -2657
rect 134 -2691 230 -2657
<< viali >>
rect -34 2519 34 2553
rect -96 1684 -62 2460
rect 62 1684 96 2460
rect -34 1591 34 1625
rect -34 1483 34 1517
rect -96 648 -62 1424
rect 62 648 96 1424
rect -34 555 34 589
rect -34 447 34 481
rect -96 -388 -62 388
rect 62 -388 96 388
rect -34 -481 34 -447
rect -34 -589 34 -555
rect -96 -1424 -62 -648
rect 62 -1424 96 -648
rect -34 -1517 34 -1483
rect -34 -1625 34 -1591
rect -96 -2460 -62 -1684
rect 62 -2460 96 -1684
rect -34 -2553 34 -2519
<< metal1 >>
rect -46 2553 46 2559
rect -46 2519 -34 2553
rect 34 2519 46 2553
rect -46 2513 46 2519
rect -102 2460 -56 2472
rect -102 1684 -96 2460
rect -62 1684 -56 2460
rect -102 1672 -56 1684
rect 56 2460 102 2472
rect 56 1684 62 2460
rect 96 1684 102 2460
rect 56 1672 102 1684
rect -46 1625 46 1631
rect -46 1591 -34 1625
rect 34 1591 46 1625
rect -46 1585 46 1591
rect -46 1517 46 1523
rect -46 1483 -34 1517
rect 34 1483 46 1517
rect -46 1477 46 1483
rect -102 1424 -56 1436
rect -102 648 -96 1424
rect -62 648 -56 1424
rect -102 636 -56 648
rect 56 1424 102 1436
rect 56 648 62 1424
rect 96 648 102 1424
rect 56 636 102 648
rect -46 589 46 595
rect -46 555 -34 589
rect 34 555 46 589
rect -46 549 46 555
rect -46 481 46 487
rect -46 447 -34 481
rect 34 447 46 481
rect -46 441 46 447
rect -102 388 -56 400
rect -102 -388 -96 388
rect -62 -388 -56 388
rect -102 -400 -56 -388
rect 56 388 102 400
rect 56 -388 62 388
rect 96 -388 102 388
rect 56 -400 102 -388
rect -46 -447 46 -441
rect -46 -481 -34 -447
rect 34 -481 46 -447
rect -46 -487 46 -481
rect -46 -555 46 -549
rect -46 -589 -34 -555
rect 34 -589 46 -555
rect -46 -595 46 -589
rect -102 -648 -56 -636
rect -102 -1424 -96 -648
rect -62 -1424 -56 -648
rect -102 -1436 -56 -1424
rect 56 -648 102 -636
rect 56 -1424 62 -648
rect 96 -1424 102 -648
rect 56 -1436 102 -1424
rect -46 -1483 46 -1477
rect -46 -1517 -34 -1483
rect 34 -1517 46 -1483
rect -46 -1523 46 -1517
rect -46 -1591 46 -1585
rect -46 -1625 -34 -1591
rect 34 -1625 46 -1591
rect -46 -1631 46 -1625
rect -102 -1684 -56 -1672
rect -102 -2460 -96 -1684
rect -62 -2460 -56 -1684
rect -102 -2472 -56 -2460
rect 56 -1684 102 -1672
rect 56 -2460 62 -1684
rect 96 -2460 102 -1684
rect 56 -2472 102 -2460
rect -46 -2519 46 -2513
rect -46 -2553 -34 -2519
rect 34 -2553 46 -2519
rect -46 -2559 46 -2553
<< properties >>
string FIXED_BBOX -213 -2674 213 2674
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 0.5 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
