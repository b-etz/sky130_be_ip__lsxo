magic
tech sky130A
magscale 1 2
timestamp 1712073300
<< metal3 >>
rect -5104 9132 -2732 9160
rect -5104 7108 -2816 9132
rect -2752 7108 -2732 9132
rect -5104 7080 -2732 7108
rect -2492 9132 -120 9160
rect -2492 7108 -204 9132
rect -140 7108 -120 9132
rect -2492 7080 -120 7108
rect 120 9132 2492 9160
rect 120 7108 2408 9132
rect 2472 7108 2492 9132
rect 120 7080 2492 7108
rect 2732 9132 5104 9160
rect 2732 7108 5020 9132
rect 5084 7108 5104 9132
rect 2732 7080 5104 7108
rect -5104 6812 -2732 6840
rect -5104 4788 -2816 6812
rect -2752 4788 -2732 6812
rect -5104 4760 -2732 4788
rect -2492 6812 -120 6840
rect -2492 4788 -204 6812
rect -140 4788 -120 6812
rect -2492 4760 -120 4788
rect 120 6812 2492 6840
rect 120 4788 2408 6812
rect 2472 4788 2492 6812
rect 120 4760 2492 4788
rect 2732 6812 5104 6840
rect 2732 4788 5020 6812
rect 5084 4788 5104 6812
rect 2732 4760 5104 4788
rect -5104 4492 -2732 4520
rect -5104 2468 -2816 4492
rect -2752 2468 -2732 4492
rect -5104 2440 -2732 2468
rect -2492 4492 -120 4520
rect -2492 2468 -204 4492
rect -140 2468 -120 4492
rect -2492 2440 -120 2468
rect 120 4492 2492 4520
rect 120 2468 2408 4492
rect 2472 2468 2492 4492
rect 120 2440 2492 2468
rect 2732 4492 5104 4520
rect 2732 2468 5020 4492
rect 5084 2468 5104 4492
rect 2732 2440 5104 2468
rect -5104 2172 -2732 2200
rect -5104 148 -2816 2172
rect -2752 148 -2732 2172
rect -5104 120 -2732 148
rect -2492 2172 -120 2200
rect -2492 148 -204 2172
rect -140 148 -120 2172
rect -2492 120 -120 148
rect 120 2172 2492 2200
rect 120 148 2408 2172
rect 2472 148 2492 2172
rect 120 120 2492 148
rect 2732 2172 5104 2200
rect 2732 148 5020 2172
rect 5084 148 5104 2172
rect 2732 120 5104 148
rect -5104 -148 -2732 -120
rect -5104 -2172 -2816 -148
rect -2752 -2172 -2732 -148
rect -5104 -2200 -2732 -2172
rect -2492 -148 -120 -120
rect -2492 -2172 -204 -148
rect -140 -2172 -120 -148
rect -2492 -2200 -120 -2172
rect 120 -148 2492 -120
rect 120 -2172 2408 -148
rect 2472 -2172 2492 -148
rect 120 -2200 2492 -2172
rect 2732 -148 5104 -120
rect 2732 -2172 5020 -148
rect 5084 -2172 5104 -148
rect 2732 -2200 5104 -2172
rect -5104 -2468 -2732 -2440
rect -5104 -4492 -2816 -2468
rect -2752 -4492 -2732 -2468
rect -5104 -4520 -2732 -4492
rect -2492 -2468 -120 -2440
rect -2492 -4492 -204 -2468
rect -140 -4492 -120 -2468
rect -2492 -4520 -120 -4492
rect 120 -2468 2492 -2440
rect 120 -4492 2408 -2468
rect 2472 -4492 2492 -2468
rect 120 -4520 2492 -4492
rect 2732 -2468 5104 -2440
rect 2732 -4492 5020 -2468
rect 5084 -4492 5104 -2468
rect 2732 -4520 5104 -4492
rect -5104 -4788 -2732 -4760
rect -5104 -6812 -2816 -4788
rect -2752 -6812 -2732 -4788
rect -5104 -6840 -2732 -6812
rect -2492 -4788 -120 -4760
rect -2492 -6812 -204 -4788
rect -140 -6812 -120 -4788
rect -2492 -6840 -120 -6812
rect 120 -4788 2492 -4760
rect 120 -6812 2408 -4788
rect 2472 -6812 2492 -4788
rect 120 -6840 2492 -6812
rect 2732 -4788 5104 -4760
rect 2732 -6812 5020 -4788
rect 5084 -6812 5104 -4788
rect 2732 -6840 5104 -6812
rect -5104 -7108 -2732 -7080
rect -5104 -9132 -2816 -7108
rect -2752 -9132 -2732 -7108
rect -5104 -9160 -2732 -9132
rect -2492 -7108 -120 -7080
rect -2492 -9132 -204 -7108
rect -140 -9132 -120 -7108
rect -2492 -9160 -120 -9132
rect 120 -7108 2492 -7080
rect 120 -9132 2408 -7108
rect 2472 -9132 2492 -7108
rect 120 -9160 2492 -9132
rect 2732 -7108 5104 -7080
rect 2732 -9132 5020 -7108
rect 5084 -9132 5104 -7108
rect 2732 -9160 5104 -9132
<< via3 >>
rect -2816 7108 -2752 9132
rect -204 7108 -140 9132
rect 2408 7108 2472 9132
rect 5020 7108 5084 9132
rect -2816 4788 -2752 6812
rect -204 4788 -140 6812
rect 2408 4788 2472 6812
rect 5020 4788 5084 6812
rect -2816 2468 -2752 4492
rect -204 2468 -140 4492
rect 2408 2468 2472 4492
rect 5020 2468 5084 4492
rect -2816 148 -2752 2172
rect -204 148 -140 2172
rect 2408 148 2472 2172
rect 5020 148 5084 2172
rect -2816 -2172 -2752 -148
rect -204 -2172 -140 -148
rect 2408 -2172 2472 -148
rect 5020 -2172 5084 -148
rect -2816 -4492 -2752 -2468
rect -204 -4492 -140 -2468
rect 2408 -4492 2472 -2468
rect 5020 -4492 5084 -2468
rect -2816 -6812 -2752 -4788
rect -204 -6812 -140 -4788
rect 2408 -6812 2472 -4788
rect 5020 -6812 5084 -4788
rect -2816 -9132 -2752 -7108
rect -204 -9132 -140 -7108
rect 2408 -9132 2472 -7108
rect 5020 -9132 5084 -7108
<< mimcap >>
rect -5064 9080 -3064 9120
rect -5064 7160 -5024 9080
rect -3104 7160 -3064 9080
rect -5064 7120 -3064 7160
rect -2452 9080 -452 9120
rect -2452 7160 -2412 9080
rect -492 7160 -452 9080
rect -2452 7120 -452 7160
rect 160 9080 2160 9120
rect 160 7160 200 9080
rect 2120 7160 2160 9080
rect 160 7120 2160 7160
rect 2772 9080 4772 9120
rect 2772 7160 2812 9080
rect 4732 7160 4772 9080
rect 2772 7120 4772 7160
rect -5064 6760 -3064 6800
rect -5064 4840 -5024 6760
rect -3104 4840 -3064 6760
rect -5064 4800 -3064 4840
rect -2452 6760 -452 6800
rect -2452 4840 -2412 6760
rect -492 4840 -452 6760
rect -2452 4800 -452 4840
rect 160 6760 2160 6800
rect 160 4840 200 6760
rect 2120 4840 2160 6760
rect 160 4800 2160 4840
rect 2772 6760 4772 6800
rect 2772 4840 2812 6760
rect 4732 4840 4772 6760
rect 2772 4800 4772 4840
rect -5064 4440 -3064 4480
rect -5064 2520 -5024 4440
rect -3104 2520 -3064 4440
rect -5064 2480 -3064 2520
rect -2452 4440 -452 4480
rect -2452 2520 -2412 4440
rect -492 2520 -452 4440
rect -2452 2480 -452 2520
rect 160 4440 2160 4480
rect 160 2520 200 4440
rect 2120 2520 2160 4440
rect 160 2480 2160 2520
rect 2772 4440 4772 4480
rect 2772 2520 2812 4440
rect 4732 2520 4772 4440
rect 2772 2480 4772 2520
rect -5064 2120 -3064 2160
rect -5064 200 -5024 2120
rect -3104 200 -3064 2120
rect -5064 160 -3064 200
rect -2452 2120 -452 2160
rect -2452 200 -2412 2120
rect -492 200 -452 2120
rect -2452 160 -452 200
rect 160 2120 2160 2160
rect 160 200 200 2120
rect 2120 200 2160 2120
rect 160 160 2160 200
rect 2772 2120 4772 2160
rect 2772 200 2812 2120
rect 4732 200 4772 2120
rect 2772 160 4772 200
rect -5064 -200 -3064 -160
rect -5064 -2120 -5024 -200
rect -3104 -2120 -3064 -200
rect -5064 -2160 -3064 -2120
rect -2452 -200 -452 -160
rect -2452 -2120 -2412 -200
rect -492 -2120 -452 -200
rect -2452 -2160 -452 -2120
rect 160 -200 2160 -160
rect 160 -2120 200 -200
rect 2120 -2120 2160 -200
rect 160 -2160 2160 -2120
rect 2772 -200 4772 -160
rect 2772 -2120 2812 -200
rect 4732 -2120 4772 -200
rect 2772 -2160 4772 -2120
rect -5064 -2520 -3064 -2480
rect -5064 -4440 -5024 -2520
rect -3104 -4440 -3064 -2520
rect -5064 -4480 -3064 -4440
rect -2452 -2520 -452 -2480
rect -2452 -4440 -2412 -2520
rect -492 -4440 -452 -2520
rect -2452 -4480 -452 -4440
rect 160 -2520 2160 -2480
rect 160 -4440 200 -2520
rect 2120 -4440 2160 -2520
rect 160 -4480 2160 -4440
rect 2772 -2520 4772 -2480
rect 2772 -4440 2812 -2520
rect 4732 -4440 4772 -2520
rect 2772 -4480 4772 -4440
rect -5064 -4840 -3064 -4800
rect -5064 -6760 -5024 -4840
rect -3104 -6760 -3064 -4840
rect -5064 -6800 -3064 -6760
rect -2452 -4840 -452 -4800
rect -2452 -6760 -2412 -4840
rect -492 -6760 -452 -4840
rect -2452 -6800 -452 -6760
rect 160 -4840 2160 -4800
rect 160 -6760 200 -4840
rect 2120 -6760 2160 -4840
rect 160 -6800 2160 -6760
rect 2772 -4840 4772 -4800
rect 2772 -6760 2812 -4840
rect 4732 -6760 4772 -4840
rect 2772 -6800 4772 -6760
rect -5064 -7160 -3064 -7120
rect -5064 -9080 -5024 -7160
rect -3104 -9080 -3064 -7160
rect -5064 -9120 -3064 -9080
rect -2452 -7160 -452 -7120
rect -2452 -9080 -2412 -7160
rect -492 -9080 -452 -7160
rect -2452 -9120 -452 -9080
rect 160 -7160 2160 -7120
rect 160 -9080 200 -7160
rect 2120 -9080 2160 -7160
rect 160 -9120 2160 -9080
rect 2772 -7160 4772 -7120
rect 2772 -9080 2812 -7160
rect 4732 -9080 4772 -7160
rect 2772 -9120 4772 -9080
<< mimcapcontact >>
rect -5024 7160 -3104 9080
rect -2412 7160 -492 9080
rect 200 7160 2120 9080
rect 2812 7160 4732 9080
rect -5024 4840 -3104 6760
rect -2412 4840 -492 6760
rect 200 4840 2120 6760
rect 2812 4840 4732 6760
rect -5024 2520 -3104 4440
rect -2412 2520 -492 4440
rect 200 2520 2120 4440
rect 2812 2520 4732 4440
rect -5024 200 -3104 2120
rect -2412 200 -492 2120
rect 200 200 2120 2120
rect 2812 200 4732 2120
rect -5024 -2120 -3104 -200
rect -2412 -2120 -492 -200
rect 200 -2120 2120 -200
rect 2812 -2120 4732 -200
rect -5024 -4440 -3104 -2520
rect -2412 -4440 -492 -2520
rect 200 -4440 2120 -2520
rect 2812 -4440 4732 -2520
rect -5024 -6760 -3104 -4840
rect -2412 -6760 -492 -4840
rect 200 -6760 2120 -4840
rect 2812 -6760 4732 -4840
rect -5024 -9080 -3104 -7160
rect -2412 -9080 -492 -7160
rect 200 -9080 2120 -7160
rect 2812 -9080 4732 -7160
<< metal4 >>
rect -4116 9081 -4012 9280
rect -2836 9132 -2732 9280
rect -5025 9080 -3103 9081
rect -5025 7160 -5024 9080
rect -3104 7160 -3103 9080
rect -5025 7159 -3103 7160
rect -4116 6761 -4012 7159
rect -2836 7108 -2816 9132
rect -2752 7108 -2732 9132
rect -1504 9081 -1400 9280
rect -224 9132 -120 9280
rect -2413 9080 -491 9081
rect -2413 7160 -2412 9080
rect -492 7160 -491 9080
rect -2413 7159 -491 7160
rect -2836 6812 -2732 7108
rect -5025 6760 -3103 6761
rect -5025 4840 -5024 6760
rect -3104 4840 -3103 6760
rect -5025 4839 -3103 4840
rect -4116 4441 -4012 4839
rect -2836 4788 -2816 6812
rect -2752 4788 -2732 6812
rect -1504 6761 -1400 7159
rect -224 7108 -204 9132
rect -140 7108 -120 9132
rect 1108 9081 1212 9280
rect 2388 9132 2492 9280
rect 199 9080 2121 9081
rect 199 7160 200 9080
rect 2120 7160 2121 9080
rect 199 7159 2121 7160
rect -224 6812 -120 7108
rect -2413 6760 -491 6761
rect -2413 4840 -2412 6760
rect -492 4840 -491 6760
rect -2413 4839 -491 4840
rect -2836 4492 -2732 4788
rect -5025 4440 -3103 4441
rect -5025 2520 -5024 4440
rect -3104 2520 -3103 4440
rect -5025 2519 -3103 2520
rect -4116 2121 -4012 2519
rect -2836 2468 -2816 4492
rect -2752 2468 -2732 4492
rect -1504 4441 -1400 4839
rect -224 4788 -204 6812
rect -140 4788 -120 6812
rect 1108 6761 1212 7159
rect 2388 7108 2408 9132
rect 2472 7108 2492 9132
rect 3720 9081 3824 9280
rect 5000 9132 5104 9280
rect 2811 9080 4733 9081
rect 2811 7160 2812 9080
rect 4732 7160 4733 9080
rect 2811 7159 4733 7160
rect 2388 6812 2492 7108
rect 199 6760 2121 6761
rect 199 4840 200 6760
rect 2120 4840 2121 6760
rect 199 4839 2121 4840
rect -224 4492 -120 4788
rect -2413 4440 -491 4441
rect -2413 2520 -2412 4440
rect -492 2520 -491 4440
rect -2413 2519 -491 2520
rect -2836 2172 -2732 2468
rect -5025 2120 -3103 2121
rect -5025 200 -5024 2120
rect -3104 200 -3103 2120
rect -5025 199 -3103 200
rect -4116 -199 -4012 199
rect -2836 148 -2816 2172
rect -2752 148 -2732 2172
rect -1504 2121 -1400 2519
rect -224 2468 -204 4492
rect -140 2468 -120 4492
rect 1108 4441 1212 4839
rect 2388 4788 2408 6812
rect 2472 4788 2492 6812
rect 3720 6761 3824 7159
rect 5000 7108 5020 9132
rect 5084 7108 5104 9132
rect 5000 6812 5104 7108
rect 2811 6760 4733 6761
rect 2811 4840 2812 6760
rect 4732 4840 4733 6760
rect 2811 4839 4733 4840
rect 2388 4492 2492 4788
rect 199 4440 2121 4441
rect 199 2520 200 4440
rect 2120 2520 2121 4440
rect 199 2519 2121 2520
rect -224 2172 -120 2468
rect -2413 2120 -491 2121
rect -2413 200 -2412 2120
rect -492 200 -491 2120
rect -2413 199 -491 200
rect -2836 -148 -2732 148
rect -5025 -200 -3103 -199
rect -5025 -2120 -5024 -200
rect -3104 -2120 -3103 -200
rect -5025 -2121 -3103 -2120
rect -4116 -2519 -4012 -2121
rect -2836 -2172 -2816 -148
rect -2752 -2172 -2732 -148
rect -1504 -199 -1400 199
rect -224 148 -204 2172
rect -140 148 -120 2172
rect 1108 2121 1212 2519
rect 2388 2468 2408 4492
rect 2472 2468 2492 4492
rect 3720 4441 3824 4839
rect 5000 4788 5020 6812
rect 5084 4788 5104 6812
rect 5000 4492 5104 4788
rect 2811 4440 4733 4441
rect 2811 2520 2812 4440
rect 4732 2520 4733 4440
rect 2811 2519 4733 2520
rect 2388 2172 2492 2468
rect 199 2120 2121 2121
rect 199 200 200 2120
rect 2120 200 2121 2120
rect 199 199 2121 200
rect -224 -148 -120 148
rect -2413 -200 -491 -199
rect -2413 -2120 -2412 -200
rect -492 -2120 -491 -200
rect -2413 -2121 -491 -2120
rect -2836 -2468 -2732 -2172
rect -5025 -2520 -3103 -2519
rect -5025 -4440 -5024 -2520
rect -3104 -4440 -3103 -2520
rect -5025 -4441 -3103 -4440
rect -4116 -4839 -4012 -4441
rect -2836 -4492 -2816 -2468
rect -2752 -4492 -2732 -2468
rect -1504 -2519 -1400 -2121
rect -224 -2172 -204 -148
rect -140 -2172 -120 -148
rect 1108 -199 1212 199
rect 2388 148 2408 2172
rect 2472 148 2492 2172
rect 3720 2121 3824 2519
rect 5000 2468 5020 4492
rect 5084 2468 5104 4492
rect 5000 2172 5104 2468
rect 2811 2120 4733 2121
rect 2811 200 2812 2120
rect 4732 200 4733 2120
rect 2811 199 4733 200
rect 2388 -148 2492 148
rect 199 -200 2121 -199
rect 199 -2120 200 -200
rect 2120 -2120 2121 -200
rect 199 -2121 2121 -2120
rect -224 -2468 -120 -2172
rect -2413 -2520 -491 -2519
rect -2413 -4440 -2412 -2520
rect -492 -4440 -491 -2520
rect -2413 -4441 -491 -4440
rect -2836 -4788 -2732 -4492
rect -5025 -4840 -3103 -4839
rect -5025 -6760 -5024 -4840
rect -3104 -6760 -3103 -4840
rect -5025 -6761 -3103 -6760
rect -4116 -7159 -4012 -6761
rect -2836 -6812 -2816 -4788
rect -2752 -6812 -2732 -4788
rect -1504 -4839 -1400 -4441
rect -224 -4492 -204 -2468
rect -140 -4492 -120 -2468
rect 1108 -2519 1212 -2121
rect 2388 -2172 2408 -148
rect 2472 -2172 2492 -148
rect 3720 -199 3824 199
rect 5000 148 5020 2172
rect 5084 148 5104 2172
rect 5000 -148 5104 148
rect 2811 -200 4733 -199
rect 2811 -2120 2812 -200
rect 4732 -2120 4733 -200
rect 2811 -2121 4733 -2120
rect 2388 -2468 2492 -2172
rect 199 -2520 2121 -2519
rect 199 -4440 200 -2520
rect 2120 -4440 2121 -2520
rect 199 -4441 2121 -4440
rect -224 -4788 -120 -4492
rect -2413 -4840 -491 -4839
rect -2413 -6760 -2412 -4840
rect -492 -6760 -491 -4840
rect -2413 -6761 -491 -6760
rect -2836 -7108 -2732 -6812
rect -5025 -7160 -3103 -7159
rect -5025 -9080 -5024 -7160
rect -3104 -9080 -3103 -7160
rect -5025 -9081 -3103 -9080
rect -4116 -9280 -4012 -9081
rect -2836 -9132 -2816 -7108
rect -2752 -9132 -2732 -7108
rect -1504 -7159 -1400 -6761
rect -224 -6812 -204 -4788
rect -140 -6812 -120 -4788
rect 1108 -4839 1212 -4441
rect 2388 -4492 2408 -2468
rect 2472 -4492 2492 -2468
rect 3720 -2519 3824 -2121
rect 5000 -2172 5020 -148
rect 5084 -2172 5104 -148
rect 5000 -2468 5104 -2172
rect 2811 -2520 4733 -2519
rect 2811 -4440 2812 -2520
rect 4732 -4440 4733 -2520
rect 2811 -4441 4733 -4440
rect 2388 -4788 2492 -4492
rect 199 -4840 2121 -4839
rect 199 -6760 200 -4840
rect 2120 -6760 2121 -4840
rect 199 -6761 2121 -6760
rect -224 -7108 -120 -6812
rect -2413 -7160 -491 -7159
rect -2413 -9080 -2412 -7160
rect -492 -9080 -491 -7160
rect -2413 -9081 -491 -9080
rect -2836 -9280 -2732 -9132
rect -1504 -9280 -1400 -9081
rect -224 -9132 -204 -7108
rect -140 -9132 -120 -7108
rect 1108 -7159 1212 -6761
rect 2388 -6812 2408 -4788
rect 2472 -6812 2492 -4788
rect 3720 -4839 3824 -4441
rect 5000 -4492 5020 -2468
rect 5084 -4492 5104 -2468
rect 5000 -4788 5104 -4492
rect 2811 -4840 4733 -4839
rect 2811 -6760 2812 -4840
rect 4732 -6760 4733 -4840
rect 2811 -6761 4733 -6760
rect 2388 -7108 2492 -6812
rect 199 -7160 2121 -7159
rect 199 -9080 200 -7160
rect 2120 -9080 2121 -7160
rect 199 -9081 2121 -9080
rect -224 -9280 -120 -9132
rect 1108 -9280 1212 -9081
rect 2388 -9132 2408 -7108
rect 2472 -9132 2492 -7108
rect 3720 -7159 3824 -6761
rect 5000 -6812 5020 -4788
rect 5084 -6812 5104 -4788
rect 5000 -7108 5104 -6812
rect 2811 -7160 4733 -7159
rect 2811 -9080 2812 -7160
rect 4732 -9080 4733 -7160
rect 2811 -9081 4733 -9080
rect 2388 -9280 2492 -9132
rect 3720 -9280 3824 -9081
rect 5000 -9132 5020 -7108
rect 5084 -9132 5104 -7108
rect 5000 -9280 5104 -9132
<< properties >>
string FIXED_BBOX 2732 7080 4812 9160
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 4 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
