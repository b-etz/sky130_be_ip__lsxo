magic
tech sky130A
magscale 1 2
timestamp 1712930846
<< nwell >>
rect -1825 -269 1825 269
<< pmos >>
rect -1629 -50 -29 50
rect 29 -50 1629 50
<< pdiff >>
rect -1687 38 -1629 50
rect -1687 -38 -1675 38
rect -1641 -38 -1629 38
rect -1687 -50 -1629 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 1629 38 1687 50
rect 1629 -38 1641 38
rect 1675 -38 1687 38
rect 1629 -50 1687 -38
<< pdiffc >>
rect -1675 -38 -1641 38
rect -17 -38 17 38
rect 1641 -38 1675 38
<< nsubdiff >>
rect -1789 199 -1693 233
rect 1693 199 1789 233
rect -1789 137 -1755 199
rect 1755 137 1789 199
rect -1789 -199 -1755 -137
rect 1755 -199 1789 -137
rect -1789 -233 -1693 -199
rect 1693 -233 1789 -199
<< nsubdiffcont >>
rect -1693 199 1693 233
rect -1789 -137 -1755 137
rect 1755 -137 1789 137
rect -1693 -233 1693 -199
<< poly >>
rect -1629 131 -29 147
rect -1629 97 -1613 131
rect -45 97 -29 131
rect -1629 50 -29 97
rect 29 131 1629 147
rect 29 97 45 131
rect 1613 97 1629 131
rect 29 50 1629 97
rect -1629 -97 -29 -50
rect -1629 -131 -1613 -97
rect -45 -131 -29 -97
rect -1629 -147 -29 -131
rect 29 -97 1629 -50
rect 29 -131 45 -97
rect 1613 -131 1629 -97
rect 29 -147 1629 -131
<< polycont >>
rect -1613 97 -45 131
rect 45 97 1613 131
rect -1613 -131 -45 -97
rect 45 -131 1613 -97
<< locali >>
rect -1789 199 -1693 233
rect 1693 199 1789 233
rect -1789 137 -1755 199
rect 1755 137 1789 199
rect -1629 97 -1613 131
rect -45 97 -29 131
rect 29 97 45 131
rect 1613 97 1629 131
rect -1675 38 -1641 54
rect -1675 -54 -1641 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 1641 38 1675 54
rect 1641 -54 1675 -38
rect -1629 -131 -1613 -97
rect -45 -131 -29 -97
rect 29 -131 45 -97
rect 1613 -131 1629 -97
rect -1789 -199 -1755 -137
rect 1755 -199 1789 -137
rect -1789 -233 -1693 -199
rect 1693 -233 1789 -199
<< viali >>
rect -1613 97 -45 131
rect 45 97 1613 131
rect -1675 -38 -1641 38
rect -17 -38 17 38
rect 1641 -38 1675 38
rect -1613 -131 -45 -97
rect 45 -131 1613 -97
<< metal1 >>
rect -1625 131 -33 137
rect -1625 97 -1613 131
rect -45 97 -33 131
rect -1625 91 -33 97
rect 33 131 1625 137
rect 33 97 45 131
rect 1613 97 1625 131
rect 33 91 1625 97
rect -1681 38 -1635 50
rect -1681 -38 -1675 38
rect -1641 -38 -1635 38
rect -1681 -50 -1635 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 1635 38 1681 50
rect 1635 -38 1641 38
rect 1675 -38 1681 38
rect 1635 -50 1681 -38
rect -1625 -97 -33 -91
rect -1625 -131 -1613 -97
rect -45 -131 -33 -97
rect -1625 -137 -33 -131
rect 33 -97 1625 -91
rect 33 -131 45 -97
rect 1613 -131 1625 -97
rect 33 -137 1625 -131
<< properties >>
string FIXED_BBOX -1772 -216 1772 216
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 8 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
