magic
tech sky130A
magscale 1 2
timestamp 1712854380
<< nwell >>
rect -425 -383 425 383
<< pmos >>
rect -229 64 -29 164
rect 29 64 229 164
rect -229 -164 -29 -64
rect 29 -164 229 -64
<< pdiff >>
rect -287 152 -229 164
rect -287 76 -275 152
rect -241 76 -229 152
rect -287 64 -229 76
rect -29 152 29 164
rect -29 76 -17 152
rect 17 76 29 152
rect -29 64 29 76
rect 229 152 287 164
rect 229 76 241 152
rect 275 76 287 152
rect 229 64 287 76
rect -287 -76 -229 -64
rect -287 -152 -275 -76
rect -241 -152 -229 -76
rect -287 -164 -229 -152
rect -29 -76 29 -64
rect -29 -152 -17 -76
rect 17 -152 29 -76
rect -29 -164 29 -152
rect 229 -76 287 -64
rect 229 -152 241 -76
rect 275 -152 287 -76
rect 229 -164 287 -152
<< pdiffc >>
rect -275 76 -241 152
rect -17 76 17 152
rect 241 76 275 152
rect -275 -152 -241 -76
rect -17 -152 17 -76
rect 241 -152 275 -76
<< nsubdiff >>
rect -389 313 -293 347
rect 293 313 389 347
rect -389 251 -355 313
rect 355 251 389 313
rect -389 -313 -355 -251
rect 355 -313 389 -251
rect -389 -347 -293 -313
rect 293 -347 389 -313
<< nsubdiffcont >>
rect -293 313 293 347
rect -389 -251 -355 251
rect 355 -251 389 251
rect -293 -347 293 -313
<< poly >>
rect -229 245 -29 261
rect -229 211 -213 245
rect -45 211 -29 245
rect -229 164 -29 211
rect 29 245 229 261
rect 29 211 45 245
rect 213 211 229 245
rect 29 164 229 211
rect -229 17 -29 64
rect -229 -17 -213 17
rect -45 -17 -29 17
rect -229 -64 -29 -17
rect 29 17 229 64
rect 29 -17 45 17
rect 213 -17 229 17
rect 29 -64 229 -17
rect -229 -211 -29 -164
rect -229 -245 -213 -211
rect -45 -245 -29 -211
rect -229 -261 -29 -245
rect 29 -211 229 -164
rect 29 -245 45 -211
rect 213 -245 229 -211
rect 29 -261 229 -245
<< polycont >>
rect -213 211 -45 245
rect 45 211 213 245
rect -213 -17 -45 17
rect 45 -17 213 17
rect -213 -245 -45 -211
rect 45 -245 213 -211
<< locali >>
rect -389 313 -293 347
rect 293 313 389 347
rect -389 251 -355 313
rect 355 251 389 313
rect -229 211 -213 245
rect -45 211 -29 245
rect 29 211 45 245
rect 213 211 229 245
rect -275 152 -241 168
rect -275 60 -241 76
rect -17 152 17 168
rect -17 60 17 76
rect 241 152 275 168
rect 241 60 275 76
rect -229 -17 -213 17
rect -45 -17 -29 17
rect 29 -17 45 17
rect 213 -17 229 17
rect -275 -76 -241 -60
rect -275 -168 -241 -152
rect -17 -76 17 -60
rect -17 -168 17 -152
rect 241 -76 275 -60
rect 241 -168 275 -152
rect -229 -245 -213 -211
rect -45 -245 -29 -211
rect 29 -245 45 -211
rect 213 -245 229 -211
rect -389 -313 -355 -251
rect 355 -313 389 -251
rect -389 -347 -293 -313
rect 293 -347 389 -313
<< viali >>
rect -213 211 -45 245
rect 45 211 213 245
rect -275 76 -241 152
rect -17 76 17 152
rect 241 76 275 152
rect -213 -17 -45 17
rect 45 -17 213 17
rect -275 -152 -241 -76
rect -17 -152 17 -76
rect 241 -152 275 -76
rect -213 -245 -45 -211
rect 45 -245 213 -211
<< metal1 >>
rect -225 245 -33 251
rect -225 211 -213 245
rect -45 211 -33 245
rect -225 205 -33 211
rect 33 245 225 251
rect 33 211 45 245
rect 213 211 225 245
rect 33 205 225 211
rect -281 152 -235 164
rect -281 76 -275 152
rect -241 76 -235 152
rect -281 64 -235 76
rect -23 152 23 164
rect -23 76 -17 152
rect 17 76 23 152
rect -23 64 23 76
rect 235 152 281 164
rect 235 76 241 152
rect 275 76 281 152
rect 235 64 281 76
rect -225 17 -33 23
rect -225 -17 -213 17
rect -45 -17 -33 17
rect -225 -23 -33 -17
rect 33 17 225 23
rect 33 -17 45 17
rect 213 -17 225 17
rect 33 -23 225 -17
rect -281 -76 -235 -64
rect -281 -152 -275 -76
rect -241 -152 -235 -76
rect -281 -164 -235 -152
rect -23 -76 23 -64
rect -23 -152 -17 -76
rect 17 -152 23 -76
rect -23 -164 23 -152
rect 235 -76 281 -64
rect 235 -152 241 -76
rect 275 -152 281 -76
rect 235 -164 281 -152
rect -225 -211 -33 -205
rect -225 -245 -213 -211
rect -45 -245 -33 -211
rect -225 -251 -33 -245
rect 33 -211 225 -205
rect 33 -245 45 -211
rect 213 -245 225 -211
rect 33 -251 225 -245
<< properties >>
string FIXED_BBOX -372 -330 372 330
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 1 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
