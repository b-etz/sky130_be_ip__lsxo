magic
tech sky130A
magscale 1 2
timestamp 1712854380
use sky130_fd_pr__pfet_01v8_CQSSVD  XM6
timestamp 1712071977
transform 1 0 13800 0 1 -10163
box -996 -269 996 269
use sky130_fd_pr__nfet_01v8_FMHZDY  XM7
timestamp 1712071977
transform 1 0 13798 0 1 -10738
box -996 -260 996 260
use sky130_fd_pr__pfet_01v8_CQSSVD  XM8
timestamp 1712071977
transform 1 0 11914 0 1 -10163
box -996 -269 996 269
use sky130_fd_pr__nfet_01v8_FMHZDY  XM9
timestamp 1712071977
transform 1 0 11912 0 1 -10738
box -996 -260 996 260
use sky130_fd_pr__pfet_01v8_FQSSVM  XM10
timestamp 1712071977
transform 1 0 15786 0 1 -10173
box -296 -269 296 269
use sky130_fd_pr__nfet_01v8_FMMQLY  XM11
timestamp 1712071977
transform 1 0 15772 0 1 -11240
box -296 -260 296 260
use sky130_fd_pr__pfet_01v8_3HMWVM  XM12
timestamp 1712071977
transform 1 0 16686 0 1 -10039
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_69TQ3K  XM13
timestamp 1712071977
transform 1 0 16672 0 1 -10976
box -296 -310 296 310
<< end >>
