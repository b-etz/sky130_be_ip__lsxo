magic
tech sky130A
magscale 1 2
timestamp 1713220443
<< nwell >>
rect -1145 -697 1145 697
<< mvpmos >>
rect -887 -400 -487 400
rect -429 -400 -29 400
rect 29 -400 429 400
rect 487 -400 887 400
<< mvpdiff >>
rect -945 388 -887 400
rect -945 -388 -933 388
rect -899 -388 -887 388
rect -945 -400 -887 -388
rect -487 388 -429 400
rect -487 -388 -475 388
rect -441 -388 -429 388
rect -487 -400 -429 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 429 388 487 400
rect 429 -388 441 388
rect 475 -388 487 388
rect 429 -400 487 -388
rect 887 388 945 400
rect 887 -388 899 388
rect 933 -388 945 388
rect 887 -400 945 -388
<< mvpdiffc >>
rect -933 -388 -899 388
rect -475 -388 -441 388
rect -17 -388 17 388
rect 441 -388 475 388
rect 899 -388 933 388
<< mvnsubdiff >>
rect -1079 619 1079 631
rect -1079 585 -971 619
rect 971 585 1079 619
rect -1079 573 1079 585
rect -1079 523 -1021 573
rect -1079 -523 -1067 523
rect -1033 -523 -1021 523
rect 1021 523 1079 573
rect -1079 -573 -1021 -523
rect 1021 -523 1033 523
rect 1067 -523 1079 523
rect 1021 -573 1079 -523
rect -1079 -585 1079 -573
rect -1079 -619 -971 -585
rect 971 -619 1079 -585
rect -1079 -631 1079 -619
<< mvnsubdiffcont >>
rect -971 585 971 619
rect -1067 -523 -1033 523
rect 1033 -523 1067 523
rect -971 -619 971 -585
<< poly >>
rect -887 481 -487 497
rect -887 447 -871 481
rect -503 447 -487 481
rect -887 400 -487 447
rect -429 481 -29 497
rect -429 447 -413 481
rect -45 447 -29 481
rect -429 400 -29 447
rect 29 481 429 497
rect 29 447 45 481
rect 413 447 429 481
rect 29 400 429 447
rect 487 481 887 497
rect 487 447 503 481
rect 871 447 887 481
rect 487 400 887 447
rect -887 -447 -487 -400
rect -887 -481 -871 -447
rect -503 -481 -487 -447
rect -887 -497 -487 -481
rect -429 -447 -29 -400
rect -429 -481 -413 -447
rect -45 -481 -29 -447
rect -429 -497 -29 -481
rect 29 -447 429 -400
rect 29 -481 45 -447
rect 413 -481 429 -447
rect 29 -497 429 -481
rect 487 -447 887 -400
rect 487 -481 503 -447
rect 871 -481 887 -447
rect 487 -497 887 -481
<< polycont >>
rect -871 447 -503 481
rect -413 447 -45 481
rect 45 447 413 481
rect 503 447 871 481
rect -871 -481 -503 -447
rect -413 -481 -45 -447
rect 45 -481 413 -447
rect 503 -481 871 -447
<< locali >>
rect -1067 585 -971 619
rect 971 585 1067 619
rect -1067 523 -1033 585
rect 1033 523 1067 585
rect -887 447 -871 481
rect -503 447 -487 481
rect -429 447 -413 481
rect -45 447 -29 481
rect 29 447 45 481
rect 413 447 429 481
rect 487 447 503 481
rect 871 447 887 481
rect -933 388 -899 404
rect -933 -404 -899 -388
rect -475 388 -441 404
rect -475 -404 -441 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 441 388 475 404
rect 441 -404 475 -388
rect 899 388 933 404
rect 899 -404 933 -388
rect -887 -481 -871 -447
rect -503 -481 -487 -447
rect -429 -481 -413 -447
rect -45 -481 -29 -447
rect 29 -481 45 -447
rect 413 -481 429 -447
rect 487 -481 503 -447
rect 871 -481 887 -447
rect -1067 -585 -1033 -523
rect 1033 -585 1067 -523
rect -1067 -619 -971 -585
rect 971 -619 1067 -585
<< properties >>
string FIXED_BBOX -1050 -602 1050 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 2 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 0 viadrn 0 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
