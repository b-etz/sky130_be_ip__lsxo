magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< metal3 >>
rect -1186 13772 1186 13800
rect -1186 11748 1102 13772
rect 1166 11748 1186 13772
rect -1186 11720 1186 11748
rect -1186 11452 1186 11480
rect -1186 9428 1102 11452
rect 1166 9428 1186 11452
rect -1186 9400 1186 9428
rect -1186 9132 1186 9160
rect -1186 7108 1102 9132
rect 1166 7108 1186 9132
rect -1186 7080 1186 7108
rect -1186 6812 1186 6840
rect -1186 4788 1102 6812
rect 1166 4788 1186 6812
rect -1186 4760 1186 4788
rect -1186 4492 1186 4520
rect -1186 2468 1102 4492
rect 1166 2468 1186 4492
rect -1186 2440 1186 2468
rect -1186 2172 1186 2200
rect -1186 148 1102 2172
rect 1166 148 1186 2172
rect -1186 120 1186 148
rect -1186 -148 1186 -120
rect -1186 -2172 1102 -148
rect 1166 -2172 1186 -148
rect -1186 -2200 1186 -2172
rect -1186 -2468 1186 -2440
rect -1186 -4492 1102 -2468
rect 1166 -4492 1186 -2468
rect -1186 -4520 1186 -4492
rect -1186 -4788 1186 -4760
rect -1186 -6812 1102 -4788
rect 1166 -6812 1186 -4788
rect -1186 -6840 1186 -6812
rect -1186 -7108 1186 -7080
rect -1186 -9132 1102 -7108
rect 1166 -9132 1186 -7108
rect -1186 -9160 1186 -9132
rect -1186 -9428 1186 -9400
rect -1186 -11452 1102 -9428
rect 1166 -11452 1186 -9428
rect -1186 -11480 1186 -11452
rect -1186 -11748 1186 -11720
rect -1186 -13772 1102 -11748
rect 1166 -13772 1186 -11748
rect -1186 -13800 1186 -13772
<< via3 >>
rect 1102 11748 1166 13772
rect 1102 9428 1166 11452
rect 1102 7108 1166 9132
rect 1102 4788 1166 6812
rect 1102 2468 1166 4492
rect 1102 148 1166 2172
rect 1102 -2172 1166 -148
rect 1102 -4492 1166 -2468
rect 1102 -6812 1166 -4788
rect 1102 -9132 1166 -7108
rect 1102 -11452 1166 -9428
rect 1102 -13772 1166 -11748
<< mimcap >>
rect -1146 13720 854 13760
rect -1146 11800 -1106 13720
rect 814 11800 854 13720
rect -1146 11760 854 11800
rect -1146 11400 854 11440
rect -1146 9480 -1106 11400
rect 814 9480 854 11400
rect -1146 9440 854 9480
rect -1146 9080 854 9120
rect -1146 7160 -1106 9080
rect 814 7160 854 9080
rect -1146 7120 854 7160
rect -1146 6760 854 6800
rect -1146 4840 -1106 6760
rect 814 4840 854 6760
rect -1146 4800 854 4840
rect -1146 4440 854 4480
rect -1146 2520 -1106 4440
rect 814 2520 854 4440
rect -1146 2480 854 2520
rect -1146 2120 854 2160
rect -1146 200 -1106 2120
rect 814 200 854 2120
rect -1146 160 854 200
rect -1146 -200 854 -160
rect -1146 -2120 -1106 -200
rect 814 -2120 854 -200
rect -1146 -2160 854 -2120
rect -1146 -2520 854 -2480
rect -1146 -4440 -1106 -2520
rect 814 -4440 854 -2520
rect -1146 -4480 854 -4440
rect -1146 -4840 854 -4800
rect -1146 -6760 -1106 -4840
rect 814 -6760 854 -4840
rect -1146 -6800 854 -6760
rect -1146 -7160 854 -7120
rect -1146 -9080 -1106 -7160
rect 814 -9080 854 -7160
rect -1146 -9120 854 -9080
rect -1146 -9480 854 -9440
rect -1146 -11400 -1106 -9480
rect 814 -11400 854 -9480
rect -1146 -11440 854 -11400
rect -1146 -11800 854 -11760
rect -1146 -13720 -1106 -11800
rect 814 -13720 854 -11800
rect -1146 -13760 854 -13720
<< mimcapcontact >>
rect -1106 11800 814 13720
rect -1106 9480 814 11400
rect -1106 7160 814 9080
rect -1106 4840 814 6760
rect -1106 2520 814 4440
rect -1106 200 814 2120
rect -1106 -2120 814 -200
rect -1106 -4440 814 -2520
rect -1106 -6760 814 -4840
rect -1106 -9080 814 -7160
rect -1106 -11400 814 -9480
rect -1106 -13720 814 -11800
<< metal4 >>
rect -198 13721 -94 13920
rect 1082 13772 1186 13920
rect -1107 13720 815 13721
rect -1107 11800 -1106 13720
rect 814 11800 815 13720
rect -1107 11799 815 11800
rect -198 11401 -94 11799
rect 1082 11748 1102 13772
rect 1166 11748 1186 13772
rect 1082 11452 1186 11748
rect -1107 11400 815 11401
rect -1107 9480 -1106 11400
rect 814 9480 815 11400
rect -1107 9479 815 9480
rect -198 9081 -94 9479
rect 1082 9428 1102 11452
rect 1166 9428 1186 11452
rect 1082 9132 1186 9428
rect -1107 9080 815 9081
rect -1107 7160 -1106 9080
rect 814 7160 815 9080
rect -1107 7159 815 7160
rect -198 6761 -94 7159
rect 1082 7108 1102 9132
rect 1166 7108 1186 9132
rect 1082 6812 1186 7108
rect -1107 6760 815 6761
rect -1107 4840 -1106 6760
rect 814 4840 815 6760
rect -1107 4839 815 4840
rect -198 4441 -94 4839
rect 1082 4788 1102 6812
rect 1166 4788 1186 6812
rect 1082 4492 1186 4788
rect -1107 4440 815 4441
rect -1107 2520 -1106 4440
rect 814 2520 815 4440
rect -1107 2519 815 2520
rect -198 2121 -94 2519
rect 1082 2468 1102 4492
rect 1166 2468 1186 4492
rect 1082 2172 1186 2468
rect -1107 2120 815 2121
rect -1107 200 -1106 2120
rect 814 200 815 2120
rect -1107 199 815 200
rect -198 -199 -94 199
rect 1082 148 1102 2172
rect 1166 148 1186 2172
rect 1082 -148 1186 148
rect -1107 -200 815 -199
rect -1107 -2120 -1106 -200
rect 814 -2120 815 -200
rect -1107 -2121 815 -2120
rect -198 -2519 -94 -2121
rect 1082 -2172 1102 -148
rect 1166 -2172 1186 -148
rect 1082 -2468 1186 -2172
rect -1107 -2520 815 -2519
rect -1107 -4440 -1106 -2520
rect 814 -4440 815 -2520
rect -1107 -4441 815 -4440
rect -198 -4839 -94 -4441
rect 1082 -4492 1102 -2468
rect 1166 -4492 1186 -2468
rect 1082 -4788 1186 -4492
rect -1107 -4840 815 -4839
rect -1107 -6760 -1106 -4840
rect 814 -6760 815 -4840
rect -1107 -6761 815 -6760
rect -198 -7159 -94 -6761
rect 1082 -6812 1102 -4788
rect 1166 -6812 1186 -4788
rect 1082 -7108 1186 -6812
rect -1107 -7160 815 -7159
rect -1107 -9080 -1106 -7160
rect 814 -9080 815 -7160
rect -1107 -9081 815 -9080
rect -198 -9479 -94 -9081
rect 1082 -9132 1102 -7108
rect 1166 -9132 1186 -7108
rect 1082 -9428 1186 -9132
rect -1107 -9480 815 -9479
rect -1107 -11400 -1106 -9480
rect 814 -11400 815 -9480
rect -1107 -11401 815 -11400
rect -198 -11799 -94 -11401
rect 1082 -11452 1102 -9428
rect 1166 -11452 1186 -9428
rect 1082 -11748 1186 -11452
rect -1107 -11800 815 -11799
rect -1107 -13720 -1106 -11800
rect 814 -13720 815 -11800
rect -1107 -13721 815 -13720
rect -198 -13920 -94 -13721
rect 1082 -13772 1102 -11748
rect 1166 -13772 1186 -11748
rect 1082 -13920 1186 -13772
<< properties >>
string FIXED_BBOX -1186 11720 894 13800
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 12 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
