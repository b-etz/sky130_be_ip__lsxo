magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< metal3 >>
rect -3798 4492 -1426 4520
rect -3798 2468 -1510 4492
rect -1446 2468 -1426 4492
rect -3798 2440 -1426 2468
rect -1186 4492 1186 4520
rect -1186 2468 1102 4492
rect 1166 2468 1186 4492
rect -1186 2440 1186 2468
rect 1426 4492 3798 4520
rect 1426 2468 3714 4492
rect 3778 2468 3798 4492
rect 1426 2440 3798 2468
rect -3798 2172 -1426 2200
rect -3798 148 -1510 2172
rect -1446 148 -1426 2172
rect -3798 120 -1426 148
rect -1186 2172 1186 2200
rect -1186 148 1102 2172
rect 1166 148 1186 2172
rect -1186 120 1186 148
rect 1426 2172 3798 2200
rect 1426 148 3714 2172
rect 3778 148 3798 2172
rect 1426 120 3798 148
rect -3798 -148 -1426 -120
rect -3798 -2172 -1510 -148
rect -1446 -2172 -1426 -148
rect -3798 -2200 -1426 -2172
rect -1186 -148 1186 -120
rect -1186 -2172 1102 -148
rect 1166 -2172 1186 -148
rect -1186 -2200 1186 -2172
rect 1426 -148 3798 -120
rect 1426 -2172 3714 -148
rect 3778 -2172 3798 -148
rect 1426 -2200 3798 -2172
rect -3798 -2468 -1426 -2440
rect -3798 -4492 -1510 -2468
rect -1446 -4492 -1426 -2468
rect -3798 -4520 -1426 -4492
rect -1186 -2468 1186 -2440
rect -1186 -4492 1102 -2468
rect 1166 -4492 1186 -2468
rect -1186 -4520 1186 -4492
rect 1426 -2468 3798 -2440
rect 1426 -4492 3714 -2468
rect 3778 -4492 3798 -2468
rect 1426 -4520 3798 -4492
<< via3 >>
rect -1510 2468 -1446 4492
rect 1102 2468 1166 4492
rect 3714 2468 3778 4492
rect -1510 148 -1446 2172
rect 1102 148 1166 2172
rect 3714 148 3778 2172
rect -1510 -2172 -1446 -148
rect 1102 -2172 1166 -148
rect 3714 -2172 3778 -148
rect -1510 -4492 -1446 -2468
rect 1102 -4492 1166 -2468
rect 3714 -4492 3778 -2468
<< mimcap >>
rect -3758 4440 -1758 4480
rect -3758 2520 -3718 4440
rect -1798 2520 -1758 4440
rect -3758 2480 -1758 2520
rect -1146 4440 854 4480
rect -1146 2520 -1106 4440
rect 814 2520 854 4440
rect -1146 2480 854 2520
rect 1466 4440 3466 4480
rect 1466 2520 1506 4440
rect 3426 2520 3466 4440
rect 1466 2480 3466 2520
rect -3758 2120 -1758 2160
rect -3758 200 -3718 2120
rect -1798 200 -1758 2120
rect -3758 160 -1758 200
rect -1146 2120 854 2160
rect -1146 200 -1106 2120
rect 814 200 854 2120
rect -1146 160 854 200
rect 1466 2120 3466 2160
rect 1466 200 1506 2120
rect 3426 200 3466 2120
rect 1466 160 3466 200
rect -3758 -200 -1758 -160
rect -3758 -2120 -3718 -200
rect -1798 -2120 -1758 -200
rect -3758 -2160 -1758 -2120
rect -1146 -200 854 -160
rect -1146 -2120 -1106 -200
rect 814 -2120 854 -200
rect -1146 -2160 854 -2120
rect 1466 -200 3466 -160
rect 1466 -2120 1506 -200
rect 3426 -2120 3466 -200
rect 1466 -2160 3466 -2120
rect -3758 -2520 -1758 -2480
rect -3758 -4440 -3718 -2520
rect -1798 -4440 -1758 -2520
rect -3758 -4480 -1758 -4440
rect -1146 -2520 854 -2480
rect -1146 -4440 -1106 -2520
rect 814 -4440 854 -2520
rect -1146 -4480 854 -4440
rect 1466 -2520 3466 -2480
rect 1466 -4440 1506 -2520
rect 3426 -4440 3466 -2520
rect 1466 -4480 3466 -4440
<< mimcapcontact >>
rect -3718 2520 -1798 4440
rect -1106 2520 814 4440
rect 1506 2520 3426 4440
rect -3718 200 -1798 2120
rect -1106 200 814 2120
rect 1506 200 3426 2120
rect -3718 -2120 -1798 -200
rect -1106 -2120 814 -200
rect 1506 -2120 3426 -200
rect -3718 -4440 -1798 -2520
rect -1106 -4440 814 -2520
rect 1506 -4440 3426 -2520
<< metal4 >>
rect -2810 4441 -2706 4640
rect -1530 4492 -1426 4640
rect -3719 4440 -1797 4441
rect -3719 2520 -3718 4440
rect -1798 2520 -1797 4440
rect -3719 2519 -1797 2520
rect -2810 2121 -2706 2519
rect -1530 2468 -1510 4492
rect -1446 2468 -1426 4492
rect -198 4441 -94 4640
rect 1082 4492 1186 4640
rect -1107 4440 815 4441
rect -1107 2520 -1106 4440
rect 814 2520 815 4440
rect -1107 2519 815 2520
rect -1530 2172 -1426 2468
rect -3719 2120 -1797 2121
rect -3719 200 -3718 2120
rect -1798 200 -1797 2120
rect -3719 199 -1797 200
rect -2810 -199 -2706 199
rect -1530 148 -1510 2172
rect -1446 148 -1426 2172
rect -198 2121 -94 2519
rect 1082 2468 1102 4492
rect 1166 2468 1186 4492
rect 2414 4441 2518 4640
rect 3694 4492 3798 4640
rect 1505 4440 3427 4441
rect 1505 2520 1506 4440
rect 3426 2520 3427 4440
rect 1505 2519 3427 2520
rect 1082 2172 1186 2468
rect -1107 2120 815 2121
rect -1107 200 -1106 2120
rect 814 200 815 2120
rect -1107 199 815 200
rect -1530 -148 -1426 148
rect -3719 -200 -1797 -199
rect -3719 -2120 -3718 -200
rect -1798 -2120 -1797 -200
rect -3719 -2121 -1797 -2120
rect -2810 -2519 -2706 -2121
rect -1530 -2172 -1510 -148
rect -1446 -2172 -1426 -148
rect -198 -199 -94 199
rect 1082 148 1102 2172
rect 1166 148 1186 2172
rect 2414 2121 2518 2519
rect 3694 2468 3714 4492
rect 3778 2468 3798 4492
rect 3694 2172 3798 2468
rect 1505 2120 3427 2121
rect 1505 200 1506 2120
rect 3426 200 3427 2120
rect 1505 199 3427 200
rect 1082 -148 1186 148
rect -1107 -200 815 -199
rect -1107 -2120 -1106 -200
rect 814 -2120 815 -200
rect -1107 -2121 815 -2120
rect -1530 -2468 -1426 -2172
rect -3719 -2520 -1797 -2519
rect -3719 -4440 -3718 -2520
rect -1798 -4440 -1797 -2520
rect -3719 -4441 -1797 -4440
rect -2810 -4640 -2706 -4441
rect -1530 -4492 -1510 -2468
rect -1446 -4492 -1426 -2468
rect -198 -2519 -94 -2121
rect 1082 -2172 1102 -148
rect 1166 -2172 1186 -148
rect 2414 -199 2518 199
rect 3694 148 3714 2172
rect 3778 148 3798 2172
rect 3694 -148 3798 148
rect 1505 -200 3427 -199
rect 1505 -2120 1506 -200
rect 3426 -2120 3427 -200
rect 1505 -2121 3427 -2120
rect 1082 -2468 1186 -2172
rect -1107 -2520 815 -2519
rect -1107 -4440 -1106 -2520
rect 814 -4440 815 -2520
rect -1107 -4441 815 -4440
rect -1530 -4640 -1426 -4492
rect -198 -4640 -94 -4441
rect 1082 -4492 1102 -2468
rect 1166 -4492 1186 -2468
rect 2414 -2519 2518 -2121
rect 3694 -2172 3714 -148
rect 3778 -2172 3798 -148
rect 3694 -2468 3798 -2172
rect 1505 -2520 3427 -2519
rect 1505 -4440 1506 -2520
rect 3426 -4440 3427 -2520
rect 1505 -4441 3427 -4440
rect 1082 -4640 1186 -4492
rect 2414 -4640 2518 -4441
rect 3694 -4492 3714 -2468
rect 3778 -4492 3798 -2468
rect 3694 -4640 3798 -4492
<< properties >>
string FIXED_BBOX 1426 2440 3506 4520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 3 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
