magic
tech sky130A
magscale 1 2
timestamp 1712854380
<< pwell >>
rect -2031 -458 2031 458
<< mvnmos >>
rect -1803 -200 -1403 200
rect -1345 -200 -945 200
rect -887 -200 -487 200
rect -429 -200 -29 200
rect 29 -200 429 200
rect 487 -200 887 200
rect 945 -200 1345 200
rect 1403 -200 1803 200
<< mvndiff >>
rect -1861 188 -1803 200
rect -1861 -188 -1849 188
rect -1815 -188 -1803 188
rect -1861 -200 -1803 -188
rect -1403 188 -1345 200
rect -1403 -188 -1391 188
rect -1357 -188 -1345 188
rect -1403 -200 -1345 -188
rect -945 188 -887 200
rect -945 -188 -933 188
rect -899 -188 -887 188
rect -945 -200 -887 -188
rect -487 188 -429 200
rect -487 -188 -475 188
rect -441 -188 -429 188
rect -487 -200 -429 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 429 188 487 200
rect 429 -188 441 188
rect 475 -188 487 188
rect 429 -200 487 -188
rect 887 188 945 200
rect 887 -188 899 188
rect 933 -188 945 188
rect 887 -200 945 -188
rect 1345 188 1403 200
rect 1345 -188 1357 188
rect 1391 -188 1403 188
rect 1345 -200 1403 -188
rect 1803 188 1861 200
rect 1803 -188 1815 188
rect 1849 -188 1861 188
rect 1803 -200 1861 -188
<< mvndiffc >>
rect -1849 -188 -1815 188
rect -1391 -188 -1357 188
rect -933 -188 -899 188
rect -475 -188 -441 188
rect -17 -188 17 188
rect 441 -188 475 188
rect 899 -188 933 188
rect 1357 -188 1391 188
rect 1815 -188 1849 188
<< mvpsubdiff >>
rect -1995 410 1995 422
rect -1995 376 -1887 410
rect 1887 376 1995 410
rect -1995 364 1995 376
rect -1995 314 -1937 364
rect -1995 -314 -1983 314
rect -1949 -314 -1937 314
rect 1937 314 1995 364
rect -1995 -364 -1937 -314
rect 1937 -314 1949 314
rect 1983 -314 1995 314
rect 1937 -364 1995 -314
rect -1995 -376 1995 -364
rect -1995 -410 -1887 -376
rect 1887 -410 1995 -376
rect -1995 -422 1995 -410
<< mvpsubdiffcont >>
rect -1887 376 1887 410
rect -1983 -314 -1949 314
rect 1949 -314 1983 314
rect -1887 -410 1887 -376
<< poly >>
rect -1803 272 -1403 288
rect -1803 238 -1787 272
rect -1419 238 -1403 272
rect -1803 200 -1403 238
rect -1345 272 -945 288
rect -1345 238 -1329 272
rect -961 238 -945 272
rect -1345 200 -945 238
rect -887 272 -487 288
rect -887 238 -871 272
rect -503 238 -487 272
rect -887 200 -487 238
rect -429 272 -29 288
rect -429 238 -413 272
rect -45 238 -29 272
rect -429 200 -29 238
rect 29 272 429 288
rect 29 238 45 272
rect 413 238 429 272
rect 29 200 429 238
rect 487 272 887 288
rect 487 238 503 272
rect 871 238 887 272
rect 487 200 887 238
rect 945 272 1345 288
rect 945 238 961 272
rect 1329 238 1345 272
rect 945 200 1345 238
rect 1403 272 1803 288
rect 1403 238 1419 272
rect 1787 238 1803 272
rect 1403 200 1803 238
rect -1803 -238 -1403 -200
rect -1803 -272 -1787 -238
rect -1419 -272 -1403 -238
rect -1803 -288 -1403 -272
rect -1345 -238 -945 -200
rect -1345 -272 -1329 -238
rect -961 -272 -945 -238
rect -1345 -288 -945 -272
rect -887 -238 -487 -200
rect -887 -272 -871 -238
rect -503 -272 -487 -238
rect -887 -288 -487 -272
rect -429 -238 -29 -200
rect -429 -272 -413 -238
rect -45 -272 -29 -238
rect -429 -288 -29 -272
rect 29 -238 429 -200
rect 29 -272 45 -238
rect 413 -272 429 -238
rect 29 -288 429 -272
rect 487 -238 887 -200
rect 487 -272 503 -238
rect 871 -272 887 -238
rect 487 -288 887 -272
rect 945 -238 1345 -200
rect 945 -272 961 -238
rect 1329 -272 1345 -238
rect 945 -288 1345 -272
rect 1403 -238 1803 -200
rect 1403 -272 1419 -238
rect 1787 -272 1803 -238
rect 1403 -288 1803 -272
<< polycont >>
rect -1787 238 -1419 272
rect -1329 238 -961 272
rect -871 238 -503 272
rect -413 238 -45 272
rect 45 238 413 272
rect 503 238 871 272
rect 961 238 1329 272
rect 1419 238 1787 272
rect -1787 -272 -1419 -238
rect -1329 -272 -961 -238
rect -871 -272 -503 -238
rect -413 -272 -45 -238
rect 45 -272 413 -238
rect 503 -272 871 -238
rect 961 -272 1329 -238
rect 1419 -272 1787 -238
<< locali >>
rect -1983 376 -1887 410
rect 1887 376 1983 410
rect -1983 314 -1949 376
rect 1949 314 1983 376
rect -1803 238 -1787 272
rect -1419 238 -1403 272
rect -1345 238 -1329 272
rect -961 238 -945 272
rect -887 238 -871 272
rect -503 238 -487 272
rect -429 238 -413 272
rect -45 238 -29 272
rect 29 238 45 272
rect 413 238 429 272
rect 487 238 503 272
rect 871 238 887 272
rect 945 238 961 272
rect 1329 238 1345 272
rect 1403 238 1419 272
rect 1787 238 1803 272
rect -1849 188 -1815 204
rect -1849 -204 -1815 -188
rect -1391 188 -1357 204
rect -1391 -204 -1357 -188
rect -933 188 -899 204
rect -933 -204 -899 -188
rect -475 188 -441 204
rect -475 -204 -441 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 441 188 475 204
rect 441 -204 475 -188
rect 899 188 933 204
rect 899 -204 933 -188
rect 1357 188 1391 204
rect 1357 -204 1391 -188
rect 1815 188 1849 204
rect 1815 -204 1849 -188
rect -1803 -272 -1787 -238
rect -1419 -272 -1403 -238
rect -1345 -272 -1329 -238
rect -961 -272 -945 -238
rect -887 -272 -871 -238
rect -503 -272 -487 -238
rect -429 -272 -413 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 413 -272 429 -238
rect 487 -272 503 -238
rect 871 -272 887 -238
rect 945 -272 961 -238
rect 1329 -272 1345 -238
rect 1403 -272 1419 -238
rect 1787 -272 1803 -238
rect -1983 -376 -1949 -314
rect 1949 -376 1983 -314
rect -1983 -410 -1887 -376
rect 1887 -410 1983 -376
<< viali >>
rect -1787 238 -1419 272
rect -1329 238 -961 272
rect -871 238 -503 272
rect -413 238 -45 272
rect 45 238 413 272
rect 503 238 871 272
rect 961 238 1329 272
rect 1419 238 1787 272
rect -1849 -188 -1815 188
rect -1391 -188 -1357 188
rect -933 -188 -899 188
rect -475 -188 -441 188
rect -17 -188 17 188
rect 441 -188 475 188
rect 899 -188 933 188
rect 1357 -188 1391 188
rect 1815 -188 1849 188
rect -1787 -272 -1419 -238
rect -1329 -272 -961 -238
rect -871 -272 -503 -238
rect -413 -272 -45 -238
rect 45 -272 413 -238
rect 503 -272 871 -238
rect 961 -272 1329 -238
rect 1419 -272 1787 -238
<< metal1 >>
rect -1799 272 -1407 278
rect -1799 238 -1787 272
rect -1419 238 -1407 272
rect -1799 232 -1407 238
rect -1341 272 -949 278
rect -1341 238 -1329 272
rect -961 238 -949 272
rect -1341 232 -949 238
rect -883 272 -491 278
rect -883 238 -871 272
rect -503 238 -491 272
rect -883 232 -491 238
rect -425 272 -33 278
rect -425 238 -413 272
rect -45 238 -33 272
rect -425 232 -33 238
rect 33 272 425 278
rect 33 238 45 272
rect 413 238 425 272
rect 33 232 425 238
rect 491 272 883 278
rect 491 238 503 272
rect 871 238 883 272
rect 491 232 883 238
rect 949 272 1341 278
rect 949 238 961 272
rect 1329 238 1341 272
rect 949 232 1341 238
rect 1407 272 1799 278
rect 1407 238 1419 272
rect 1787 238 1799 272
rect 1407 232 1799 238
rect -1855 188 -1809 200
rect -1855 -188 -1849 188
rect -1815 -188 -1809 188
rect -1855 -200 -1809 -188
rect -1397 188 -1351 200
rect -1397 -188 -1391 188
rect -1357 -188 -1351 188
rect -1397 -200 -1351 -188
rect -939 188 -893 200
rect -939 -188 -933 188
rect -899 -188 -893 188
rect -939 -200 -893 -188
rect -481 188 -435 200
rect -481 -188 -475 188
rect -441 -188 -435 188
rect -481 -200 -435 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 435 188 481 200
rect 435 -188 441 188
rect 475 -188 481 188
rect 435 -200 481 -188
rect 893 188 939 200
rect 893 -188 899 188
rect 933 -188 939 188
rect 893 -200 939 -188
rect 1351 188 1397 200
rect 1351 -188 1357 188
rect 1391 -188 1397 188
rect 1351 -200 1397 -188
rect 1809 188 1855 200
rect 1809 -188 1815 188
rect 1849 -188 1855 188
rect 1809 -200 1855 -188
rect -1799 -238 -1407 -232
rect -1799 -272 -1787 -238
rect -1419 -272 -1407 -238
rect -1799 -278 -1407 -272
rect -1341 -238 -949 -232
rect -1341 -272 -1329 -238
rect -961 -272 -949 -238
rect -1341 -278 -949 -272
rect -883 -238 -491 -232
rect -883 -272 -871 -238
rect -503 -272 -491 -238
rect -883 -278 -491 -272
rect -425 -238 -33 -232
rect -425 -272 -413 -238
rect -45 -272 -33 -238
rect -425 -278 -33 -272
rect 33 -238 425 -232
rect 33 -272 45 -238
rect 413 -272 425 -238
rect 33 -278 425 -272
rect 491 -238 883 -232
rect 491 -272 503 -238
rect 871 -272 883 -238
rect 491 -278 883 -272
rect 949 -238 1341 -232
rect 949 -272 961 -238
rect 1329 -272 1341 -238
rect 949 -278 1341 -272
rect 1407 -238 1799 -232
rect 1407 -272 1419 -238
rect 1787 -272 1799 -238
rect 1407 -278 1799 -272
<< properties >>
string FIXED_BBOX -1966 -393 1966 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 2 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
