magic
tech sky130A
magscale 1 2
timestamp 1712544943
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 3364 -7142 3370 -6962
rect 2500 -7222 3370 -7142
rect 3478 -7222 3484 -6962
rect 3614 -7214 3620 -6954
rect 3728 -7134 3734 -6954
rect 3728 -7214 4600 -7134
rect 2406 -8054 2412 -7254
rect 2520 -8054 2526 -7254
rect 2564 -8054 2570 -7254
rect 2678 -8054 2684 -7254
rect 2722 -8054 2728 -7254
rect 2836 -8054 2842 -7254
rect 2880 -8054 2886 -7254
rect 2994 -8054 3000 -7254
rect 3036 -8054 3042 -7254
rect 3150 -8054 3156 -7254
rect 3196 -8054 3202 -7254
rect 3310 -8054 3316 -7254
rect 3364 -8086 3370 -7906
rect 2500 -8166 3370 -8086
rect 3478 -8086 3484 -7906
rect 3478 -8166 3486 -8086
rect 3614 -8176 3620 -7916
rect 3728 -8096 3734 -7916
rect 3782 -8054 3790 -7254
rect 3894 -8054 3902 -7254
rect 3940 -8054 3946 -7254
rect 4054 -8054 4060 -7254
rect 4098 -8054 4104 -7254
rect 4212 -8054 4218 -7254
rect 4256 -8054 4262 -7254
rect 4370 -8054 4376 -7254
rect 4414 -8054 4420 -7254
rect 4528 -8054 4534 -7254
rect 4572 -8054 4578 -7254
rect 4686 -8054 4692 -7254
rect 3728 -8176 4600 -8096
<< via1 >>
rect 3370 -7222 3478 -6962
rect 3620 -7214 3728 -6954
rect 2412 -8054 2520 -7254
rect 2570 -8054 2678 -7254
rect 2728 -8054 2836 -7254
rect 2886 -8054 2994 -7254
rect 3042 -8054 3150 -7254
rect 3202 -8054 3310 -7254
rect 3370 -8166 3478 -7906
rect 3620 -8176 3728 -7916
rect 3790 -8054 3894 -7254
rect 3946 -8054 4054 -7254
rect 4104 -8054 4212 -7254
rect 4262 -8054 4370 -7254
rect 4420 -8054 4528 -7254
rect 4578 -8054 4686 -7254
<< metal2 >>
rect 2610 -6860 3484 -6740
rect 3364 -6962 3484 -6860
rect 2406 -7174 3158 -6974
rect 2406 -7254 2526 -7174
rect 2722 -7254 2842 -7174
rect 3036 -7254 3158 -7174
rect 3364 -7222 3370 -6962
rect 3478 -7222 3484 -6962
rect 2406 -8054 2412 -7254
rect 2520 -8054 2526 -7254
rect 2564 -8054 2570 -7254
rect 2678 -8054 2684 -7254
rect 2722 -8054 2728 -7254
rect 2836 -8054 2842 -7254
rect 2880 -8054 2886 -7254
rect 2994 -8054 3000 -7254
rect 3036 -8054 3042 -7254
rect 3150 -7554 3158 -7254
rect 3150 -8054 3156 -7554
rect 3196 -8054 3202 -7254
rect 3310 -8054 3316 -7254
rect 2564 -8134 2684 -8054
rect 2880 -8134 3000 -8054
rect 3196 -8134 3316 -8054
rect 2564 -8334 3316 -8134
rect 3364 -7906 3484 -7222
rect 3364 -8166 3370 -7906
rect 3478 -8166 3484 -7906
rect 3614 -6954 3734 -6750
rect 3614 -7214 3620 -6954
rect 3728 -7214 3734 -6954
rect 3614 -7916 3734 -7214
rect 3940 -7174 4692 -6974
rect 3940 -7254 4060 -7174
rect 4256 -7254 4376 -7174
rect 4572 -7254 4692 -7174
rect 3614 -8176 3620 -7916
rect 3728 -8176 3734 -7916
rect 3782 -8054 3790 -7254
rect 3894 -8054 3902 -7254
rect 3940 -8054 3946 -7254
rect 4054 -8054 4060 -7254
rect 4098 -8054 4104 -7254
rect 4212 -8054 4218 -7254
rect 4256 -8054 4262 -7254
rect 4370 -8054 4376 -7254
rect 4414 -8054 4420 -7254
rect 4528 -8054 4534 -7254
rect 4572 -8054 4578 -7254
rect 4686 -8054 4692 -7254
rect 3782 -8134 3902 -8054
rect 4098 -8134 4218 -8054
rect 4414 -8134 4534 -8054
rect 3782 -8334 4534 -8134
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 0 1 2848 -1 0 -1286
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x2
timestamp 1707688321
transform 0 -1 5492 -1 0 -1286
box -38 -48 314 592
use level_shift  x3
timestamp 1712539951
transform 0 1 4250 -1 0 -1190
box 652 -1950 5670 -128
use level_shift  x4
timestamp 1712539951
transform 0 -1 4086 -1 0 -1190
box 652 -1950 5670 -128
use bias_gen  x5
timestamp 1712250795
transform 1 0 1962 0 1 -15524
box -450 -14480 16732 3256
use dout_amp  x6
timestamp 1712087189
transform 1 0 20214 0 1 -2274
box -1220 -12900 16982 200
use ripl_dly_clk_buf  x7
timestamp 1712544943
transform 1 0 38260 0 1 -6068
box 872 -3046 9184 598
use sky130_fd_pr__cap_mim_m3_1_KAF84V  XC1
timestamp 1712073300
transform -1 0 17850 0 -1 -24526
box -886 -3440 886 3440
use sky130_fd_pr__cap_mim_m3_1_4HJTN9  XC2
timestamp 1712437813
transform 1 0 33062 0 1 -21822
box -7716 -4640 7716 4640
use sky130_fd_pr__cap_mim_m3_1_3DMTNZ  XC3
timestamp 1712540964
transform 1 0 9184 0 1 -4434
box -2492 -2320 2492 2320
use sky130_fd_pr__cap_mim_m3_1_4HHTN9  XC4
timestamp 1712073300
transform 0 -1 42836 1 0 -10682
box -1186 -4640 1186 4640
use sky130_fd_pr__nfet_g5v0d10v5_MHWJF7  XM1
timestamp 1712250795
transform 1 0 20755 0 1 -24504
box -989 -658 989 658
use sky130_fd_pr__pfet_g5v0d10v5_28EAA9  XM2
timestamp 1712250795
transform 0 1 20849 -1 0 -21271
box -2519 -697 2519 697
use sky130_fd_pr__nfet_01v8_AHZR5K  XM3
timestamp 1712071977
transform 1 0 39782 0 1 -9680
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_HZ6WG7  XM4
timestamp 1712071977
transform 1 0 46948 0 1 -11363
box -296 -285 296 285
use sky130_fd_pr__nfet_g5v0d10v5_ZPGQJT  XM5
timestamp 1712087189
transform -1 0 2862 0 1 -7654
box -594 -658 594 658
use sky130_fd_pr__pfet_g5v0d10v5_KLKQZ5  XM6
timestamp 1712087189
transform 1 0 4238 0 -1 -7655
box -624 -697 624 697
use sky130_fd_pr__pfet_01v8_3H68VM  XM7
timestamp 1712071977
transform 1 0 46810 0 1 -10257
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_XPHWY6  XM8
timestamp 1712087189
transform 1 0 16278 0 1 -1749
box -562 -1137 562 1137
use sky130_fd_pr__pfet_g5v0d10v5_KL3SY6  XM9
timestamp 1712071977
transform -1 0 16514 0 -1 -6935
box -308 -697 308 697
use sky130_fd_pr__nfet_01v8_Y5BWKS  XM11
timestamp 1712087189
transform 1 0 16360 0 1 -4521
box -562 -1119 562 1119
use sky130_fd_pr__res_xhigh_po_0p35_27M88N  XR2
timestamp 1712437813
transform 0 1 12474 -1 0 -27691
box -2359 -10982 2359 10982
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 dvdd
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 dvss
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 ibias
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 ena
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 standby
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 dout
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 xin
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 xout
port 9 nsew
<< end >>
