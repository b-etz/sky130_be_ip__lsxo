magic
tech sky130A
magscale 1 2
timestamp 1712875330
<< error_s >>
rect 3109 -1600 3430 -1248
rect 4910 -1600 5231 -1248
rect 12659 -3154 12980 -1974
rect 13188 -2839 20072 -2273
rect 12856 -3378 13170 -3364
rect 13406 -3398 13440 -3350
rect 13566 -3390 14044 -3364
rect 12890 -3412 14010 -3398
rect 12986 -3432 14010 -3412
rect 13406 -3668 13440 -3432
rect 13520 -3469 13558 -3462
rect 13508 -3484 13558 -3469
rect 13508 -3500 13566 -3484
rect 13834 -3500 13872 -3462
rect 13508 -3528 13872 -3500
rect 13516 -3532 13834 -3528
rect 13516 -3534 13850 -3532
rect 13542 -3540 13846 -3534
rect 13828 -3560 13930 -3550
rect 13570 -3566 13930 -3560
rect 13566 -3568 13900 -3566
rect 13582 -3572 13900 -3568
rect 13582 -3600 13908 -3572
rect 13850 -3616 13908 -3600
rect 13893 -3631 13908 -3616
rect 13862 -3660 13896 -3634
rect 13976 -3668 14010 -3432
rect 13406 -3702 14430 -3668
rect 13372 -3736 13850 -3710
rect 13976 -3750 14010 -3702
<< locali >>
rect 3872 -7142 4600 -7134
rect 2500 -7152 3228 -7142
rect 2500 -7216 2512 -7152
rect 3872 -7208 3888 -7142
rect 4588 -7208 4600 -7142
rect 2406 -7266 2526 -7254
rect 2406 -8042 2420 -7266
rect 2512 -8042 2526 -7266
rect 2406 -8054 2526 -8042
rect 2564 -7266 2684 -7254
rect 2564 -8042 2578 -7266
rect 2670 -8042 2684 -7266
rect 2564 -8054 2684 -8042
rect 2722 -7266 2842 -7254
rect 2722 -8042 2736 -7266
rect 2828 -8042 2842 -7266
rect 2722 -8054 2842 -8042
rect 2880 -7266 3000 -7254
rect 2880 -8042 2894 -7266
rect 2986 -8042 3000 -7266
rect 2880 -8054 3000 -8042
rect 3036 -7266 3156 -7254
rect 3036 -8042 3050 -7266
rect 3142 -8042 3156 -7266
rect 3036 -8054 3156 -8042
rect 3196 -7266 3316 -7254
rect 3196 -8042 3210 -7266
rect 3302 -8042 3316 -7266
rect 3196 -8054 3316 -8042
rect 3782 -7266 3902 -7254
rect 3782 -8044 3796 -7266
rect 3888 -8044 3902 -7266
rect 3782 -8054 3902 -8044
rect 3940 -7266 4060 -7254
rect 3940 -8044 3954 -7266
rect 4046 -8044 4060 -7266
rect 3940 -8054 4060 -8044
rect 4098 -7266 4218 -7254
rect 4098 -8044 4112 -7266
rect 4204 -8044 4218 -7266
rect 4098 -8054 4218 -8044
rect 4256 -7266 4376 -7254
rect 4256 -8044 4270 -7266
rect 4362 -8044 4376 -7266
rect 4256 -8054 4376 -8044
rect 4414 -7266 4534 -7254
rect 4414 -8044 4428 -7266
rect 4520 -8044 4534 -7266
rect 4414 -8054 4534 -8044
rect 4572 -7266 4692 -7254
rect 4572 -8044 4586 -7266
rect 4678 -8044 4692 -7266
rect 4572 -8054 4692 -8044
rect 2500 -8158 2512 -8092
rect 3212 -8158 3228 -8092
rect 2500 -8166 3228 -8158
rect 3872 -8168 3888 -8102
rect 4588 -8168 4600 -8102
rect 3872 -8176 4600 -8168
<< viali >>
rect 2512 -7216 3230 -7152
rect 3888 -7208 4588 -7142
rect 2420 -8042 2512 -7266
rect 2578 -8042 2670 -7266
rect 2736 -8042 2828 -7266
rect 2894 -8042 2986 -7266
rect 3050 -8042 3142 -7266
rect 3210 -8042 3302 -7266
rect 3796 -8044 3888 -7266
rect 3954 -8044 4046 -7266
rect 4112 -8044 4204 -7266
rect 4270 -8044 4362 -7266
rect 4428 -8044 4520 -7266
rect 4586 -8044 4678 -7266
rect 2512 -8158 3212 -8092
rect 3888 -8168 4588 -8102
<< metal1 >>
rect 1782 -1202 1982 -1002
rect 2242 -1202 2442 -1002
rect 2974 -1214 3174 -1014
rect 5136 -1192 5336 -992
rect 7066 -1128 7266 -928
rect 9806 -958 10006 -758
rect 11378 -950 11578 -750
rect 22408 -870 22608 -670
rect 3364 -7142 3370 -6962
rect 2500 -7152 3370 -7142
rect 2500 -7216 2512 -7152
rect 3230 -7216 3370 -7152
rect 2500 -7222 3370 -7216
rect 3478 -7222 3484 -6962
rect 3614 -7214 3620 -6954
rect 3728 -7134 3734 -6954
rect 3728 -7142 4600 -7134
rect 3728 -7208 3888 -7142
rect 4588 -7208 4600 -7142
rect 3728 -7214 4600 -7208
rect 2406 -8054 2412 -7254
rect 2520 -8054 2526 -7254
rect 2564 -8054 2570 -7254
rect 2678 -8054 2684 -7254
rect 2722 -8054 2728 -7254
rect 2836 -8054 2842 -7254
rect 2880 -8054 2886 -7254
rect 2994 -8054 3000 -7254
rect 3036 -8054 3042 -7254
rect 3150 -8054 3156 -7254
rect 3196 -8054 3202 -7254
rect 3310 -8054 3316 -7254
rect 3364 -8086 3370 -7906
rect 2500 -8092 3370 -8086
rect 2500 -8158 2512 -8092
rect 3212 -8158 3370 -8092
rect 2500 -8166 3370 -8158
rect 3478 -8086 3484 -7906
rect 3478 -8166 3486 -8086
rect 3614 -8176 3620 -7916
rect 3728 -8096 3734 -7916
rect 3782 -8054 3790 -7254
rect 3894 -8054 3902 -7254
rect 3940 -8054 3946 -7254
rect 4054 -8054 4060 -7254
rect 4098 -8054 4104 -7254
rect 4212 -8054 4218 -7254
rect 4256 -8054 4262 -7254
rect 4370 -8054 4376 -7254
rect 4414 -8054 4420 -7254
rect 4528 -8054 4534 -7254
rect 4572 -8054 4578 -7254
rect 4686 -8054 4692 -7254
rect 3728 -8102 4600 -8096
rect 3728 -8168 3888 -8102
rect 4588 -8168 4600 -8102
rect 3728 -8176 4600 -8168
rect 23936 -23898 24136 -23698
rect 1510 -24172 1710 -23972
<< via1 >>
rect 3370 -7222 3478 -6962
rect 3620 -7214 3728 -6954
rect 2412 -7266 2520 -7254
rect 2412 -8042 2420 -7266
rect 2420 -8042 2512 -7266
rect 2512 -8042 2520 -7266
rect 2412 -8054 2520 -8042
rect 2570 -7266 2678 -7254
rect 2570 -8042 2578 -7266
rect 2578 -8042 2670 -7266
rect 2670 -8042 2678 -7266
rect 2570 -8054 2678 -8042
rect 2728 -7266 2836 -7254
rect 2728 -8042 2736 -7266
rect 2736 -8042 2828 -7266
rect 2828 -8042 2836 -7266
rect 2728 -8054 2836 -8042
rect 2886 -7266 2994 -7254
rect 2886 -8042 2894 -7266
rect 2894 -8042 2986 -7266
rect 2986 -8042 2994 -7266
rect 2886 -8054 2994 -8042
rect 3042 -7266 3150 -7254
rect 3042 -8042 3050 -7266
rect 3050 -8042 3142 -7266
rect 3142 -8042 3150 -7266
rect 3042 -8054 3150 -8042
rect 3202 -7266 3310 -7254
rect 3202 -8042 3210 -7266
rect 3210 -8042 3302 -7266
rect 3302 -8042 3310 -7266
rect 3202 -8054 3310 -8042
rect 3370 -8166 3478 -7906
rect 3620 -8176 3728 -7916
rect 3790 -7266 3894 -7254
rect 3790 -8044 3796 -7266
rect 3796 -8044 3888 -7266
rect 3888 -8044 3894 -7266
rect 3790 -8054 3894 -8044
rect 3946 -7266 4054 -7254
rect 3946 -8044 3954 -7266
rect 3954 -8044 4046 -7266
rect 4046 -8044 4054 -7266
rect 3946 -8054 4054 -8044
rect 4104 -7266 4212 -7254
rect 4104 -8044 4112 -7266
rect 4112 -8044 4204 -7266
rect 4204 -8044 4212 -7266
rect 4104 -8054 4212 -8044
rect 4262 -7266 4370 -7254
rect 4262 -8044 4270 -7266
rect 4270 -8044 4362 -7266
rect 4362 -8044 4370 -7266
rect 4262 -8054 4370 -8044
rect 4420 -7266 4528 -7254
rect 4420 -8044 4428 -7266
rect 4428 -8044 4520 -7266
rect 4520 -8044 4528 -7266
rect 4420 -8054 4528 -8044
rect 4578 -7266 4686 -7254
rect 4578 -8044 4586 -7266
rect 4586 -8044 4678 -7266
rect 4678 -8044 4686 -7266
rect 4578 -8054 4686 -8044
<< metal2 >>
rect 2610 -6860 3484 -6740
rect 3364 -6962 3484 -6860
rect 2406 -7174 3158 -6974
rect 2406 -7254 2526 -7174
rect 2722 -7254 2842 -7174
rect 3036 -7254 3158 -7174
rect 3364 -7222 3370 -6962
rect 3478 -7222 3484 -6962
rect 2406 -8054 2412 -7254
rect 2520 -8054 2526 -7254
rect 2564 -8054 2570 -7254
rect 2678 -8054 2684 -7254
rect 2722 -8054 2728 -7254
rect 2836 -8054 2842 -7254
rect 2880 -8054 2886 -7254
rect 2994 -8054 3000 -7254
rect 3036 -8054 3042 -7254
rect 3150 -7554 3158 -7254
rect 3150 -8054 3156 -7554
rect 3196 -8054 3202 -7254
rect 3310 -8054 3316 -7254
rect 2564 -8134 2684 -8054
rect 2880 -8134 3000 -8054
rect 3196 -8134 3316 -8054
rect 2564 -8334 3316 -8134
rect 3364 -7906 3484 -7222
rect 3364 -8166 3370 -7906
rect 3478 -8166 3484 -7906
rect 3614 -6954 3734 -6750
rect 3614 -7214 3620 -6954
rect 3728 -7214 3734 -6954
rect 3614 -7916 3734 -7214
rect 3940 -7174 4692 -6974
rect 3940 -7254 4060 -7174
rect 4256 -7254 4376 -7174
rect 4572 -7254 4692 -7174
rect 3614 -8176 3620 -7916
rect 3728 -8176 3734 -7916
rect 3782 -8054 3790 -7254
rect 3894 -8054 3902 -7254
rect 3940 -8054 3946 -7254
rect 4054 -8054 4060 -7254
rect 4098 -8054 4104 -7254
rect 4212 -8054 4218 -7254
rect 4256 -8054 4262 -7254
rect 4370 -8054 4376 -7254
rect 4414 -8054 4420 -7254
rect 4528 -8054 4534 -7254
rect 4572 -8054 4578 -7254
rect 4686 -8054 4692 -7254
rect 3782 -8134 3902 -8054
rect 4098 -8134 4218 -8054
rect 4414 -8134 4534 -8054
rect 3782 -8334 4534 -8134
use sky130_fd_pr__cap_mim_m3_1_67RTNB  amp_XC1
timestamp 1712856537
transform 0 1 11932 -1 0 -7478
box -3798 -4640 3798 4640
use sky130_fd_pr__nfet_g5v0d10v5_554GUR  amp_XM1_2
timestamp 1712854380
transform 1 0 12515 0 1 -5116
box -2031 -458 2031 458
use sky130_fd_pr__pfet_01v8_T2YKL7  amp_XM3_5
timestamp 1712854380
transform 1 0 22729 0 1 -4817
box -1083 -619 1083 619
use sky130_fd_pr__nfet_01v8_8DG47J  amp_XM4_18
timestamp 1712854380
transform 1 0 22683 0 1 -6264
box -1083 -610 1083 610
use sky130_fd_pr__pfet_01v8_ED4X7U  amp_XM6_8
timestamp 1712854380
transform 0 1 9383 -1 0 -7765
box -1825 -269 1825 269
use sky130_fd_pr__nfet_01v8_YD343X  amp_XM7_9
timestamp 1712854380
transform 0 1 8460 -1 0 -7811
box -1825 -260 1825 260
use sky130_fd_pr__pfet_01v8_8D4V8N  amp_XM10_12
timestamp 1712854380
transform 1 0 19605 0 1 -6629
box -425 -383 425 383
use sky130_fd_pr__nfet_01v8_U59KY9  amp_XM11_13
timestamp 1712854380
transform 1 0 18395 0 1 -6669
box -425 -365 425 365
use sky130_fd_pr__pfet_g5v0d10v5_QS5HKK  amp_XM16_17
timestamp 1712854380
transform 1 0 12453 0 1 -6501
box -2061 -761 2061 761
use sky130_fd_pr__res_xhigh_po_0p35_F7SPRR  amp_XR1
timestamp 1712856537
transform 0 1 17212 -1 0 -9206
box -1612 -6832 1612 6832
use sky130_fd_pr__cap_mim_m3_1_VMUSDZ  bias_XC1
timestamp 1712851378
transform 0 -1 13238 1 0 -21322
box -2386 -11800 2386 11800
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  bias_XC2
timestamp 1712848480
transform 1 0 4112 0 1 -11804
box -2186 -2040 2186 2040
use sky130_fd_pr__cap_mim_m3_1_F5PPB9  bias_XC3
timestamp 1712849042
transform 0 1 9280 -1 0 -16342
box -1986 -7840 1986 7840
use sky130_fd_pr__nfet_g5v0d10v5_QNESWN  bias_XM1_2
timestamp 1712848480
transform 0 1 19622 -1 0 -15316
box -1802 -658 1802 658
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  bias_XM5
timestamp 1712848480
transform 1 0 6934 0 1 -12416
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_H6M2KM  bias_XM6_7_8
timestamp 1712851378
transform -1 0 10114 0 -1 -12418
box -2686 -300 2686 300
use sky130_fd_pr__res_xhigh_po_0p35_7UAGMY  bias_XR2
timestamp 1712849042
transform 0 1 10022 -1 0 -16453
box -2359 -8582 2359 8582
use sky130_fd_pr__res_xhigh_po_0p35_VTNT3C  bias_XR3
timestamp 1712851378
transform 0 1 10474 -1 0 -13400
box -450 -8082 450 8082
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712500979
transform 0 1 2848 -1 0 -1286
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x2
timestamp 1712500979
transform 0 -1 5492 -1 0 -1286
box -38 -48 314 592
use level_shift  x3
timestamp 1712539951
transform 0 1 4250 -1 0 -1190
box 652 -1950 5670 -128
use level_shift  x4
timestamp 1712539951
transform 0 -1 4086 -1 0 -1190
box 652 -1950 5670 -128
use ripl_dly_clk_buf  x7
timestamp 1712875330
transform 1 0 11856 0 1 -1322
box 216 -2416 8478 -290
use sky130_fd_pr__cap_mim_m3_1_KAF84V  XC1
timestamp 1712073300
transform 0 -1 10690 1 0 -12540
box -886 -3440 886 3440
use sky130_fd_pr__cap_mim_m3_1_4RGTN9  XC2
timestamp 1712848480
transform 1 0 21230 0 1 -9232
box -3798 -9280 3798 9280
use sky130_fd_pr__cap_mim_m3_1_3DMTNZ  XC3
timestamp 1712866372
transform 1 0 -2430 0 1 -3906
box -2492 -2320 2492 2320
use sky130_fd_pr__cap_mim_m3_1_4HHTN9  XC4
timestamp 1712866372
transform 0 -1 12224 1 0 -2198
box -1186 -4640 1186 4640
use sky130_fd_pr__nfet_g5v0d10v5_AB4DGB  XM1
timestamp 1712851712
transform 1 0 21667 0 1 -18058
box -1147 -658 1147 658
use sky130_fd_pr__pfet_g5v0d10v5_V6TMVM  XM2_bias_XM3_4
timestamp 1712848480
transform 0 1 21689 -1 0 -15091
box -2061 -1161 2061 1161
use sky130_fd_pr__nfet_01v8_AHZR5K  XM3
timestamp 1712867472
transform 1 0 13450 0 1 -3622
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_HZ6WG7  XM4
timestamp 1712071977
transform 1 0 21986 0 1 -1371
box -296 -285 296 285
use sky130_fd_pr__nfet_g5v0d10v5_ZPGQJT  XM5
timestamp 1712087189
transform -1 0 2862 0 1 -7654
box -594 -658 594 658
use sky130_fd_pr__pfet_g5v0d10v5_KLKQZ5  XM6
timestamp 1712087189
transform 1 0 4238 0 -1 -7655
box -624 -697 624 697
use sky130_fd_pr__pfet_01v8_3H68VM  XM7
timestamp 1712071977
transform 0 1 23155 -1 0 -1360
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_EDP4SU  XM8
timestamp 1712694485
transform 1 0 9915 0 1 -2827
box -957 -619 957 619
use sky130_fd_pr__pfet_g5v0d10v5_KL3SY6  XM9
timestamp 1712866372
transform -1 0 11588 0 -1 -2791
box -308 -697 308 697
use sky130_fd_pr__nfet_01v8_MLR4K3  XM11
timestamp 1712694485
transform 1 0 7837 0 1 -2836
box -957 -610 957 610
use sky130_fd_pr__res_xhigh_po_0p35_27M88N  XR2
timestamp 1712437813
transform 0 1 12478 -1 0 -21583
box -2359 -10982 2359 10982
<< labels >>
flabel metal1 23936 -23898 24136 -23698 0 FreeSans 256 0 0 0 xout
port 9 nsew
flabel metal1 22408 -870 22608 -670 0 FreeSans 256 0 0 0 dout
port 7 nsew
flabel metal1 5136 -1192 5336 -992 0 FreeSans 256 0 0 0 standby
port 6 nsew
flabel metal1 2974 -1214 3174 -1014 0 FreeSans 256 0 0 0 ena
port 5 nsew
flabel metal1 11378 -950 11578 -750 0 FreeSans 256 0 0 0 ibias
port 4 nsew
flabel metal1 7066 -1128 7266 -928 0 FreeSans 256 0 0 0 dvss
port 3 nsew
flabel metal1 9806 -958 10006 -758 0 FreeSans 256 0 0 0 dvdd
port 2 nsew
flabel metal1 2242 -1202 2442 -1002 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 1782 -1202 1982 -1002 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal1 1510 -24172 1710 -23972 0 FreeSans 256 0 0 0 xin
port 8 nsew
<< end >>
