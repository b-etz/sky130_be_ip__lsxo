magic
tech sky130A
magscale 1 2
timestamp 1712855660
<< pwell >>
rect -1114 -10582 1114 10582
<< psubdiff >>
rect -1078 10512 -982 10546
rect 982 10512 1078 10546
rect -1078 10450 -1044 10512
rect 1044 10450 1078 10512
rect -1078 -10512 -1044 -10450
rect 1044 -10512 1078 -10450
rect -1078 -10546 -982 -10512
rect 982 -10546 1078 -10512
<< psubdiffcont >>
rect -982 10512 982 10546
rect -1078 -10450 -1044 10450
rect 1044 -10450 1078 10450
rect -982 -10546 982 -10512
<< xpolycontact >>
rect -948 9984 -878 10416
rect -948 -10416 -878 -9984
rect -782 9984 -712 10416
rect -782 -10416 -712 -9984
rect -616 9984 -546 10416
rect -616 -10416 -546 -9984
rect -450 9984 -380 10416
rect -450 -10416 -380 -9984
rect -284 9984 -214 10416
rect -284 -10416 -214 -9984
rect -118 9984 -48 10416
rect -118 -10416 -48 -9984
rect 48 9984 118 10416
rect 48 -10416 118 -9984
rect 214 9984 284 10416
rect 214 -10416 284 -9984
rect 380 9984 450 10416
rect 380 -10416 450 -9984
rect 546 9984 616 10416
rect 546 -10416 616 -9984
rect 712 9984 782 10416
rect 712 -10416 782 -9984
rect 878 9984 948 10416
rect 878 -10416 948 -9984
<< xpolyres >>
rect -948 -9984 -878 9984
rect -782 -9984 -712 9984
rect -616 -9984 -546 9984
rect -450 -9984 -380 9984
rect -284 -9984 -214 9984
rect -118 -9984 -48 9984
rect 48 -9984 118 9984
rect 214 -9984 284 9984
rect 380 -9984 450 9984
rect 546 -9984 616 9984
rect 712 -9984 782 9984
rect 878 -9984 948 9984
<< locali >>
rect -1078 10512 -982 10546
rect 982 10512 1078 10546
rect -1078 10450 -1044 10512
rect 1044 10450 1078 10512
rect -1078 -10512 -1044 -10450
rect 1044 -10512 1078 -10450
rect -1078 -10546 -982 -10512
rect 982 -10546 1078 -10512
<< viali >>
rect -932 10001 -894 10398
rect -766 10001 -728 10398
rect -600 10001 -562 10398
rect -434 10001 -396 10398
rect -268 10001 -230 10398
rect -102 10001 -64 10398
rect 64 10001 102 10398
rect 230 10001 268 10398
rect 396 10001 434 10398
rect 562 10001 600 10398
rect 728 10001 766 10398
rect 894 10001 932 10398
rect -932 -10398 -894 -10001
rect -766 -10398 -728 -10001
rect -600 -10398 -562 -10001
rect -434 -10398 -396 -10001
rect -268 -10398 -230 -10001
rect -102 -10398 -64 -10001
rect 64 -10398 102 -10001
rect 230 -10398 268 -10001
rect 396 -10398 434 -10001
rect 562 -10398 600 -10001
rect 728 -10398 766 -10001
rect 894 -10398 932 -10001
<< metal1 >>
rect -938 10398 -888 10410
rect -938 10001 -932 10398
rect -894 10001 -888 10398
rect -938 9989 -888 10001
rect -772 10398 -722 10410
rect -772 10001 -766 10398
rect -728 10001 -722 10398
rect -772 9989 -722 10001
rect -606 10398 -556 10410
rect -606 10001 -600 10398
rect -562 10001 -556 10398
rect -606 9989 -556 10001
rect -440 10398 -390 10410
rect -440 10001 -434 10398
rect -396 10001 -390 10398
rect -440 9989 -390 10001
rect -274 10398 -224 10410
rect -274 10001 -268 10398
rect -230 10001 -224 10398
rect -274 9989 -224 10001
rect -108 10398 -58 10410
rect -108 10001 -102 10398
rect -64 10001 -58 10398
rect -108 9989 -58 10001
rect 58 10398 108 10410
rect 58 10001 64 10398
rect 102 10001 108 10398
rect 58 9989 108 10001
rect 224 10398 274 10410
rect 224 10001 230 10398
rect 268 10001 274 10398
rect 224 9989 274 10001
rect 390 10398 440 10410
rect 390 10001 396 10398
rect 434 10001 440 10398
rect 390 9989 440 10001
rect 556 10398 606 10410
rect 556 10001 562 10398
rect 600 10001 606 10398
rect 556 9989 606 10001
rect 722 10398 772 10410
rect 722 10001 728 10398
rect 766 10001 772 10398
rect 722 9989 772 10001
rect 888 10398 938 10410
rect 888 10001 894 10398
rect 932 10001 938 10398
rect 888 9989 938 10001
rect -938 -10001 -888 -9989
rect -938 -10398 -932 -10001
rect -894 -10398 -888 -10001
rect -938 -10410 -888 -10398
rect -772 -10001 -722 -9989
rect -772 -10398 -766 -10001
rect -728 -10398 -722 -10001
rect -772 -10410 -722 -10398
rect -606 -10001 -556 -9989
rect -606 -10398 -600 -10001
rect -562 -10398 -556 -10001
rect -606 -10410 -556 -10398
rect -440 -10001 -390 -9989
rect -440 -10398 -434 -10001
rect -396 -10398 -390 -10001
rect -440 -10410 -390 -10398
rect -274 -10001 -224 -9989
rect -274 -10398 -268 -10001
rect -230 -10398 -224 -10001
rect -274 -10410 -224 -10398
rect -108 -10001 -58 -9989
rect -108 -10398 -102 -10001
rect -64 -10398 -58 -10001
rect -108 -10410 -58 -10398
rect 58 -10001 108 -9989
rect 58 -10398 64 -10001
rect 102 -10398 108 -10001
rect 58 -10410 108 -10398
rect 224 -10001 274 -9989
rect 224 -10398 230 -10001
rect 268 -10398 274 -10001
rect 224 -10410 274 -10398
rect 390 -10001 440 -9989
rect 390 -10398 396 -10001
rect 434 -10398 440 -10001
rect 390 -10410 440 -10398
rect 556 -10001 606 -9989
rect 556 -10398 562 -10001
rect 600 -10398 606 -10001
rect 556 -10410 606 -10398
rect 722 -10001 772 -9989
rect 722 -10398 728 -10001
rect 766 -10398 772 -10001
rect 722 -10410 772 -10398
rect 888 -10001 938 -9989
rect 888 -10398 894 -10001
rect 932 -10398 938 -10001
rect 888 -10410 938 -10398
<< properties >>
string FIXED_BBOX -1061 -10529 1061 10529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 100 m 1 nx 12 wmin 0.350 lmin 0.50 rho 2000 val 572.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
