magic
tech sky130A
magscale 1 2
timestamp 1713105616
<< metal3 >>
rect -886 1840 586 3320
rect -886 120 586 1600
rect -886 -1600 586 -120
rect -886 -3320 586 -1840
<< mimcap >>
rect -846 3240 554 3280
rect -846 1920 -806 3240
rect 514 1920 554 3240
rect -846 1880 554 1920
rect -846 1520 554 1560
rect -846 200 -806 1520
rect 514 200 554 1520
rect -846 160 554 200
rect -846 -200 554 -160
rect -846 -1520 -806 -200
rect 514 -1520 554 -200
rect -846 -1560 554 -1520
rect -846 -1920 554 -1880
rect -846 -3240 -806 -1920
rect 514 -3240 554 -1920
rect -846 -3280 554 -3240
<< mimcapcontact >>
rect -806 1920 514 3240
rect -806 200 514 1520
rect -806 -1520 514 -200
rect -806 -3240 514 -1920
<< metal4 >>
rect -198 3241 -94 3440
rect -807 3240 515 3241
rect -807 1920 -806 3240
rect 514 1920 515 3240
rect -807 1919 515 1920
rect -198 1521 -94 1919
rect -807 1520 515 1521
rect -807 200 -806 1520
rect 514 200 515 1520
rect -807 199 515 200
rect -198 -199 -94 199
rect -807 -200 515 -199
rect -807 -1520 -806 -200
rect 514 -1520 515 -200
rect -807 -1521 515 -1520
rect -198 -1919 -94 -1521
rect -807 -1920 515 -1919
rect -807 -3240 -806 -1920
rect 514 -3240 515 -1920
rect -807 -3241 515 -3240
rect -198 -3440 -94 -3241
<< properties >>
string FIXED_BBOX -886 1840 594 3320
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 7.0 l 7.0 val 103.32 carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
