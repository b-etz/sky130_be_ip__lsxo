magic
tech sky130A
timestamp 1713017924
<< psubdiff >>
rect 236 -847 266 -835
rect 236 -889 266 -877
<< psubdiffcont >>
rect 236 -877 266 -847
<< locali >>
rect 108 -260 399 -253
rect 108 -346 115 -260
rect 201 -278 399 -260
rect 201 -346 208 -278
rect 108 -353 208 -346
rect 379 -388 399 -278
rect 371 -706 443 -695
rect 371 -730 381 -706
rect 431 -730 443 -706
rect 236 -847 266 -839
rect 236 -885 266 -877
rect 297 -914 330 -830
rect 297 -921 347 -914
rect 383 -978 433 -864
rect 484 -914 517 -830
rect 484 -921 534 -914
rect 607 -978 657 -476
rect 245 -1028 657 -978
rect 245 -1034 345 -1028
rect 245 -1200 252 -1034
rect 338 -1200 345 -1034
rect 245 -1208 345 -1200
<< viali >>
rect 115 -346 201 -260
rect 379 -450 398 -406
rect 346 -507 392 -490
rect 345 -565 391 -548
rect 379 -634 398 -595
rect 381 -756 431 -706
rect 297 -961 347 -921
rect 484 -961 534 -921
rect 252 -1200 338 -1034
<< metal1 >>
rect 247 -128 735 -78
rect 108 -258 208 -253
rect 108 -348 113 -258
rect 203 -348 208 -258
rect 108 -353 208 -348
rect 247 -355 295 -128
rect 494 -152 594 -145
rect 494 -239 501 -152
rect 587 -239 594 -152
rect 494 -245 594 -239
rect 519 -345 567 -245
rect 685 -369 735 -128
rect 4345 -369 4495 -321
rect 371 -406 495 -399
rect 371 -452 378 -406
rect 488 -452 495 -406
rect 371 -459 495 -452
rect 339 -482 399 -479
rect 339 -508 343 -482
rect 396 -508 399 -482
rect 339 -511 399 -508
rect 339 -545 399 -542
rect 339 -571 343 -545
rect 396 -571 399 -545
rect 339 -574 399 -571
rect 4345 -587 4415 -582
rect 370 -595 494 -592
rect 370 -599 379 -595
rect 398 -599 494 -595
rect 370 -645 377 -599
rect 487 -645 494 -599
rect 543 -641 717 -593
rect 370 -652 494 -645
rect 4345 -647 4350 -587
rect 4410 -647 4415 -587
rect 4345 -652 4415 -647
rect 370 -706 443 -695
rect 370 -756 381 -706
rect 431 -756 443 -706
rect 370 -778 443 -756
rect 370 -844 410 -778
rect 370 -878 373 -844
rect 407 -878 410 -844
rect 4445 -865 4495 -369
rect 370 -881 410 -878
rect 288 -921 543 -913
rect 288 -961 297 -921
rect 347 -961 484 -921
rect 534 -961 543 -921
rect 288 -969 543 -961
rect 245 -1034 345 -1028
rect 245 -1200 252 -1034
rect 338 -1200 345 -1034
rect 245 -1208 345 -1200
rect 443 -1053 543 -969
rect 857 -994 1252 -988
rect 857 -1033 863 -994
rect 1246 -1033 1252 -994
rect 857 -1037 1252 -1033
rect 1303 -1053 1353 -896
rect 4345 -913 4495 -865
rect 443 -1103 852 -1053
rect 1258 -1103 1353 -1053
rect 443 -1208 543 -1103
<< via1 >>
rect 113 -260 203 -258
rect 113 -346 115 -260
rect 115 -346 201 -260
rect 201 -346 203 -260
rect 113 -348 203 -346
rect 501 -239 587 -152
rect 378 -450 379 -406
rect 379 -450 398 -406
rect 398 -450 488 -406
rect 378 -452 488 -450
rect 343 -490 396 -482
rect 343 -507 346 -490
rect 346 -507 392 -490
rect 392 -507 396 -490
rect 343 -508 396 -507
rect 343 -548 396 -545
rect 343 -565 345 -548
rect 345 -565 391 -548
rect 391 -565 396 -548
rect 343 -571 396 -565
rect 377 -634 379 -599
rect 379 -634 398 -599
rect 398 -634 487 -599
rect 377 -645 487 -634
rect 4350 -647 4410 -587
rect 373 -878 407 -844
rect 863 -1033 1246 -994
<< metal2 >>
rect 494 -152 594 -145
rect 494 -239 501 -152
rect 587 -239 594 -152
rect 494 -245 594 -239
rect 108 -258 208 -253
rect 108 -348 113 -258
rect 203 -348 208 -258
rect 108 -353 208 -348
rect 455 -321 899 -271
rect 455 -399 495 -321
rect 371 -406 495 -399
rect 108 -475 208 -415
rect 371 -452 378 -406
rect 488 -452 495 -406
rect 371 -459 495 -452
rect 640 -475 680 -434
rect 849 -456 899 -321
rect 108 -482 680 -475
rect 108 -508 343 -482
rect 396 -508 680 -482
rect 108 -515 680 -508
rect 108 -545 680 -538
rect 108 -571 343 -545
rect 396 -571 680 -545
rect 108 -578 680 -571
rect 108 -638 208 -578
rect 370 -599 494 -592
rect 370 -645 377 -599
rect 487 -645 494 -599
rect 370 -652 494 -645
rect 370 -844 410 -841
rect 370 -878 373 -844
rect 407 -878 410 -844
rect 370 -989 410 -878
rect 454 -913 494 -652
rect 640 -804 680 -578
rect 4345 -587 4415 -582
rect 4345 -647 4350 -587
rect 4410 -647 4415 -587
rect 4345 -652 4415 -647
rect 849 -913 899 -778
rect 454 -963 899 -913
rect 370 -994 1252 -989
rect 370 -1019 863 -994
rect 857 -1033 863 -1019
rect 1246 -1033 1252 -994
rect 857 -1037 1252 -1033
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1713017924
transform 0 1 271 -1 0 -299
box -19 -24 65 296
use ripple_dly_4  x1
timestamp 1713017924
transform 1 0 689 0 -1 -935
box -49 -614 3675 -294
use ripple_dly_4  x2
timestamp 1713017924
transform 1 0 689 0 1 -299
box -49 -614 3675 -294
use sky130_fd_sc_hd__a221o_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1713017924
transform 0 1 271 -1 0 -345
box -19 -24 387 296
use sky130_fd_sc_hd__einvn_0  x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1713017924
transform 0 1 271 -1 0 -713
box -19 -24 203 296
use sky130_fd_pr__nfet_01v8_AHZR5K  XM3
timestamp 1713017924
transform 1 0 1055 0 1 -1078
box -298 -130 298 130
<< labels >>
flabel metal1 443 -1208 543 -961 0 FreeSans 400 0 0 0 clkout
port 4 nsew
flabel metal1 245 -1208 345 -1028 0 FreeSans 400 0 0 0 clkin
port 3 nsew
flabel metal2 108 -515 208 -415 0 FreeSans 400 0 0 0 ena
port 5 nsew
flabel metal2 108 -638 208 -538 0 FreeSans 400 0 0 0 stby_b
port 8 nsew
flabel metal2 494 -245 594 -145 0 FreeSans 400 0 0 0 dvdd
port 1 nsew
flabel metal2 108 -353 208 -253 0 FreeSans 400 0 0 0 stby
port 6 nsew
flabel metal1 4445 -913 4495 -321 0 FreeSans 400 0 0 0 dvss
port 2 nsew
<< end >>
