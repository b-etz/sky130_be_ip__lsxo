magic
tech sky130A
magscale 1 2
timestamp 1712250795
<< pwell >>
rect -2276 -10582 2276 10582
<< psubdiff >>
rect -2240 10512 -2144 10546
rect 2144 10512 2240 10546
rect -2240 10450 -2206 10512
rect 2206 10450 2240 10512
rect -2240 -10512 -2206 -10450
rect 2206 -10512 2240 -10450
rect -2240 -10546 -2144 -10512
rect 2144 -10546 2240 -10512
<< psubdiffcont >>
rect -2144 10512 2144 10546
rect -2240 -10450 -2206 10450
rect 2206 -10450 2240 10450
rect -2144 -10546 2144 -10512
<< xpolycontact >>
rect -2110 9984 -2040 10416
rect -2110 -10416 -2040 -9984
rect -1944 9984 -1874 10416
rect -1944 -10416 -1874 -9984
rect -1778 9984 -1708 10416
rect -1778 -10416 -1708 -9984
rect -1612 9984 -1542 10416
rect -1612 -10416 -1542 -9984
rect -1446 9984 -1376 10416
rect -1446 -10416 -1376 -9984
rect -1280 9984 -1210 10416
rect -1280 -10416 -1210 -9984
rect -1114 9984 -1044 10416
rect -1114 -10416 -1044 -9984
rect -948 9984 -878 10416
rect -948 -10416 -878 -9984
rect -782 9984 -712 10416
rect -782 -10416 -712 -9984
rect -616 9984 -546 10416
rect -616 -10416 -546 -9984
rect -450 9984 -380 10416
rect -450 -10416 -380 -9984
rect -284 9984 -214 10416
rect -284 -10416 -214 -9984
rect -118 9984 -48 10416
rect -118 -10416 -48 -9984
rect 48 9984 118 10416
rect 48 -10416 118 -9984
rect 214 9984 284 10416
rect 214 -10416 284 -9984
rect 380 9984 450 10416
rect 380 -10416 450 -9984
rect 546 9984 616 10416
rect 546 -10416 616 -9984
rect 712 9984 782 10416
rect 712 -10416 782 -9984
rect 878 9984 948 10416
rect 878 -10416 948 -9984
rect 1044 9984 1114 10416
rect 1044 -10416 1114 -9984
rect 1210 9984 1280 10416
rect 1210 -10416 1280 -9984
rect 1376 9984 1446 10416
rect 1376 -10416 1446 -9984
rect 1542 9984 1612 10416
rect 1542 -10416 1612 -9984
rect 1708 9984 1778 10416
rect 1708 -10416 1778 -9984
rect 1874 9984 1944 10416
rect 1874 -10416 1944 -9984
rect 2040 9984 2110 10416
rect 2040 -10416 2110 -9984
<< xpolyres >>
rect -2110 -9984 -2040 9984
rect -1944 -9984 -1874 9984
rect -1778 -9984 -1708 9984
rect -1612 -9984 -1542 9984
rect -1446 -9984 -1376 9984
rect -1280 -9984 -1210 9984
rect -1114 -9984 -1044 9984
rect -948 -9984 -878 9984
rect -782 -9984 -712 9984
rect -616 -9984 -546 9984
rect -450 -9984 -380 9984
rect -284 -9984 -214 9984
rect -118 -9984 -48 9984
rect 48 -9984 118 9984
rect 214 -9984 284 9984
rect 380 -9984 450 9984
rect 546 -9984 616 9984
rect 712 -9984 782 9984
rect 878 -9984 948 9984
rect 1044 -9984 1114 9984
rect 1210 -9984 1280 9984
rect 1376 -9984 1446 9984
rect 1542 -9984 1612 9984
rect 1708 -9984 1778 9984
rect 1874 -9984 1944 9984
rect 2040 -9984 2110 9984
<< locali >>
rect -2240 10512 -2144 10546
rect 2144 10512 2240 10546
rect -2240 10450 -2206 10512
rect 2206 10450 2240 10512
rect -2240 -10512 -2206 -10450
rect 2206 -10512 2240 -10450
rect -2240 -10546 -2144 -10512
rect 2144 -10546 2240 -10512
<< viali >>
rect -2094 10001 -2056 10398
rect -1928 10001 -1890 10398
rect -1762 10001 -1724 10398
rect -1596 10001 -1558 10398
rect -1430 10001 -1392 10398
rect -1264 10001 -1226 10398
rect -1098 10001 -1060 10398
rect -932 10001 -894 10398
rect -766 10001 -728 10398
rect -600 10001 -562 10398
rect -434 10001 -396 10398
rect -268 10001 -230 10398
rect -102 10001 -64 10398
rect 64 10001 102 10398
rect 230 10001 268 10398
rect 396 10001 434 10398
rect 562 10001 600 10398
rect 728 10001 766 10398
rect 894 10001 932 10398
rect 1060 10001 1098 10398
rect 1226 10001 1264 10398
rect 1392 10001 1430 10398
rect 1558 10001 1596 10398
rect 1724 10001 1762 10398
rect 1890 10001 1928 10398
rect 2056 10001 2094 10398
rect -2094 -10398 -2056 -10001
rect -1928 -10398 -1890 -10001
rect -1762 -10398 -1724 -10001
rect -1596 -10398 -1558 -10001
rect -1430 -10398 -1392 -10001
rect -1264 -10398 -1226 -10001
rect -1098 -10398 -1060 -10001
rect -932 -10398 -894 -10001
rect -766 -10398 -728 -10001
rect -600 -10398 -562 -10001
rect -434 -10398 -396 -10001
rect -268 -10398 -230 -10001
rect -102 -10398 -64 -10001
rect 64 -10398 102 -10001
rect 230 -10398 268 -10001
rect 396 -10398 434 -10001
rect 562 -10398 600 -10001
rect 728 -10398 766 -10001
rect 894 -10398 932 -10001
rect 1060 -10398 1098 -10001
rect 1226 -10398 1264 -10001
rect 1392 -10398 1430 -10001
rect 1558 -10398 1596 -10001
rect 1724 -10398 1762 -10001
rect 1890 -10398 1928 -10001
rect 2056 -10398 2094 -10001
<< metal1 >>
rect -2100 10398 -2050 10410
rect -2100 10001 -2094 10398
rect -2056 10001 -2050 10398
rect -2100 9989 -2050 10001
rect -1934 10398 -1884 10410
rect -1934 10001 -1928 10398
rect -1890 10001 -1884 10398
rect -1934 9989 -1884 10001
rect -1768 10398 -1718 10410
rect -1768 10001 -1762 10398
rect -1724 10001 -1718 10398
rect -1768 9989 -1718 10001
rect -1602 10398 -1552 10410
rect -1602 10001 -1596 10398
rect -1558 10001 -1552 10398
rect -1602 9989 -1552 10001
rect -1436 10398 -1386 10410
rect -1436 10001 -1430 10398
rect -1392 10001 -1386 10398
rect -1436 9989 -1386 10001
rect -1270 10398 -1220 10410
rect -1270 10001 -1264 10398
rect -1226 10001 -1220 10398
rect -1270 9989 -1220 10001
rect -1104 10398 -1054 10410
rect -1104 10001 -1098 10398
rect -1060 10001 -1054 10398
rect -1104 9989 -1054 10001
rect -938 10398 -888 10410
rect -938 10001 -932 10398
rect -894 10001 -888 10398
rect -938 9989 -888 10001
rect -772 10398 -722 10410
rect -772 10001 -766 10398
rect -728 10001 -722 10398
rect -772 9989 -722 10001
rect -606 10398 -556 10410
rect -606 10001 -600 10398
rect -562 10001 -556 10398
rect -606 9989 -556 10001
rect -440 10398 -390 10410
rect -440 10001 -434 10398
rect -396 10001 -390 10398
rect -440 9989 -390 10001
rect -274 10398 -224 10410
rect -274 10001 -268 10398
rect -230 10001 -224 10398
rect -274 9989 -224 10001
rect -108 10398 -58 10410
rect -108 10001 -102 10398
rect -64 10001 -58 10398
rect -108 9989 -58 10001
rect 58 10398 108 10410
rect 58 10001 64 10398
rect 102 10001 108 10398
rect 58 9989 108 10001
rect 224 10398 274 10410
rect 224 10001 230 10398
rect 268 10001 274 10398
rect 224 9989 274 10001
rect 390 10398 440 10410
rect 390 10001 396 10398
rect 434 10001 440 10398
rect 390 9989 440 10001
rect 556 10398 606 10410
rect 556 10001 562 10398
rect 600 10001 606 10398
rect 556 9989 606 10001
rect 722 10398 772 10410
rect 722 10001 728 10398
rect 766 10001 772 10398
rect 722 9989 772 10001
rect 888 10398 938 10410
rect 888 10001 894 10398
rect 932 10001 938 10398
rect 888 9989 938 10001
rect 1054 10398 1104 10410
rect 1054 10001 1060 10398
rect 1098 10001 1104 10398
rect 1054 9989 1104 10001
rect 1220 10398 1270 10410
rect 1220 10001 1226 10398
rect 1264 10001 1270 10398
rect 1220 9989 1270 10001
rect 1386 10398 1436 10410
rect 1386 10001 1392 10398
rect 1430 10001 1436 10398
rect 1386 9989 1436 10001
rect 1552 10398 1602 10410
rect 1552 10001 1558 10398
rect 1596 10001 1602 10398
rect 1552 9989 1602 10001
rect 1718 10398 1768 10410
rect 1718 10001 1724 10398
rect 1762 10001 1768 10398
rect 1718 9989 1768 10001
rect 1884 10398 1934 10410
rect 1884 10001 1890 10398
rect 1928 10001 1934 10398
rect 1884 9989 1934 10001
rect 2050 10398 2100 10410
rect 2050 10001 2056 10398
rect 2094 10001 2100 10398
rect 2050 9989 2100 10001
rect -2100 -10001 -2050 -9989
rect -2100 -10398 -2094 -10001
rect -2056 -10398 -2050 -10001
rect -2100 -10410 -2050 -10398
rect -1934 -10001 -1884 -9989
rect -1934 -10398 -1928 -10001
rect -1890 -10398 -1884 -10001
rect -1934 -10410 -1884 -10398
rect -1768 -10001 -1718 -9989
rect -1768 -10398 -1762 -10001
rect -1724 -10398 -1718 -10001
rect -1768 -10410 -1718 -10398
rect -1602 -10001 -1552 -9989
rect -1602 -10398 -1596 -10001
rect -1558 -10398 -1552 -10001
rect -1602 -10410 -1552 -10398
rect -1436 -10001 -1386 -9989
rect -1436 -10398 -1430 -10001
rect -1392 -10398 -1386 -10001
rect -1436 -10410 -1386 -10398
rect -1270 -10001 -1220 -9989
rect -1270 -10398 -1264 -10001
rect -1226 -10398 -1220 -10001
rect -1270 -10410 -1220 -10398
rect -1104 -10001 -1054 -9989
rect -1104 -10398 -1098 -10001
rect -1060 -10398 -1054 -10001
rect -1104 -10410 -1054 -10398
rect -938 -10001 -888 -9989
rect -938 -10398 -932 -10001
rect -894 -10398 -888 -10001
rect -938 -10410 -888 -10398
rect -772 -10001 -722 -9989
rect -772 -10398 -766 -10001
rect -728 -10398 -722 -10001
rect -772 -10410 -722 -10398
rect -606 -10001 -556 -9989
rect -606 -10398 -600 -10001
rect -562 -10398 -556 -10001
rect -606 -10410 -556 -10398
rect -440 -10001 -390 -9989
rect -440 -10398 -434 -10001
rect -396 -10398 -390 -10001
rect -440 -10410 -390 -10398
rect -274 -10001 -224 -9989
rect -274 -10398 -268 -10001
rect -230 -10398 -224 -10001
rect -274 -10410 -224 -10398
rect -108 -10001 -58 -9989
rect -108 -10398 -102 -10001
rect -64 -10398 -58 -10001
rect -108 -10410 -58 -10398
rect 58 -10001 108 -9989
rect 58 -10398 64 -10001
rect 102 -10398 108 -10001
rect 58 -10410 108 -10398
rect 224 -10001 274 -9989
rect 224 -10398 230 -10001
rect 268 -10398 274 -10001
rect 224 -10410 274 -10398
rect 390 -10001 440 -9989
rect 390 -10398 396 -10001
rect 434 -10398 440 -10001
rect 390 -10410 440 -10398
rect 556 -10001 606 -9989
rect 556 -10398 562 -10001
rect 600 -10398 606 -10001
rect 556 -10410 606 -10398
rect 722 -10001 772 -9989
rect 722 -10398 728 -10001
rect 766 -10398 772 -10001
rect 722 -10410 772 -10398
rect 888 -10001 938 -9989
rect 888 -10398 894 -10001
rect 932 -10398 938 -10001
rect 888 -10410 938 -10398
rect 1054 -10001 1104 -9989
rect 1054 -10398 1060 -10001
rect 1098 -10398 1104 -10001
rect 1054 -10410 1104 -10398
rect 1220 -10001 1270 -9989
rect 1220 -10398 1226 -10001
rect 1264 -10398 1270 -10001
rect 1220 -10410 1270 -10398
rect 1386 -10001 1436 -9989
rect 1386 -10398 1392 -10001
rect 1430 -10398 1436 -10001
rect 1386 -10410 1436 -10398
rect 1552 -10001 1602 -9989
rect 1552 -10398 1558 -10001
rect 1596 -10398 1602 -10001
rect 1552 -10410 1602 -10398
rect 1718 -10001 1768 -9989
rect 1718 -10398 1724 -10001
rect 1762 -10398 1768 -10001
rect 1718 -10410 1768 -10398
rect 1884 -10001 1934 -9989
rect 1884 -10398 1890 -10001
rect 1928 -10398 1934 -10001
rect 1884 -10410 1934 -10398
rect 2050 -10001 2100 -9989
rect 2050 -10398 2056 -10001
rect 2094 -10398 2100 -10001
rect 2050 -10410 2100 -10398
<< properties >>
string FIXED_BBOX -2223 -10529 2223 10529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 100 m 1 nx 26 wmin 0.350 lmin 0.50 rho 2000 val 572.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
