magic
tech sky130A
magscale 1 2
timestamp 1713225924
<< pwell >>
rect -2451 -458 2451 458
<< mvnmos >>
rect -2223 -200 -1823 200
rect -1645 -200 -1245 200
rect -1067 -200 -667 200
rect -489 -200 -89 200
rect 89 -200 489 200
rect 667 -200 1067 200
rect 1245 -200 1645 200
rect 1823 -200 2223 200
<< mvndiff >>
rect -2281 188 -2223 200
rect -2281 -188 -2269 188
rect -2235 -188 -2223 188
rect -2281 -200 -2223 -188
rect -1823 188 -1765 200
rect -1823 -188 -1811 188
rect -1777 -188 -1765 188
rect -1823 -200 -1765 -188
rect -1703 188 -1645 200
rect -1703 -188 -1691 188
rect -1657 -188 -1645 188
rect -1703 -200 -1645 -188
rect -1245 188 -1187 200
rect -1245 -188 -1233 188
rect -1199 -188 -1187 188
rect -1245 -200 -1187 -188
rect -1125 188 -1067 200
rect -1125 -188 -1113 188
rect -1079 -188 -1067 188
rect -1125 -200 -1067 -188
rect -667 188 -609 200
rect -667 -188 -655 188
rect -621 -188 -609 188
rect -667 -200 -609 -188
rect -547 188 -489 200
rect -547 -188 -535 188
rect -501 -188 -489 188
rect -547 -200 -489 -188
rect -89 188 -31 200
rect -89 -188 -77 188
rect -43 -188 -31 188
rect -89 -200 -31 -188
rect 31 188 89 200
rect 31 -188 43 188
rect 77 -188 89 188
rect 31 -200 89 -188
rect 489 188 547 200
rect 489 -188 501 188
rect 535 -188 547 188
rect 489 -200 547 -188
rect 609 188 667 200
rect 609 -188 621 188
rect 655 -188 667 188
rect 609 -200 667 -188
rect 1067 188 1125 200
rect 1067 -188 1079 188
rect 1113 -188 1125 188
rect 1067 -200 1125 -188
rect 1187 188 1245 200
rect 1187 -188 1199 188
rect 1233 -188 1245 188
rect 1187 -200 1245 -188
rect 1645 188 1703 200
rect 1645 -188 1657 188
rect 1691 -188 1703 188
rect 1645 -200 1703 -188
rect 1765 188 1823 200
rect 1765 -188 1777 188
rect 1811 -188 1823 188
rect 1765 -200 1823 -188
rect 2223 188 2281 200
rect 2223 -188 2235 188
rect 2269 -188 2281 188
rect 2223 -200 2281 -188
<< mvndiffc >>
rect -2269 -188 -2235 188
rect -1811 -188 -1777 188
rect -1691 -188 -1657 188
rect -1233 -188 -1199 188
rect -1113 -188 -1079 188
rect -655 -188 -621 188
rect -535 -188 -501 188
rect -77 -188 -43 188
rect 43 -188 77 188
rect 501 -188 535 188
rect 621 -188 655 188
rect 1079 -188 1113 188
rect 1199 -188 1233 188
rect 1657 -188 1691 188
rect 1777 -188 1811 188
rect 2235 -188 2269 188
<< mvpsubdiff >>
rect -2415 410 2415 422
rect -2415 376 -2307 410
rect 2307 376 2415 410
rect -2415 364 2415 376
rect -2415 314 -2357 364
rect -2415 -314 -2403 314
rect -2369 -314 -2357 314
rect 2357 314 2415 364
rect -2415 -364 -2357 -314
rect 2357 -314 2369 314
rect 2403 -314 2415 314
rect 2357 -364 2415 -314
rect -2415 -376 2415 -364
rect -2415 -410 -2307 -376
rect 2307 -410 2415 -376
rect -2415 -422 2415 -410
<< mvpsubdiffcont >>
rect -2307 376 2307 410
rect -2403 -314 -2369 314
rect 2369 -314 2403 314
rect -2307 -410 2307 -376
<< poly >>
rect -2223 272 -1823 288
rect -2223 238 -2207 272
rect -1839 238 -1823 272
rect -2223 200 -1823 238
rect -1645 272 -1245 288
rect -1645 238 -1629 272
rect -1261 238 -1245 272
rect -1645 200 -1245 238
rect -1067 272 -667 288
rect -1067 238 -1051 272
rect -683 238 -667 272
rect -1067 200 -667 238
rect -489 272 -89 288
rect -489 238 -473 272
rect -105 238 -89 272
rect -489 200 -89 238
rect 89 272 489 288
rect 89 238 105 272
rect 473 238 489 272
rect 89 200 489 238
rect 667 272 1067 288
rect 667 238 683 272
rect 1051 238 1067 272
rect 667 200 1067 238
rect 1245 272 1645 288
rect 1245 238 1261 272
rect 1629 238 1645 272
rect 1245 200 1645 238
rect 1823 272 2223 288
rect 1823 238 1839 272
rect 2207 238 2223 272
rect 1823 200 2223 238
rect -2223 -238 -1823 -200
rect -2223 -272 -2207 -238
rect -1839 -272 -1823 -238
rect -2223 -288 -1823 -272
rect -1645 -238 -1245 -200
rect -1645 -272 -1629 -238
rect -1261 -272 -1245 -238
rect -1645 -288 -1245 -272
rect -1067 -238 -667 -200
rect -1067 -272 -1051 -238
rect -683 -272 -667 -238
rect -1067 -288 -667 -272
rect -489 -238 -89 -200
rect -489 -272 -473 -238
rect -105 -272 -89 -238
rect -489 -288 -89 -272
rect 89 -238 489 -200
rect 89 -272 105 -238
rect 473 -272 489 -238
rect 89 -288 489 -272
rect 667 -238 1067 -200
rect 667 -272 683 -238
rect 1051 -272 1067 -238
rect 667 -288 1067 -272
rect 1245 -238 1645 -200
rect 1245 -272 1261 -238
rect 1629 -272 1645 -238
rect 1245 -288 1645 -272
rect 1823 -238 2223 -200
rect 1823 -272 1839 -238
rect 2207 -272 2223 -238
rect 1823 -288 2223 -272
<< polycont >>
rect -2207 238 -1839 272
rect -1629 238 -1261 272
rect -1051 238 -683 272
rect -473 238 -105 272
rect 105 238 473 272
rect 683 238 1051 272
rect 1261 238 1629 272
rect 1839 238 2207 272
rect -2207 -272 -1839 -238
rect -1629 -272 -1261 -238
rect -1051 -272 -683 -238
rect -473 -272 -105 -238
rect 105 -272 473 -238
rect 683 -272 1051 -238
rect 1261 -272 1629 -238
rect 1839 -272 2207 -238
<< locali >>
rect -2403 376 -2307 410
rect 2307 376 2403 410
rect -2403 314 -2369 376
rect 2369 314 2403 376
rect -2223 238 -2207 272
rect -1839 238 -1823 272
rect -1645 238 -1629 272
rect -1261 238 -1245 272
rect -1067 238 -1051 272
rect -683 238 -667 272
rect -489 238 -473 272
rect -105 238 -89 272
rect 89 238 105 272
rect 473 238 489 272
rect 667 238 683 272
rect 1051 238 1067 272
rect 1245 238 1261 272
rect 1629 238 1645 272
rect 1823 238 1839 272
rect 2207 238 2223 272
rect -2269 188 -2235 204
rect -2269 -204 -2235 -188
rect -1811 188 -1777 204
rect -1811 -204 -1777 -188
rect -1691 188 -1657 204
rect -1691 -204 -1657 -188
rect -1233 188 -1199 204
rect -1233 -204 -1199 -188
rect -1113 188 -1079 204
rect -1113 -204 -1079 -188
rect -655 188 -621 204
rect -655 -204 -621 -188
rect -535 188 -501 204
rect -535 -204 -501 -188
rect -77 188 -43 204
rect -77 -204 -43 -188
rect 43 188 77 204
rect 43 -204 77 -188
rect 501 188 535 204
rect 501 -204 535 -188
rect 621 188 655 204
rect 621 -204 655 -188
rect 1079 188 1113 204
rect 1079 -204 1113 -188
rect 1199 188 1233 204
rect 1199 -204 1233 -188
rect 1657 188 1691 204
rect 1657 -204 1691 -188
rect 1777 188 1811 204
rect 1777 -204 1811 -188
rect 2235 188 2269 204
rect 2235 -204 2269 -188
rect -2223 -272 -2207 -238
rect -1839 -272 -1823 -238
rect -1645 -272 -1629 -238
rect -1261 -272 -1245 -238
rect -1067 -272 -1051 -238
rect -683 -272 -667 -238
rect -489 -272 -473 -238
rect -105 -272 -89 -238
rect 89 -272 105 -238
rect 473 -272 489 -238
rect 667 -272 683 -238
rect 1051 -272 1067 -238
rect 1245 -272 1261 -238
rect 1629 -272 1645 -238
rect 1823 -272 1839 -238
rect 2207 -272 2223 -238
rect -2403 -376 -2369 -314
rect 2369 -376 2403 -314
rect -2403 -410 -2307 -376
rect 2307 -410 2403 -376
<< viali >>
rect -2207 238 -1839 272
rect -1629 238 -1261 272
rect -1051 238 -683 272
rect -473 238 -105 272
rect 105 238 473 272
rect 683 238 1051 272
rect 1261 238 1629 272
rect 1839 238 2207 272
rect -2207 -272 -1839 -238
rect -1629 -272 -1261 -238
rect -1051 -272 -683 -238
rect -473 -272 -105 -238
rect 105 -272 473 -238
rect 683 -272 1051 -238
rect 1261 -272 1629 -238
rect 1839 -272 2207 -238
<< metal1 >>
rect -2219 272 -1827 278
rect -2219 238 -2207 272
rect -1839 238 -1827 272
rect -2219 232 -1827 238
rect -1641 272 -1249 278
rect -1641 238 -1629 272
rect -1261 238 -1249 272
rect -1641 232 -1249 238
rect -1063 272 -671 278
rect -1063 238 -1051 272
rect -683 238 -671 272
rect -1063 232 -671 238
rect -485 272 -93 278
rect -485 238 -473 272
rect -105 238 -93 272
rect -485 232 -93 238
rect 93 272 485 278
rect 93 238 105 272
rect 473 238 485 272
rect 93 232 485 238
rect 671 272 1063 278
rect 671 238 683 272
rect 1051 238 1063 272
rect 671 232 1063 238
rect 1249 272 1641 278
rect 1249 238 1261 272
rect 1629 238 1641 272
rect 1249 232 1641 238
rect 1827 272 2219 278
rect 1827 238 1839 272
rect 2207 238 2219 272
rect 1827 232 2219 238
rect -2219 -238 -1827 -232
rect -2219 -272 -2207 -238
rect -1839 -272 -1827 -238
rect -2219 -278 -1827 -272
rect -1641 -238 -1249 -232
rect -1641 -272 -1629 -238
rect -1261 -272 -1249 -238
rect -1641 -278 -1249 -272
rect -1063 -238 -671 -232
rect -1063 -272 -1051 -238
rect -683 -272 -671 -238
rect -1063 -278 -671 -272
rect -485 -238 -93 -232
rect -485 -272 -473 -238
rect -105 -272 -93 -238
rect -485 -278 -93 -272
rect 93 -238 485 -232
rect 93 -272 105 -238
rect 473 -272 485 -238
rect 93 -278 485 -272
rect 671 -238 1063 -232
rect 671 -272 683 -238
rect 1051 -272 1063 -238
rect 671 -278 1063 -272
rect 1249 -238 1641 -232
rect 1249 -272 1261 -238
rect 1629 -272 1641 -238
rect 1249 -278 1641 -272
rect 1827 -238 2219 -232
rect 1827 -272 1839 -238
rect 2207 -272 2219 -238
rect 1827 -278 2219 -272
<< properties >>
string FIXED_BBOX -2386 -393 2386 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 2 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
