magic
tech sky130A
magscale 1 2
timestamp 1712851378
<< metal3 >>
rect -1186 3012 1186 3040
rect -1186 -3012 1102 3012
rect 1166 -3012 1186 3012
rect -1186 -3040 1186 -3012
<< via3 >>
rect 1102 -3012 1166 3012
<< mimcap >>
rect -1146 2960 854 3000
rect -1146 -2960 -1106 2960
rect 814 -2960 854 2960
rect -1146 -3000 854 -2960
<< mimcapcontact >>
rect -1106 -2960 814 2960
<< metal4 >>
rect 1086 3012 1182 3028
rect -1107 2960 815 2961
rect -1107 -2960 -1106 2960
rect 814 -2960 815 2960
rect -1107 -2961 815 -2960
rect 1086 -3012 1102 3012
rect 1166 -3012 1182 3012
rect 1086 -3028 1182 -3012
<< properties >>
string FIXED_BBOX -1186 -3040 894 3040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10 l 30.0 val 615.2 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
