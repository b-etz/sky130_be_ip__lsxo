magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< error_s >>
rect 2878 -46 2893 -39
rect 2906 -46 2921 -36
rect 5016 -46 5022 -36
rect 5044 -46 5050 -36
rect 2868 -49 7198 -46
rect 241 -367 7198 -49
rect 241 -370 2931 -367
rect 1706 -500 1756 -456
rect 319 -584 372 -500
rect 402 -584 444 -500
rect 474 -584 566 -500
rect 596 -584 649 -500
rect 804 -584 856 -500
rect 886 -584 940 -500
rect 970 -584 1022 -500
rect 1090 -584 1195 -500
rect 1225 -512 1275 -500
rect 1434 -512 1552 -500
rect 1225 -584 1290 -512
rect 1320 -584 1386 -512
rect 1416 -584 1552 -512
rect 1582 -584 1624 -500
rect 1654 -584 1756 -500
rect 1786 -512 1840 -456
rect 2010 -512 2060 -500
rect 1786 -584 1855 -512
rect 1885 -584 1964 -512
rect 1994 -584 2060 -512
rect 2090 -584 2209 -500
rect 2239 -584 2300 -500
rect 2330 -584 2382 -500
rect 2436 -584 2488 -454
rect 2518 -584 2570 -454
rect 2721 -500 2773 -454
rect 2624 -584 2676 -500
rect 2706 -584 2773 -500
rect 2803 -584 2855 -454
rect 3835 -497 3885 -453
rect 2878 -614 2893 -583
rect 2872 -648 2893 -614
rect 2878 -679 2893 -648
rect 2906 -611 2921 -580
rect 2933 -581 2985 -497
rect 3015 -581 3069 -497
rect 3099 -581 3151 -497
rect 3219 -581 3324 -497
rect 3354 -509 3404 -497
rect 3563 -509 3681 -497
rect 3354 -581 3419 -509
rect 3449 -581 3515 -509
rect 3545 -581 3681 -509
rect 3711 -581 3753 -497
rect 3783 -581 3885 -497
rect 3915 -509 3969 -453
rect 4139 -509 4189 -497
rect 3915 -581 3984 -509
rect 4014 -581 4093 -509
rect 4123 -581 4189 -509
rect 4219 -581 4338 -497
rect 4368 -581 4429 -497
rect 4459 -581 4511 -497
rect 4565 -581 4617 -451
rect 4647 -581 4699 -451
rect 4850 -497 4902 -451
rect 4753 -581 4805 -497
rect 4835 -581 4902 -497
rect 4932 -581 4984 -451
rect 5973 -497 6023 -453
rect 5016 -611 5022 -580
rect 2906 -645 2927 -611
rect 5010 -645 5022 -611
rect 2906 -676 2921 -645
rect 5016 -676 5022 -645
rect 5044 -611 5050 -580
rect 5071 -581 5123 -497
rect 5153 -581 5207 -497
rect 5237 -581 5289 -497
rect 5357 -581 5462 -497
rect 5492 -509 5542 -497
rect 5701 -509 5819 -497
rect 5492 -581 5557 -509
rect 5587 -581 5653 -509
rect 5683 -581 5819 -509
rect 5849 -581 5891 -497
rect 5921 -581 6023 -497
rect 6053 -509 6107 -453
rect 6277 -509 6327 -497
rect 6053 -581 6122 -509
rect 6152 -581 6231 -509
rect 6261 -581 6327 -509
rect 6357 -581 6476 -497
rect 6506 -581 6567 -497
rect 6597 -581 6649 -497
rect 6703 -581 6755 -451
rect 6785 -581 6837 -451
rect 6988 -497 7040 -451
rect 6891 -581 6943 -497
rect 6973 -581 7040 -497
rect 7070 -581 7122 -451
rect 5044 -645 5056 -611
rect 5044 -676 5050 -645
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_sc_hd__and2_0  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 279 0 1 -631
box -38 -48 498 592
use sky130_fd_sc_hd__dfrbp_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 777 0 1 -631
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  x3
timestamp 1707688321
transform 1 0 2906 0 1 -628
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  x4
timestamp 1707688321
transform 1 0 5044 0 1 -628
box -38 -48 2154 592
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 128 0 0 0 dvdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 128 0 0 0 dvss
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 128 0 0 0 clkin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 128 0 0 0 done
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 128 0 0 0 doneb
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 128 0 0 0 ena
port 5 nsew
<< end >>
