magic
tech sky130A
timestamp 1712544943
<< metal1 >>
rect 436 61 536 161
rect 2344 -48 2444 52
rect 446 -219 546 -119
rect 4492 -127 4592 -27
rect 444 -812 544 -712
rect 489 -1031 589 -931
rect 2349 -1523 2449 -1423
use ripple_dly_4  x1
timestamp 1712544943
transform 1 0 505 0 1 -38
box 116 -613 3637 -293
use ripple_dly_4  x2
timestamp 1712544943
transform 1 0 506 0 -1 -1542
box 116 -613 3637 -293
use sky130_fd_sc_hd__a221o_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 708 0 1 3
box -19 -24 387 296
use sky130_fd_sc_hd__einvn_0  x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 1114 0 1 3
box -19 -24 203 296
use sky130_fd_pr__nfet_01v8_AHZR5K  XM3
timestamp 1712071977
transform 1 0 4008 0 1 -51
box -298 -130 298 130
<< labels >>
flabel metal1 2344 -48 2444 52 0 FreeSans 64 0 0 0 dvdd
port 0 nsew
flabel metal1 2349 -1523 2449 -1423 0 FreeSans 64 0 0 0 dvss
port 1 nsew
flabel metal1 444 -812 544 -712 0 FreeSans 64 0 0 0 clkin
port 2 nsew
flabel metal1 4492 -127 4592 -27 0 FreeSans 64 0 0 0 clkout
port 3 nsew
flabel metal1 446 -219 546 -119 0 FreeSans 64 0 0 0 ena
port 4 nsew
flabel metal1 436 61 536 161 0 FreeSans 64 0 0 0 stby
port 6 nsew
flabel metal1 489 -1031 589 -931 0 FreeSans 64 0 0 0 stby_b
port 7 nsew
<< end >>
