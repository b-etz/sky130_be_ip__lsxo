magic
tech sky130A
magscale 1 2
timestamp 1712087189
<< nwell >>
rect -624 -697 624 697
<< mvpmos >>
rect -366 -400 -266 400
rect -208 -400 -108 400
rect -50 -400 50 400
rect 108 -400 208 400
rect 266 -400 366 400
<< mvpdiff >>
rect -424 388 -366 400
rect -424 -388 -412 388
rect -378 -388 -366 388
rect -424 -400 -366 -388
rect -266 388 -208 400
rect -266 -388 -254 388
rect -220 -388 -208 388
rect -266 -400 -208 -388
rect -108 388 -50 400
rect -108 -388 -96 388
rect -62 -388 -50 388
rect -108 -400 -50 -388
rect 50 388 108 400
rect 50 -388 62 388
rect 96 -388 108 388
rect 50 -400 108 -388
rect 208 388 266 400
rect 208 -388 220 388
rect 254 -388 266 388
rect 208 -400 266 -388
rect 366 388 424 400
rect 366 -388 378 388
rect 412 -388 424 388
rect 366 -400 424 -388
<< mvpdiffc >>
rect -412 -388 -378 388
rect -254 -388 -220 388
rect -96 -388 -62 388
rect 62 -388 96 388
rect 220 -388 254 388
rect 378 -388 412 388
<< mvnsubdiff >>
rect -558 619 558 631
rect -558 585 -450 619
rect 450 585 558 619
rect -558 573 558 585
rect -558 523 -500 573
rect -558 -523 -546 523
rect -512 -523 -500 523
rect 500 523 558 573
rect -558 -573 -500 -523
rect 500 -523 512 523
rect 546 -523 558 523
rect 500 -573 558 -523
rect -558 -585 558 -573
rect -558 -619 -450 -585
rect 450 -619 558 -585
rect -558 -631 558 -619
<< mvnsubdiffcont >>
rect -450 585 450 619
rect -546 -523 -512 523
rect 512 -523 546 523
rect -450 -619 450 -585
<< poly >>
rect -366 481 -266 497
rect -366 447 -350 481
rect -282 447 -266 481
rect -366 400 -266 447
rect -208 481 -108 497
rect -208 447 -192 481
rect -124 447 -108 481
rect -208 400 -108 447
rect -50 481 50 497
rect -50 447 -34 481
rect 34 447 50 481
rect -50 400 50 447
rect 108 481 208 497
rect 108 447 124 481
rect 192 447 208 481
rect 108 400 208 447
rect 266 481 366 497
rect 266 447 282 481
rect 350 447 366 481
rect 266 400 366 447
rect -366 -447 -266 -400
rect -366 -481 -350 -447
rect -282 -481 -266 -447
rect -366 -497 -266 -481
rect -208 -447 -108 -400
rect -208 -481 -192 -447
rect -124 -481 -108 -447
rect -208 -497 -108 -481
rect -50 -447 50 -400
rect -50 -481 -34 -447
rect 34 -481 50 -447
rect -50 -497 50 -481
rect 108 -447 208 -400
rect 108 -481 124 -447
rect 192 -481 208 -447
rect 108 -497 208 -481
rect 266 -447 366 -400
rect 266 -481 282 -447
rect 350 -481 366 -447
rect 266 -497 366 -481
<< polycont >>
rect -350 447 -282 481
rect -192 447 -124 481
rect -34 447 34 481
rect 124 447 192 481
rect 282 447 350 481
rect -350 -481 -282 -447
rect -192 -481 -124 -447
rect -34 -481 34 -447
rect 124 -481 192 -447
rect 282 -481 350 -447
<< locali >>
rect -546 585 -450 619
rect 450 585 546 619
rect -546 523 -512 585
rect 512 523 546 585
rect -366 447 -350 481
rect -282 447 -266 481
rect -208 447 -192 481
rect -124 447 -108 481
rect -50 447 -34 481
rect 34 447 50 481
rect 108 447 124 481
rect 192 447 208 481
rect 266 447 282 481
rect 350 447 366 481
rect -412 388 -378 404
rect -412 -404 -378 -388
rect -254 388 -220 404
rect -254 -404 -220 -388
rect -96 388 -62 404
rect -96 -404 -62 -388
rect 62 388 96 404
rect 62 -404 96 -388
rect 220 388 254 404
rect 220 -404 254 -388
rect 378 388 412 404
rect 378 -404 412 -388
rect -366 -481 -350 -447
rect -282 -481 -266 -447
rect -208 -481 -192 -447
rect -124 -481 -108 -447
rect -50 -481 -34 -447
rect 34 -481 50 -447
rect 108 -481 124 -447
rect 192 -481 208 -447
rect 266 -481 282 -447
rect 350 -481 366 -447
rect -546 -585 -512 -523
rect 512 -585 546 -523
rect -546 -619 -450 -585
rect 450 -619 546 -585
<< viali >>
rect -350 447 -282 481
rect -192 447 -124 481
rect -34 447 34 481
rect 124 447 192 481
rect 282 447 350 481
rect -412 -388 -378 388
rect -254 -388 -220 388
rect -96 -388 -62 388
rect 62 -388 96 388
rect 220 -388 254 388
rect 378 -388 412 388
rect -350 -481 -282 -447
rect -192 -481 -124 -447
rect -34 -481 34 -447
rect 124 -481 192 -447
rect 282 -481 350 -447
<< metal1 >>
rect -362 481 -270 487
rect -362 447 -350 481
rect -282 447 -270 481
rect -362 441 -270 447
rect -204 481 -112 487
rect -204 447 -192 481
rect -124 447 -112 481
rect -204 441 -112 447
rect -46 481 46 487
rect -46 447 -34 481
rect 34 447 46 481
rect -46 441 46 447
rect 112 481 204 487
rect 112 447 124 481
rect 192 447 204 481
rect 112 441 204 447
rect 270 481 362 487
rect 270 447 282 481
rect 350 447 362 481
rect 270 441 362 447
rect -418 388 -372 400
rect -418 -388 -412 388
rect -378 -388 -372 388
rect -418 -400 -372 -388
rect -260 388 -214 400
rect -260 -388 -254 388
rect -220 -388 -214 388
rect -260 -400 -214 -388
rect -102 388 -56 400
rect -102 -388 -96 388
rect -62 -388 -56 388
rect -102 -400 -56 -388
rect 56 388 102 400
rect 56 -388 62 388
rect 96 -388 102 388
rect 56 -400 102 -388
rect 214 388 260 400
rect 214 -388 220 388
rect 254 -388 260 388
rect 214 -400 260 -388
rect 372 388 418 400
rect 372 -388 378 388
rect 412 -388 418 388
rect 372 -400 418 -388
rect -362 -447 -270 -441
rect -362 -481 -350 -447
rect -282 -481 -270 -447
rect -362 -487 -270 -481
rect -204 -447 -112 -441
rect -204 -481 -192 -447
rect -124 -481 -112 -447
rect -204 -487 -112 -481
rect -46 -447 46 -441
rect -46 -481 -34 -447
rect 34 -481 46 -447
rect -46 -487 46 -481
rect 112 -447 204 -441
rect 112 -481 124 -447
rect 192 -481 204 -447
rect 112 -487 204 -481
rect 270 -447 362 -441
rect 270 -481 282 -447
rect 350 -481 362 -447
rect 270 -487 362 -481
<< properties >>
string FIXED_BBOX -529 -602 529 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 0.5 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
