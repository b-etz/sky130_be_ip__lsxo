magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< pwell >>
rect -428 -2185 428 2185
<< mvnmos >>
rect -200 1127 200 1927
rect -200 109 200 909
rect -200 -909 200 -109
rect -200 -1927 200 -1127
<< mvndiff >>
rect -258 1915 -200 1927
rect -258 1139 -246 1915
rect -212 1139 -200 1915
rect -258 1127 -200 1139
rect 200 1915 258 1927
rect 200 1139 212 1915
rect 246 1139 258 1915
rect 200 1127 258 1139
rect -258 897 -200 909
rect -258 121 -246 897
rect -212 121 -200 897
rect -258 109 -200 121
rect 200 897 258 909
rect 200 121 212 897
rect 246 121 258 897
rect 200 109 258 121
rect -258 -121 -200 -109
rect -258 -897 -246 -121
rect -212 -897 -200 -121
rect -258 -909 -200 -897
rect 200 -121 258 -109
rect 200 -897 212 -121
rect 246 -897 258 -121
rect 200 -909 258 -897
rect -258 -1139 -200 -1127
rect -258 -1915 -246 -1139
rect -212 -1915 -200 -1139
rect -258 -1927 -200 -1915
rect 200 -1139 258 -1127
rect 200 -1915 212 -1139
rect 246 -1915 258 -1139
rect 200 -1927 258 -1915
<< mvndiffc >>
rect -246 1139 -212 1915
rect 212 1139 246 1915
rect -246 121 -212 897
rect 212 121 246 897
rect -246 -897 -212 -121
rect 212 -897 246 -121
rect -246 -1915 -212 -1139
rect 212 -1915 246 -1139
<< mvpsubdiff >>
rect -392 2137 392 2149
rect -392 2103 -284 2137
rect 284 2103 392 2137
rect -392 2091 392 2103
rect -392 2041 -334 2091
rect -392 -2041 -380 2041
rect -346 -2041 -334 2041
rect 334 2041 392 2091
rect -392 -2091 -334 -2041
rect 334 -2041 346 2041
rect 380 -2041 392 2041
rect 334 -2091 392 -2041
rect -392 -2103 392 -2091
rect -392 -2137 -284 -2103
rect 284 -2137 392 -2103
rect -392 -2149 392 -2137
<< mvpsubdiffcont >>
rect -284 2103 284 2137
rect -380 -2041 -346 2041
rect 346 -2041 380 2041
rect -284 -2137 284 -2103
<< poly >>
rect -200 1999 200 2015
rect -200 1965 -184 1999
rect 184 1965 200 1999
rect -200 1927 200 1965
rect -200 1089 200 1127
rect -200 1055 -184 1089
rect 184 1055 200 1089
rect -200 1039 200 1055
rect -200 981 200 997
rect -200 947 -184 981
rect 184 947 200 981
rect -200 909 200 947
rect -200 71 200 109
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -109 200 -71
rect -200 -947 200 -909
rect -200 -981 -184 -947
rect 184 -981 200 -947
rect -200 -997 200 -981
rect -200 -1055 200 -1039
rect -200 -1089 -184 -1055
rect 184 -1089 200 -1055
rect -200 -1127 200 -1089
rect -200 -1965 200 -1927
rect -200 -1999 -184 -1965
rect 184 -1999 200 -1965
rect -200 -2015 200 -1999
<< polycont >>
rect -184 1965 184 1999
rect -184 1055 184 1089
rect -184 947 184 981
rect -184 37 184 71
rect -184 -71 184 -37
rect -184 -981 184 -947
rect -184 -1089 184 -1055
rect -184 -1999 184 -1965
<< locali >>
rect -380 2103 -284 2137
rect 284 2103 380 2137
rect -380 2041 -346 2103
rect 346 2041 380 2103
rect -200 1965 -184 1999
rect 184 1965 200 1999
rect -246 1915 -212 1931
rect -246 1123 -212 1139
rect 212 1915 246 1931
rect 212 1123 246 1139
rect -200 1055 -184 1089
rect 184 1055 200 1089
rect -200 947 -184 981
rect 184 947 200 981
rect -246 897 -212 913
rect -246 105 -212 121
rect 212 897 246 913
rect 212 105 246 121
rect -200 37 -184 71
rect 184 37 200 71
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -246 -121 -212 -105
rect -246 -913 -212 -897
rect 212 -121 246 -105
rect 212 -913 246 -897
rect -200 -981 -184 -947
rect 184 -981 200 -947
rect -200 -1089 -184 -1055
rect 184 -1089 200 -1055
rect -246 -1139 -212 -1123
rect -246 -1931 -212 -1915
rect 212 -1139 246 -1123
rect 212 -1931 246 -1915
rect -200 -1999 -184 -1965
rect 184 -1999 200 -1965
rect -380 -2103 -346 -2041
rect 346 -2103 380 -2041
rect -380 -2137 -284 -2103
rect 284 -2137 380 -2103
<< viali >>
rect -184 1965 184 1999
rect -246 1139 -212 1915
rect 212 1139 246 1915
rect -184 1055 184 1089
rect -184 947 184 981
rect -246 121 -212 897
rect 212 121 246 897
rect -184 37 184 71
rect -184 -71 184 -37
rect -246 -897 -212 -121
rect 212 -897 246 -121
rect -184 -981 184 -947
rect -184 -1089 184 -1055
rect -246 -1915 -212 -1139
rect 212 -1915 246 -1139
rect -184 -1999 184 -1965
<< metal1 >>
rect -196 1999 196 2005
rect -196 1965 -184 1999
rect 184 1965 196 1999
rect -196 1959 196 1965
rect -252 1915 -206 1927
rect -252 1139 -246 1915
rect -212 1139 -206 1915
rect -252 1127 -206 1139
rect 206 1915 252 1927
rect 206 1139 212 1915
rect 246 1139 252 1915
rect 206 1127 252 1139
rect -196 1089 196 1095
rect -196 1055 -184 1089
rect 184 1055 196 1089
rect -196 1049 196 1055
rect -196 981 196 987
rect -196 947 -184 981
rect 184 947 196 981
rect -196 941 196 947
rect -252 897 -206 909
rect -252 121 -246 897
rect -212 121 -206 897
rect -252 109 -206 121
rect 206 897 252 909
rect 206 121 212 897
rect 246 121 252 897
rect 206 109 252 121
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect -252 -121 -206 -109
rect -252 -897 -246 -121
rect -212 -897 -206 -121
rect -252 -909 -206 -897
rect 206 -121 252 -109
rect 206 -897 212 -121
rect 246 -897 252 -121
rect 206 -909 252 -897
rect -196 -947 196 -941
rect -196 -981 -184 -947
rect 184 -981 196 -947
rect -196 -987 196 -981
rect -196 -1055 196 -1049
rect -196 -1089 -184 -1055
rect 184 -1089 196 -1055
rect -196 -1095 196 -1089
rect -252 -1139 -206 -1127
rect -252 -1915 -246 -1139
rect -212 -1915 -206 -1139
rect -252 -1927 -206 -1915
rect 206 -1139 252 -1127
rect 206 -1915 212 -1139
rect 246 -1915 252 -1139
rect 206 -1927 252 -1915
rect -196 -1965 196 -1959
rect -196 -1999 -184 -1965
rect 184 -1999 196 -1965
rect -196 -2005 196 -1999
<< properties >>
string FIXED_BBOX -363 -2120 363 2120
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 2.0 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
