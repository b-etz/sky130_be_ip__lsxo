magic
tech sky130A
magscale 1 2
timestamp 1712250795
<< pwell >>
rect -2193 -8582 2193 8582
<< psubdiff >>
rect -2157 8512 -2061 8546
rect 2061 8512 2157 8546
rect -2157 8450 -2123 8512
rect 2123 8450 2157 8512
rect -2157 -8512 -2123 -8450
rect 2123 -8512 2157 -8450
rect -2157 -8546 -2061 -8512
rect 2061 -8546 2157 -8512
<< psubdiffcont >>
rect -2061 8512 2061 8546
rect -2157 -8450 -2123 8450
rect 2123 -8450 2157 8450
rect -2061 -8546 2061 -8512
<< xpolycontact >>
rect -2027 7984 -1957 8416
rect -2027 -8416 -1957 -7984
rect -1861 7984 -1791 8416
rect -1861 -8416 -1791 -7984
rect -1695 7984 -1625 8416
rect -1695 -8416 -1625 -7984
rect -1529 7984 -1459 8416
rect -1529 -8416 -1459 -7984
rect -1363 7984 -1293 8416
rect -1363 -8416 -1293 -7984
rect -1197 7984 -1127 8416
rect -1197 -8416 -1127 -7984
rect -1031 7984 -961 8416
rect -1031 -8416 -961 -7984
rect -865 7984 -795 8416
rect -865 -8416 -795 -7984
rect -699 7984 -629 8416
rect -699 -8416 -629 -7984
rect -533 7984 -463 8416
rect -533 -8416 -463 -7984
rect -367 7984 -297 8416
rect -367 -8416 -297 -7984
rect -201 7984 -131 8416
rect -201 -8416 -131 -7984
rect -35 7984 35 8416
rect -35 -8416 35 -7984
rect 131 7984 201 8416
rect 131 -8416 201 -7984
rect 297 7984 367 8416
rect 297 -8416 367 -7984
rect 463 7984 533 8416
rect 463 -8416 533 -7984
rect 629 7984 699 8416
rect 629 -8416 699 -7984
rect 795 7984 865 8416
rect 795 -8416 865 -7984
rect 961 7984 1031 8416
rect 961 -8416 1031 -7984
rect 1127 7984 1197 8416
rect 1127 -8416 1197 -7984
rect 1293 7984 1363 8416
rect 1293 -8416 1363 -7984
rect 1459 7984 1529 8416
rect 1459 -8416 1529 -7984
rect 1625 7984 1695 8416
rect 1625 -8416 1695 -7984
rect 1791 7984 1861 8416
rect 1791 -8416 1861 -7984
rect 1957 7984 2027 8416
rect 1957 -8416 2027 -7984
<< xpolyres >>
rect -2027 -7984 -1957 7984
rect -1861 -7984 -1791 7984
rect -1695 -7984 -1625 7984
rect -1529 -7984 -1459 7984
rect -1363 -7984 -1293 7984
rect -1197 -7984 -1127 7984
rect -1031 -7984 -961 7984
rect -865 -7984 -795 7984
rect -699 -7984 -629 7984
rect -533 -7984 -463 7984
rect -367 -7984 -297 7984
rect -201 -7984 -131 7984
rect -35 -7984 35 7984
rect 131 -7984 201 7984
rect 297 -7984 367 7984
rect 463 -7984 533 7984
rect 629 -7984 699 7984
rect 795 -7984 865 7984
rect 961 -7984 1031 7984
rect 1127 -7984 1197 7984
rect 1293 -7984 1363 7984
rect 1459 -7984 1529 7984
rect 1625 -7984 1695 7984
rect 1791 -7984 1861 7984
rect 1957 -7984 2027 7984
<< locali >>
rect -2157 8512 -2061 8546
rect 2061 8512 2157 8546
rect -2157 8450 -2123 8512
rect 2123 8450 2157 8512
rect -2157 -8512 -2123 -8450
rect 2123 -8512 2157 -8450
rect -2157 -8546 -2061 -8512
rect 2061 -8546 2157 -8512
<< viali >>
rect -2011 8001 -1973 8398
rect -1845 8001 -1807 8398
rect -1679 8001 -1641 8398
rect -1513 8001 -1475 8398
rect -1347 8001 -1309 8398
rect -1181 8001 -1143 8398
rect -1015 8001 -977 8398
rect -849 8001 -811 8398
rect -683 8001 -645 8398
rect -517 8001 -479 8398
rect -351 8001 -313 8398
rect -185 8001 -147 8398
rect -19 8001 19 8398
rect 147 8001 185 8398
rect 313 8001 351 8398
rect 479 8001 517 8398
rect 645 8001 683 8398
rect 811 8001 849 8398
rect 977 8001 1015 8398
rect 1143 8001 1181 8398
rect 1309 8001 1347 8398
rect 1475 8001 1513 8398
rect 1641 8001 1679 8398
rect 1807 8001 1845 8398
rect 1973 8001 2011 8398
rect -2011 -8398 -1973 -8001
rect -1845 -8398 -1807 -8001
rect -1679 -8398 -1641 -8001
rect -1513 -8398 -1475 -8001
rect -1347 -8398 -1309 -8001
rect -1181 -8398 -1143 -8001
rect -1015 -8398 -977 -8001
rect -849 -8398 -811 -8001
rect -683 -8398 -645 -8001
rect -517 -8398 -479 -8001
rect -351 -8398 -313 -8001
rect -185 -8398 -147 -8001
rect -19 -8398 19 -8001
rect 147 -8398 185 -8001
rect 313 -8398 351 -8001
rect 479 -8398 517 -8001
rect 645 -8398 683 -8001
rect 811 -8398 849 -8001
rect 977 -8398 1015 -8001
rect 1143 -8398 1181 -8001
rect 1309 -8398 1347 -8001
rect 1475 -8398 1513 -8001
rect 1641 -8398 1679 -8001
rect 1807 -8398 1845 -8001
rect 1973 -8398 2011 -8001
<< metal1 >>
rect -2017 8398 -1967 8410
rect -2017 8001 -2011 8398
rect -1973 8001 -1967 8398
rect -2017 7989 -1967 8001
rect -1851 8398 -1801 8410
rect -1851 8001 -1845 8398
rect -1807 8001 -1801 8398
rect -1851 7989 -1801 8001
rect -1685 8398 -1635 8410
rect -1685 8001 -1679 8398
rect -1641 8001 -1635 8398
rect -1685 7989 -1635 8001
rect -1519 8398 -1469 8410
rect -1519 8001 -1513 8398
rect -1475 8001 -1469 8398
rect -1519 7989 -1469 8001
rect -1353 8398 -1303 8410
rect -1353 8001 -1347 8398
rect -1309 8001 -1303 8398
rect -1353 7989 -1303 8001
rect -1187 8398 -1137 8410
rect -1187 8001 -1181 8398
rect -1143 8001 -1137 8398
rect -1187 7989 -1137 8001
rect -1021 8398 -971 8410
rect -1021 8001 -1015 8398
rect -977 8001 -971 8398
rect -1021 7989 -971 8001
rect -855 8398 -805 8410
rect -855 8001 -849 8398
rect -811 8001 -805 8398
rect -855 7989 -805 8001
rect -689 8398 -639 8410
rect -689 8001 -683 8398
rect -645 8001 -639 8398
rect -689 7989 -639 8001
rect -523 8398 -473 8410
rect -523 8001 -517 8398
rect -479 8001 -473 8398
rect -523 7989 -473 8001
rect -357 8398 -307 8410
rect -357 8001 -351 8398
rect -313 8001 -307 8398
rect -357 7989 -307 8001
rect -191 8398 -141 8410
rect -191 8001 -185 8398
rect -147 8001 -141 8398
rect -191 7989 -141 8001
rect -25 8398 25 8410
rect -25 8001 -19 8398
rect 19 8001 25 8398
rect -25 7989 25 8001
rect 141 8398 191 8410
rect 141 8001 147 8398
rect 185 8001 191 8398
rect 141 7989 191 8001
rect 307 8398 357 8410
rect 307 8001 313 8398
rect 351 8001 357 8398
rect 307 7989 357 8001
rect 473 8398 523 8410
rect 473 8001 479 8398
rect 517 8001 523 8398
rect 473 7989 523 8001
rect 639 8398 689 8410
rect 639 8001 645 8398
rect 683 8001 689 8398
rect 639 7989 689 8001
rect 805 8398 855 8410
rect 805 8001 811 8398
rect 849 8001 855 8398
rect 805 7989 855 8001
rect 971 8398 1021 8410
rect 971 8001 977 8398
rect 1015 8001 1021 8398
rect 971 7989 1021 8001
rect 1137 8398 1187 8410
rect 1137 8001 1143 8398
rect 1181 8001 1187 8398
rect 1137 7989 1187 8001
rect 1303 8398 1353 8410
rect 1303 8001 1309 8398
rect 1347 8001 1353 8398
rect 1303 7989 1353 8001
rect 1469 8398 1519 8410
rect 1469 8001 1475 8398
rect 1513 8001 1519 8398
rect 1469 7989 1519 8001
rect 1635 8398 1685 8410
rect 1635 8001 1641 8398
rect 1679 8001 1685 8398
rect 1635 7989 1685 8001
rect 1801 8398 1851 8410
rect 1801 8001 1807 8398
rect 1845 8001 1851 8398
rect 1801 7989 1851 8001
rect 1967 8398 2017 8410
rect 1967 8001 1973 8398
rect 2011 8001 2017 8398
rect 1967 7989 2017 8001
rect -2017 -8001 -1967 -7989
rect -2017 -8398 -2011 -8001
rect -1973 -8398 -1967 -8001
rect -2017 -8410 -1967 -8398
rect -1851 -8001 -1801 -7989
rect -1851 -8398 -1845 -8001
rect -1807 -8398 -1801 -8001
rect -1851 -8410 -1801 -8398
rect -1685 -8001 -1635 -7989
rect -1685 -8398 -1679 -8001
rect -1641 -8398 -1635 -8001
rect -1685 -8410 -1635 -8398
rect -1519 -8001 -1469 -7989
rect -1519 -8398 -1513 -8001
rect -1475 -8398 -1469 -8001
rect -1519 -8410 -1469 -8398
rect -1353 -8001 -1303 -7989
rect -1353 -8398 -1347 -8001
rect -1309 -8398 -1303 -8001
rect -1353 -8410 -1303 -8398
rect -1187 -8001 -1137 -7989
rect -1187 -8398 -1181 -8001
rect -1143 -8398 -1137 -8001
rect -1187 -8410 -1137 -8398
rect -1021 -8001 -971 -7989
rect -1021 -8398 -1015 -8001
rect -977 -8398 -971 -8001
rect -1021 -8410 -971 -8398
rect -855 -8001 -805 -7989
rect -855 -8398 -849 -8001
rect -811 -8398 -805 -8001
rect -855 -8410 -805 -8398
rect -689 -8001 -639 -7989
rect -689 -8398 -683 -8001
rect -645 -8398 -639 -8001
rect -689 -8410 -639 -8398
rect -523 -8001 -473 -7989
rect -523 -8398 -517 -8001
rect -479 -8398 -473 -8001
rect -523 -8410 -473 -8398
rect -357 -8001 -307 -7989
rect -357 -8398 -351 -8001
rect -313 -8398 -307 -8001
rect -357 -8410 -307 -8398
rect -191 -8001 -141 -7989
rect -191 -8398 -185 -8001
rect -147 -8398 -141 -8001
rect -191 -8410 -141 -8398
rect -25 -8001 25 -7989
rect -25 -8398 -19 -8001
rect 19 -8398 25 -8001
rect -25 -8410 25 -8398
rect 141 -8001 191 -7989
rect 141 -8398 147 -8001
rect 185 -8398 191 -8001
rect 141 -8410 191 -8398
rect 307 -8001 357 -7989
rect 307 -8398 313 -8001
rect 351 -8398 357 -8001
rect 307 -8410 357 -8398
rect 473 -8001 523 -7989
rect 473 -8398 479 -8001
rect 517 -8398 523 -8001
rect 473 -8410 523 -8398
rect 639 -8001 689 -7989
rect 639 -8398 645 -8001
rect 683 -8398 689 -8001
rect 639 -8410 689 -8398
rect 805 -8001 855 -7989
rect 805 -8398 811 -8001
rect 849 -8398 855 -8001
rect 805 -8410 855 -8398
rect 971 -8001 1021 -7989
rect 971 -8398 977 -8001
rect 1015 -8398 1021 -8001
rect 971 -8410 1021 -8398
rect 1137 -8001 1187 -7989
rect 1137 -8398 1143 -8001
rect 1181 -8398 1187 -8001
rect 1137 -8410 1187 -8398
rect 1303 -8001 1353 -7989
rect 1303 -8398 1309 -8001
rect 1347 -8398 1353 -8001
rect 1303 -8410 1353 -8398
rect 1469 -8001 1519 -7989
rect 1469 -8398 1475 -8001
rect 1513 -8398 1519 -8001
rect 1469 -8410 1519 -8398
rect 1635 -8001 1685 -7989
rect 1635 -8398 1641 -8001
rect 1679 -8398 1685 -8001
rect 1635 -8410 1685 -8398
rect 1801 -8001 1851 -7989
rect 1801 -8398 1807 -8001
rect 1845 -8398 1851 -8001
rect 1801 -8410 1851 -8398
rect 1967 -8001 2017 -7989
rect 1967 -8398 1973 -8001
rect 2011 -8398 2017 -8001
rect 1967 -8410 2017 -8398
<< properties >>
string FIXED_BBOX -2140 -8529 2140 8529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 80 m 1 nx 25 wmin 0.350 lmin 0.50 rho 2000 val 458.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
