magic
tech sky130A
magscale 1 2
timestamp 1713142410
<< pwell >>
rect -450 -8082 450 8082
<< psubdiff >>
rect -414 8012 -318 8046
rect 318 8012 414 8046
rect -414 7950 -380 8012
rect 380 7950 414 8012
rect -414 -8012 -380 -7950
rect 380 -8012 414 -7950
rect -414 -8046 -318 -8012
rect 318 -8046 414 -8012
<< psubdiffcont >>
rect -318 8012 318 8046
rect -414 -7950 -380 7950
rect 380 -7950 414 7950
rect -318 -8046 318 -8012
<< xpolycontact >>
rect -284 7484 -214 7916
rect -284 -7916 -214 -7484
rect -118 7484 -48 7916
rect -118 -7916 -48 -7484
rect 48 7484 118 7916
rect 48 -7916 118 -7484
rect 214 7484 284 7916
rect 214 -7916 284 -7484
<< xpolyres >>
rect -284 -7484 -214 7484
rect -118 -7484 -48 7484
rect 48 -7484 118 7484
rect 214 -7484 284 7484
<< locali >>
rect -414 8012 -318 8046
rect 318 8012 414 8046
rect -414 7950 -380 8012
rect 380 7950 414 8012
rect -414 -8012 -380 -7950
rect 380 -8012 414 -7950
rect -414 -8046 -318 -8012
rect 318 -8046 414 -8012
<< viali >>
rect -268 7501 -230 7898
rect -102 7501 -64 7898
rect 64 7501 102 7898
rect 230 7501 268 7898
rect -268 -7898 -230 -7501
rect -102 -7898 -64 -7501
rect 64 -7898 102 -7501
rect 230 -7898 268 -7501
<< metal1 >>
rect -274 7898 -224 7910
rect -274 7501 -268 7898
rect -230 7501 -224 7898
rect -274 7489 -224 7501
rect -108 7898 -58 7910
rect -108 7501 -102 7898
rect -64 7501 -58 7898
rect -108 7489 -58 7501
rect 58 7898 108 7910
rect 58 7501 64 7898
rect 102 7501 108 7898
rect 58 7489 108 7501
rect 224 7898 274 7910
rect 224 7501 230 7898
rect 268 7501 274 7898
rect 224 7489 274 7501
rect -274 -7501 -224 -7489
rect -274 -7898 -268 -7501
rect -230 -7898 -224 -7501
rect -274 -7910 -224 -7898
rect -108 -7501 -58 -7489
rect -108 -7898 -102 -7501
rect -64 -7898 -58 -7501
rect -108 -7910 -58 -7898
rect 58 -7501 108 -7489
rect 58 -7898 64 -7501
rect 102 -7898 108 -7501
rect 58 -7910 108 -7898
rect 224 -7501 274 -7489
rect 224 -7898 230 -7501
rect 268 -7898 274 -7501
rect 224 -7910 274 -7898
<< properties >>
string FIXED_BBOX -397 -8029 397 8029
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 75 m 1 nx 4 wmin 0.350 lmin 0.50 rho 2000 val 429.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
