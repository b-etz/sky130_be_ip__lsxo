magic
tech sky130A
timestamp 1712071977
<< pwell >>
rect -214 -229 214 229
<< mvnmos >>
rect -100 -100 100 100
<< mvndiff >>
rect -129 94 -100 100
rect -129 -94 -123 94
rect -106 -94 -100 94
rect -129 -100 -100 -94
rect 100 94 129 100
rect 100 -94 106 94
rect 123 -94 129 94
rect 100 -100 129 -94
<< mvndiffc >>
rect -123 -94 -106 94
rect 106 -94 123 94
<< mvpsubdiff >>
rect -196 205 196 211
rect -196 188 -142 205
rect 142 188 196 205
rect -196 182 196 188
rect -196 157 -167 182
rect -196 -157 -190 157
rect -173 -157 -167 157
rect 167 157 196 182
rect -196 -182 -167 -157
rect 167 -157 173 157
rect 190 -157 196 157
rect 167 -182 196 -157
rect -196 -188 196 -182
rect -196 -205 -142 -188
rect 142 -205 196 -188
rect -196 -211 196 -205
<< mvpsubdiffcont >>
rect -142 188 142 205
rect -190 -157 -173 157
rect 173 -157 190 157
rect -142 -205 142 -188
<< poly >>
rect -100 136 100 144
rect -100 119 -92 136
rect 92 119 100 136
rect -100 100 100 119
rect -100 -119 100 -100
rect -100 -136 -92 -119
rect 92 -136 100 -119
rect -100 -144 100 -136
<< polycont >>
rect -92 119 92 136
rect -92 -136 92 -119
<< locali >>
rect -190 188 -142 205
rect 142 188 190 205
rect -190 157 -173 188
rect 173 157 190 188
rect -100 119 -92 136
rect 92 119 100 136
rect -123 94 -106 102
rect -123 -102 -106 -94
rect 106 94 123 102
rect 106 -102 123 -94
rect -100 -136 -92 -119
rect 92 -136 100 -119
rect -190 -188 -173 -157
rect 173 -188 190 -157
rect -190 -205 -142 -188
rect 142 -205 190 -188
<< viali >>
rect -92 119 92 136
rect -123 -94 -106 94
rect 106 -94 123 94
rect -92 -136 92 -119
<< metal1 >>
rect -98 136 98 139
rect -98 119 -92 136
rect 92 119 98 136
rect -98 116 98 119
rect -126 94 -103 100
rect -126 -94 -123 94
rect -106 -94 -103 94
rect -126 -100 -103 -94
rect 103 94 126 100
rect 103 -94 106 94
rect 123 -94 126 94
rect 103 -100 126 -94
rect -98 -119 98 -116
rect -98 -136 -92 -119
rect 92 -136 98 -119
rect -98 -139 98 -136
<< properties >>
string FIXED_BBOX -181 -196 181 196
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
