magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< metal4 >>
rect -1349 35839 1349 35880
rect -1349 33761 1093 35839
rect 1329 33761 1349 35839
rect -1349 33720 1349 33761
rect -1349 33439 1349 33480
rect -1349 31361 1093 33439
rect 1329 31361 1349 33439
rect -1349 31320 1349 31361
rect -1349 31039 1349 31080
rect -1349 28961 1093 31039
rect 1329 28961 1349 31039
rect -1349 28920 1349 28961
rect -1349 28639 1349 28680
rect -1349 26561 1093 28639
rect 1329 26561 1349 28639
rect -1349 26520 1349 26561
rect -1349 26239 1349 26280
rect -1349 24161 1093 26239
rect 1329 24161 1349 26239
rect -1349 24120 1349 24161
rect -1349 23839 1349 23880
rect -1349 21761 1093 23839
rect 1329 21761 1349 23839
rect -1349 21720 1349 21761
rect -1349 21439 1349 21480
rect -1349 19361 1093 21439
rect 1329 19361 1349 21439
rect -1349 19320 1349 19361
rect -1349 19039 1349 19080
rect -1349 16961 1093 19039
rect 1329 16961 1349 19039
rect -1349 16920 1349 16961
rect -1349 16639 1349 16680
rect -1349 14561 1093 16639
rect 1329 14561 1349 16639
rect -1349 14520 1349 14561
rect -1349 14239 1349 14280
rect -1349 12161 1093 14239
rect 1329 12161 1349 14239
rect -1349 12120 1349 12161
rect -1349 11839 1349 11880
rect -1349 9761 1093 11839
rect 1329 9761 1349 11839
rect -1349 9720 1349 9761
rect -1349 9439 1349 9480
rect -1349 7361 1093 9439
rect 1329 7361 1349 9439
rect -1349 7320 1349 7361
rect -1349 7039 1349 7080
rect -1349 4961 1093 7039
rect 1329 4961 1349 7039
rect -1349 4920 1349 4961
rect -1349 4639 1349 4680
rect -1349 2561 1093 4639
rect 1329 2561 1349 4639
rect -1349 2520 1349 2561
rect -1349 2239 1349 2280
rect -1349 161 1093 2239
rect 1329 161 1349 2239
rect -1349 120 1349 161
rect -1349 -161 1349 -120
rect -1349 -2239 1093 -161
rect 1329 -2239 1349 -161
rect -1349 -2280 1349 -2239
rect -1349 -2561 1349 -2520
rect -1349 -4639 1093 -2561
rect 1329 -4639 1349 -2561
rect -1349 -4680 1349 -4639
rect -1349 -4961 1349 -4920
rect -1349 -7039 1093 -4961
rect 1329 -7039 1349 -4961
rect -1349 -7080 1349 -7039
rect -1349 -7361 1349 -7320
rect -1349 -9439 1093 -7361
rect 1329 -9439 1349 -7361
rect -1349 -9480 1349 -9439
rect -1349 -9761 1349 -9720
rect -1349 -11839 1093 -9761
rect 1329 -11839 1349 -9761
rect -1349 -11880 1349 -11839
rect -1349 -12161 1349 -12120
rect -1349 -14239 1093 -12161
rect 1329 -14239 1349 -12161
rect -1349 -14280 1349 -14239
rect -1349 -14561 1349 -14520
rect -1349 -16639 1093 -14561
rect 1329 -16639 1349 -14561
rect -1349 -16680 1349 -16639
rect -1349 -16961 1349 -16920
rect -1349 -19039 1093 -16961
rect 1329 -19039 1349 -16961
rect -1349 -19080 1349 -19039
rect -1349 -19361 1349 -19320
rect -1349 -21439 1093 -19361
rect 1329 -21439 1349 -19361
rect -1349 -21480 1349 -21439
rect -1349 -21761 1349 -21720
rect -1349 -23839 1093 -21761
rect 1329 -23839 1349 -21761
rect -1349 -23880 1349 -23839
rect -1349 -24161 1349 -24120
rect -1349 -26239 1093 -24161
rect 1329 -26239 1349 -24161
rect -1349 -26280 1349 -26239
rect -1349 -26561 1349 -26520
rect -1349 -28639 1093 -26561
rect 1329 -28639 1349 -26561
rect -1349 -28680 1349 -28639
rect -1349 -28961 1349 -28920
rect -1349 -31039 1093 -28961
rect 1329 -31039 1349 -28961
rect -1349 -31080 1349 -31039
rect -1349 -31361 1349 -31320
rect -1349 -33439 1093 -31361
rect 1329 -33439 1349 -31361
rect -1349 -33480 1349 -33439
rect -1349 -33761 1349 -33720
rect -1349 -35839 1093 -33761
rect 1329 -35839 1349 -33761
rect -1349 -35880 1349 -35839
<< via4 >>
rect 1093 33761 1329 35839
rect 1093 31361 1329 33439
rect 1093 28961 1329 31039
rect 1093 26561 1329 28639
rect 1093 24161 1329 26239
rect 1093 21761 1329 23839
rect 1093 19361 1329 21439
rect 1093 16961 1329 19039
rect 1093 14561 1329 16639
rect 1093 12161 1329 14239
rect 1093 9761 1329 11839
rect 1093 7361 1329 9439
rect 1093 4961 1329 7039
rect 1093 2561 1329 4639
rect 1093 161 1329 2239
rect 1093 -2239 1329 -161
rect 1093 -4639 1329 -2561
rect 1093 -7039 1329 -4961
rect 1093 -9439 1329 -7361
rect 1093 -11839 1329 -9761
rect 1093 -14239 1329 -12161
rect 1093 -16639 1329 -14561
rect 1093 -19039 1329 -16961
rect 1093 -21439 1329 -19361
rect 1093 -23839 1329 -21761
rect 1093 -26239 1329 -24161
rect 1093 -28639 1329 -26561
rect 1093 -31039 1329 -28961
rect 1093 -33439 1329 -31361
rect 1093 -35839 1329 -33761
<< mimcap2 >>
rect -1269 35760 731 35800
rect -1269 33840 -1229 35760
rect 691 33840 731 35760
rect -1269 33800 731 33840
rect -1269 33360 731 33400
rect -1269 31440 -1229 33360
rect 691 31440 731 33360
rect -1269 31400 731 31440
rect -1269 30960 731 31000
rect -1269 29040 -1229 30960
rect 691 29040 731 30960
rect -1269 29000 731 29040
rect -1269 28560 731 28600
rect -1269 26640 -1229 28560
rect 691 26640 731 28560
rect -1269 26600 731 26640
rect -1269 26160 731 26200
rect -1269 24240 -1229 26160
rect 691 24240 731 26160
rect -1269 24200 731 24240
rect -1269 23760 731 23800
rect -1269 21840 -1229 23760
rect 691 21840 731 23760
rect -1269 21800 731 21840
rect -1269 21360 731 21400
rect -1269 19440 -1229 21360
rect 691 19440 731 21360
rect -1269 19400 731 19440
rect -1269 18960 731 19000
rect -1269 17040 -1229 18960
rect 691 17040 731 18960
rect -1269 17000 731 17040
rect -1269 16560 731 16600
rect -1269 14640 -1229 16560
rect 691 14640 731 16560
rect -1269 14600 731 14640
rect -1269 14160 731 14200
rect -1269 12240 -1229 14160
rect 691 12240 731 14160
rect -1269 12200 731 12240
rect -1269 11760 731 11800
rect -1269 9840 -1229 11760
rect 691 9840 731 11760
rect -1269 9800 731 9840
rect -1269 9360 731 9400
rect -1269 7440 -1229 9360
rect 691 7440 731 9360
rect -1269 7400 731 7440
rect -1269 6960 731 7000
rect -1269 5040 -1229 6960
rect 691 5040 731 6960
rect -1269 5000 731 5040
rect -1269 4560 731 4600
rect -1269 2640 -1229 4560
rect 691 2640 731 4560
rect -1269 2600 731 2640
rect -1269 2160 731 2200
rect -1269 240 -1229 2160
rect 691 240 731 2160
rect -1269 200 731 240
rect -1269 -240 731 -200
rect -1269 -2160 -1229 -240
rect 691 -2160 731 -240
rect -1269 -2200 731 -2160
rect -1269 -2640 731 -2600
rect -1269 -4560 -1229 -2640
rect 691 -4560 731 -2640
rect -1269 -4600 731 -4560
rect -1269 -5040 731 -5000
rect -1269 -6960 -1229 -5040
rect 691 -6960 731 -5040
rect -1269 -7000 731 -6960
rect -1269 -7440 731 -7400
rect -1269 -9360 -1229 -7440
rect 691 -9360 731 -7440
rect -1269 -9400 731 -9360
rect -1269 -9840 731 -9800
rect -1269 -11760 -1229 -9840
rect 691 -11760 731 -9840
rect -1269 -11800 731 -11760
rect -1269 -12240 731 -12200
rect -1269 -14160 -1229 -12240
rect 691 -14160 731 -12240
rect -1269 -14200 731 -14160
rect -1269 -14640 731 -14600
rect -1269 -16560 -1229 -14640
rect 691 -16560 731 -14640
rect -1269 -16600 731 -16560
rect -1269 -17040 731 -17000
rect -1269 -18960 -1229 -17040
rect 691 -18960 731 -17040
rect -1269 -19000 731 -18960
rect -1269 -19440 731 -19400
rect -1269 -21360 -1229 -19440
rect 691 -21360 731 -19440
rect -1269 -21400 731 -21360
rect -1269 -21840 731 -21800
rect -1269 -23760 -1229 -21840
rect 691 -23760 731 -21840
rect -1269 -23800 731 -23760
rect -1269 -24240 731 -24200
rect -1269 -26160 -1229 -24240
rect 691 -26160 731 -24240
rect -1269 -26200 731 -26160
rect -1269 -26640 731 -26600
rect -1269 -28560 -1229 -26640
rect 691 -28560 731 -26640
rect -1269 -28600 731 -28560
rect -1269 -29040 731 -29000
rect -1269 -30960 -1229 -29040
rect 691 -30960 731 -29040
rect -1269 -31000 731 -30960
rect -1269 -31440 731 -31400
rect -1269 -33360 -1229 -31440
rect 691 -33360 731 -31440
rect -1269 -33400 731 -33360
rect -1269 -33840 731 -33800
rect -1269 -35760 -1229 -33840
rect 691 -35760 731 -33840
rect -1269 -35800 731 -35760
<< mimcap2contact >>
rect -1229 33840 691 35760
rect -1229 31440 691 33360
rect -1229 29040 691 30960
rect -1229 26640 691 28560
rect -1229 24240 691 26160
rect -1229 21840 691 23760
rect -1229 19440 691 21360
rect -1229 17040 691 18960
rect -1229 14640 691 16560
rect -1229 12240 691 14160
rect -1229 9840 691 11760
rect -1229 7440 691 9360
rect -1229 5040 691 6960
rect -1229 2640 691 4560
rect -1229 240 691 2160
rect -1229 -2160 691 -240
rect -1229 -4560 691 -2640
rect -1229 -6960 691 -5040
rect -1229 -9360 691 -7440
rect -1229 -11760 691 -9840
rect -1229 -14160 691 -12240
rect -1229 -16560 691 -14640
rect -1229 -18960 691 -17040
rect -1229 -21360 691 -19440
rect -1229 -23760 691 -21840
rect -1229 -26160 691 -24240
rect -1229 -28560 691 -26640
rect -1229 -30960 691 -29040
rect -1229 -33360 691 -31440
rect -1229 -35760 691 -33840
<< metal5 >>
rect -429 35784 -109 36000
rect 1051 35839 1371 36000
rect -1253 35760 715 35784
rect -1253 33840 -1229 35760
rect 691 33840 715 35760
rect -1253 33816 715 33840
rect -429 33384 -109 33816
rect 1051 33761 1093 35839
rect 1329 33761 1371 35839
rect 1051 33439 1371 33761
rect -1253 33360 715 33384
rect -1253 31440 -1229 33360
rect 691 31440 715 33360
rect -1253 31416 715 31440
rect -429 30984 -109 31416
rect 1051 31361 1093 33439
rect 1329 31361 1371 33439
rect 1051 31039 1371 31361
rect -1253 30960 715 30984
rect -1253 29040 -1229 30960
rect 691 29040 715 30960
rect -1253 29016 715 29040
rect -429 28584 -109 29016
rect 1051 28961 1093 31039
rect 1329 28961 1371 31039
rect 1051 28639 1371 28961
rect -1253 28560 715 28584
rect -1253 26640 -1229 28560
rect 691 26640 715 28560
rect -1253 26616 715 26640
rect -429 26184 -109 26616
rect 1051 26561 1093 28639
rect 1329 26561 1371 28639
rect 1051 26239 1371 26561
rect -1253 26160 715 26184
rect -1253 24240 -1229 26160
rect 691 24240 715 26160
rect -1253 24216 715 24240
rect -429 23784 -109 24216
rect 1051 24161 1093 26239
rect 1329 24161 1371 26239
rect 1051 23839 1371 24161
rect -1253 23760 715 23784
rect -1253 21840 -1229 23760
rect 691 21840 715 23760
rect -1253 21816 715 21840
rect -429 21384 -109 21816
rect 1051 21761 1093 23839
rect 1329 21761 1371 23839
rect 1051 21439 1371 21761
rect -1253 21360 715 21384
rect -1253 19440 -1229 21360
rect 691 19440 715 21360
rect -1253 19416 715 19440
rect -429 18984 -109 19416
rect 1051 19361 1093 21439
rect 1329 19361 1371 21439
rect 1051 19039 1371 19361
rect -1253 18960 715 18984
rect -1253 17040 -1229 18960
rect 691 17040 715 18960
rect -1253 17016 715 17040
rect -429 16584 -109 17016
rect 1051 16961 1093 19039
rect 1329 16961 1371 19039
rect 1051 16639 1371 16961
rect -1253 16560 715 16584
rect -1253 14640 -1229 16560
rect 691 14640 715 16560
rect -1253 14616 715 14640
rect -429 14184 -109 14616
rect 1051 14561 1093 16639
rect 1329 14561 1371 16639
rect 1051 14239 1371 14561
rect -1253 14160 715 14184
rect -1253 12240 -1229 14160
rect 691 12240 715 14160
rect -1253 12216 715 12240
rect -429 11784 -109 12216
rect 1051 12161 1093 14239
rect 1329 12161 1371 14239
rect 1051 11839 1371 12161
rect -1253 11760 715 11784
rect -1253 9840 -1229 11760
rect 691 9840 715 11760
rect -1253 9816 715 9840
rect -429 9384 -109 9816
rect 1051 9761 1093 11839
rect 1329 9761 1371 11839
rect 1051 9439 1371 9761
rect -1253 9360 715 9384
rect -1253 7440 -1229 9360
rect 691 7440 715 9360
rect -1253 7416 715 7440
rect -429 6984 -109 7416
rect 1051 7361 1093 9439
rect 1329 7361 1371 9439
rect 1051 7039 1371 7361
rect -1253 6960 715 6984
rect -1253 5040 -1229 6960
rect 691 5040 715 6960
rect -1253 5016 715 5040
rect -429 4584 -109 5016
rect 1051 4961 1093 7039
rect 1329 4961 1371 7039
rect 1051 4639 1371 4961
rect -1253 4560 715 4584
rect -1253 2640 -1229 4560
rect 691 2640 715 4560
rect -1253 2616 715 2640
rect -429 2184 -109 2616
rect 1051 2561 1093 4639
rect 1329 2561 1371 4639
rect 1051 2239 1371 2561
rect -1253 2160 715 2184
rect -1253 240 -1229 2160
rect 691 240 715 2160
rect -1253 216 715 240
rect -429 -216 -109 216
rect 1051 161 1093 2239
rect 1329 161 1371 2239
rect 1051 -161 1371 161
rect -1253 -240 715 -216
rect -1253 -2160 -1229 -240
rect 691 -2160 715 -240
rect -1253 -2184 715 -2160
rect -429 -2616 -109 -2184
rect 1051 -2239 1093 -161
rect 1329 -2239 1371 -161
rect 1051 -2561 1371 -2239
rect -1253 -2640 715 -2616
rect -1253 -4560 -1229 -2640
rect 691 -4560 715 -2640
rect -1253 -4584 715 -4560
rect -429 -5016 -109 -4584
rect 1051 -4639 1093 -2561
rect 1329 -4639 1371 -2561
rect 1051 -4961 1371 -4639
rect -1253 -5040 715 -5016
rect -1253 -6960 -1229 -5040
rect 691 -6960 715 -5040
rect -1253 -6984 715 -6960
rect -429 -7416 -109 -6984
rect 1051 -7039 1093 -4961
rect 1329 -7039 1371 -4961
rect 1051 -7361 1371 -7039
rect -1253 -7440 715 -7416
rect -1253 -9360 -1229 -7440
rect 691 -9360 715 -7440
rect -1253 -9384 715 -9360
rect -429 -9816 -109 -9384
rect 1051 -9439 1093 -7361
rect 1329 -9439 1371 -7361
rect 1051 -9761 1371 -9439
rect -1253 -9840 715 -9816
rect -1253 -11760 -1229 -9840
rect 691 -11760 715 -9840
rect -1253 -11784 715 -11760
rect -429 -12216 -109 -11784
rect 1051 -11839 1093 -9761
rect 1329 -11839 1371 -9761
rect 1051 -12161 1371 -11839
rect -1253 -12240 715 -12216
rect -1253 -14160 -1229 -12240
rect 691 -14160 715 -12240
rect -1253 -14184 715 -14160
rect -429 -14616 -109 -14184
rect 1051 -14239 1093 -12161
rect 1329 -14239 1371 -12161
rect 1051 -14561 1371 -14239
rect -1253 -14640 715 -14616
rect -1253 -16560 -1229 -14640
rect 691 -16560 715 -14640
rect -1253 -16584 715 -16560
rect -429 -17016 -109 -16584
rect 1051 -16639 1093 -14561
rect 1329 -16639 1371 -14561
rect 1051 -16961 1371 -16639
rect -1253 -17040 715 -17016
rect -1253 -18960 -1229 -17040
rect 691 -18960 715 -17040
rect -1253 -18984 715 -18960
rect -429 -19416 -109 -18984
rect 1051 -19039 1093 -16961
rect 1329 -19039 1371 -16961
rect 1051 -19361 1371 -19039
rect -1253 -19440 715 -19416
rect -1253 -21360 -1229 -19440
rect 691 -21360 715 -19440
rect -1253 -21384 715 -21360
rect -429 -21816 -109 -21384
rect 1051 -21439 1093 -19361
rect 1329 -21439 1371 -19361
rect 1051 -21761 1371 -21439
rect -1253 -21840 715 -21816
rect -1253 -23760 -1229 -21840
rect 691 -23760 715 -21840
rect -1253 -23784 715 -23760
rect -429 -24216 -109 -23784
rect 1051 -23839 1093 -21761
rect 1329 -23839 1371 -21761
rect 1051 -24161 1371 -23839
rect -1253 -24240 715 -24216
rect -1253 -26160 -1229 -24240
rect 691 -26160 715 -24240
rect -1253 -26184 715 -26160
rect -429 -26616 -109 -26184
rect 1051 -26239 1093 -24161
rect 1329 -26239 1371 -24161
rect 1051 -26561 1371 -26239
rect -1253 -26640 715 -26616
rect -1253 -28560 -1229 -26640
rect 691 -28560 715 -26640
rect -1253 -28584 715 -28560
rect -429 -29016 -109 -28584
rect 1051 -28639 1093 -26561
rect 1329 -28639 1371 -26561
rect 1051 -28961 1371 -28639
rect -1253 -29040 715 -29016
rect -1253 -30960 -1229 -29040
rect 691 -30960 715 -29040
rect -1253 -30984 715 -30960
rect -429 -31416 -109 -30984
rect 1051 -31039 1093 -28961
rect 1329 -31039 1371 -28961
rect 1051 -31361 1371 -31039
rect -1253 -31440 715 -31416
rect -1253 -33360 -1229 -31440
rect 691 -33360 715 -31440
rect -1253 -33384 715 -33360
rect -429 -33816 -109 -33384
rect 1051 -33439 1093 -31361
rect 1329 -33439 1371 -31361
rect 1051 -33761 1371 -33439
rect -1253 -33840 715 -33816
rect -1253 -35760 -1229 -33840
rect 691 -35760 715 -33840
rect -1253 -35784 715 -35760
rect -429 -36000 -109 -35784
rect 1051 -35839 1093 -33761
rect 1329 -35839 1371 -33761
rect 1051 -36000 1371 -35839
<< properties >>
string FIXED_BBOX -1349 33720 811 35880
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 30 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
