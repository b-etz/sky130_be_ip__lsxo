magic
tech sky130A
magscale 1 2
timestamp 1712250795
<< metal3 >>
rect -14916 2212 -10144 2240
rect -14916 -2212 -10228 2212
rect -10164 -2212 -10144 2212
rect -14916 -2240 -10144 -2212
rect -9904 2212 -5132 2240
rect -9904 -2212 -5216 2212
rect -5152 -2212 -5132 2212
rect -9904 -2240 -5132 -2212
rect -4892 2212 -120 2240
rect -4892 -2212 -204 2212
rect -140 -2212 -120 2212
rect -4892 -2240 -120 -2212
rect 120 2212 4892 2240
rect 120 -2212 4808 2212
rect 4872 -2212 4892 2212
rect 120 -2240 4892 -2212
rect 5132 2212 9904 2240
rect 5132 -2212 9820 2212
rect 9884 -2212 9904 2212
rect 5132 -2240 9904 -2212
rect 10144 2212 14916 2240
rect 10144 -2212 14832 2212
rect 14896 -2212 14916 2212
rect 10144 -2240 14916 -2212
<< via3 >>
rect -10228 -2212 -10164 2212
rect -5216 -2212 -5152 2212
rect -204 -2212 -140 2212
rect 4808 -2212 4872 2212
rect 9820 -2212 9884 2212
rect 14832 -2212 14896 2212
<< mimcap >>
rect -14876 2160 -10476 2200
rect -14876 -2160 -14836 2160
rect -10516 -2160 -10476 2160
rect -14876 -2200 -10476 -2160
rect -9864 2160 -5464 2200
rect -9864 -2160 -9824 2160
rect -5504 -2160 -5464 2160
rect -9864 -2200 -5464 -2160
rect -4852 2160 -452 2200
rect -4852 -2160 -4812 2160
rect -492 -2160 -452 2160
rect -4852 -2200 -452 -2160
rect 160 2160 4560 2200
rect 160 -2160 200 2160
rect 4520 -2160 4560 2160
rect 160 -2200 4560 -2160
rect 5172 2160 9572 2200
rect 5172 -2160 5212 2160
rect 9532 -2160 9572 2160
rect 5172 -2200 9572 -2160
rect 10184 2160 14584 2200
rect 10184 -2160 10224 2160
rect 14544 -2160 14584 2160
rect 10184 -2200 14584 -2160
<< mimcapcontact >>
rect -14836 -2160 -10516 2160
rect -9824 -2160 -5504 2160
rect -4812 -2160 -492 2160
rect 200 -2160 4520 2160
rect 5212 -2160 9532 2160
rect 10224 -2160 14544 2160
<< metal4 >>
rect -10244 2212 -10148 2228
rect -14837 2160 -10515 2161
rect -14837 -2160 -14836 2160
rect -10516 -2160 -10515 2160
rect -14837 -2161 -10515 -2160
rect -10244 -2212 -10228 2212
rect -10164 -2212 -10148 2212
rect -5232 2212 -5136 2228
rect -9825 2160 -5503 2161
rect -9825 -2160 -9824 2160
rect -5504 -2160 -5503 2160
rect -9825 -2161 -5503 -2160
rect -10244 -2228 -10148 -2212
rect -5232 -2212 -5216 2212
rect -5152 -2212 -5136 2212
rect -220 2212 -124 2228
rect -4813 2160 -491 2161
rect -4813 -2160 -4812 2160
rect -492 -2160 -491 2160
rect -4813 -2161 -491 -2160
rect -5232 -2228 -5136 -2212
rect -220 -2212 -204 2212
rect -140 -2212 -124 2212
rect 4792 2212 4888 2228
rect 199 2160 4521 2161
rect 199 -2160 200 2160
rect 4520 -2160 4521 2160
rect 199 -2161 4521 -2160
rect -220 -2228 -124 -2212
rect 4792 -2212 4808 2212
rect 4872 -2212 4888 2212
rect 9804 2212 9900 2228
rect 5211 2160 9533 2161
rect 5211 -2160 5212 2160
rect 9532 -2160 9533 2160
rect 5211 -2161 9533 -2160
rect 4792 -2228 4888 -2212
rect 9804 -2212 9820 2212
rect 9884 -2212 9900 2212
rect 14816 2212 14912 2228
rect 10223 2160 14545 2161
rect 10223 -2160 10224 2160
rect 14544 -2160 14545 2160
rect 10223 -2161 14545 -2160
rect 9804 -2228 9900 -2212
rect 14816 -2212 14832 2212
rect 14896 -2212 14912 2212
rect 14816 -2228 14912 -2212
<< properties >>
string FIXED_BBOX 10144 -2240 14624 2240
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 22 l 22 val 984.72 carea 2.00 cperi 0.19 nx 6 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
