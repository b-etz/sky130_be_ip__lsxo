magic
tech sky130A
magscale 1 2
timestamp 1712088150
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 2060 0 1 -1966
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x2
timestamp 1707688321
transform 1 0 2128 0 1 -6994
box -38 -48 314 592
use level_shift  x3
timestamp 1712071977
transform 1 0 3450 0 1 -836
box 0 -2800 3195 480
use level_shift  x4
timestamp 1712071977
transform 1 0 3306 0 1 -5912
box 0 -2800 3195 480
use bias_gen  x5
timestamp 1712073863
transform 1 0 22450 0 1 -13914
box 0 -3410 15466 14020
use dout_amp  x6
timestamp 1712087189
transform 1 0 8616 0 1 -19538
box -1220 -12900 16982 200
use ripl_dly_clk_buf  x7
timestamp 1712087189
transform 1 0 39172 0 1 -19356
box 872 -3046 9184 598
use sky130_fd_pr__cap_mim_m3_1_KAF84V  XC1
timestamp 1712073300
transform 1 0 20978 0 1 -11888
box -886 -3440 886 3440
use sky130_fd_pr__cap_mim_m3_1_4RVTN9  XC2
timestamp 1712073300
transform 1 0 33690 0 1 -27026
box -5104 -9280 5104 9280
use sky130_fd_pr__cap_mim_m3_1_4HHTN9  XC3
timestamp 1712073300
transform 1 0 4652 0 1 -14256
box -1186 -4640 1186 4640
use sky130_fd_pr__cap_mim_m3_1_4HHTN9  XC4
timestamp 1712073300
transform 0 -1 44532 1 0 -23604
box -1186 -4640 1186 4640
use sky130_fd_pr__nfet_g5v0d10v5_GRGQJT  XM1
timestamp 1712087189
transform 1 0 17784 0 1 -9505
box -594 -1167 594 1167
use sky130_fd_pr__pfet_g5v0d10v5_47PSVV  XM2
timestamp 1712087189
transform 1 0 17988 0 1 -6949
box -1374 -1215 1374 1215
use sky130_fd_pr__nfet_01v8_AHZR5K  XM3
timestamp 1712071977
transform 1 0 26702 0 1 -22898
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_HZ6WG7  XM4
timestamp 1712071977
transform 1 0 48834 0 1 -21391
box -296 -285 296 285
use sky130_fd_pr__nfet_g5v0d10v5_ZPGQJT  XM5
timestamp 1712087189
transform 1 0 6508 0 1 -17572
box -594 -658 594 658
use sky130_fd_pr__pfet_g5v0d10v5_KLKQZ5  XM6
timestamp 1712087189
transform 1 0 6658 0 1 -10399
box -624 -697 624 697
use sky130_fd_pr__pfet_01v8_3H68VM  XM7
timestamp 1712071977
transform 1 0 48834 0 1 -20241
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_XPHWY6  XM8
timestamp 1712087189
transform 1 0 5810 0 1 -21175
box -562 -1137 562 1137
use sky130_fd_pr__pfet_g5v0d10v5_KL3SY6  XM9
timestamp 1712071977
transform 1 0 10998 0 1 -18743
box -308 -697 308 697
use sky130_fd_pr__nfet_01v8_Y5BWKS  XM11
timestamp 1712087189
transform 1 0 5690 0 1 -28839
box -562 -1119 562 1119
use sky130_fd_pr__res_xhigh_po_0p35_LKPHWV  XR2
timestamp 1712073300
transform 1 0 11706 0 1 -11556
box -4268 -5782 4268 5782
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 dvdd
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 dvss
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 ibias
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 ena
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 standby
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 dout
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 xin
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 xout
port 9 nsew
<< end >>
