magic
tech sky130A
magscale 1 2
timestamp 1712867472
<< error_s >>
rect 308 -917 7192 -596
rect 1735 -1047 1785 -1003
rect 386 -1131 439 -1047
rect 469 -1131 511 -1047
rect 541 -1131 633 -1047
rect 663 -1131 716 -1047
rect 833 -1131 885 -1047
rect 915 -1131 969 -1047
rect 999 -1131 1051 -1047
rect 1119 -1131 1224 -1047
rect 1254 -1059 1304 -1047
rect 1463 -1059 1581 -1047
rect 1254 -1131 1319 -1059
rect 1349 -1131 1415 -1059
rect 1445 -1131 1581 -1059
rect 1611 -1131 1653 -1047
rect 1683 -1131 1785 -1047
rect 1815 -1059 1869 -1003
rect 2039 -1059 2089 -1047
rect 1815 -1131 1884 -1059
rect 1914 -1131 1993 -1059
rect 2023 -1131 2089 -1059
rect 2119 -1131 2238 -1047
rect 2268 -1131 2329 -1047
rect 2359 -1131 2411 -1047
rect 2465 -1131 2517 -1001
rect 2547 -1131 2599 -1001
rect 2750 -1047 2802 -1001
rect 2653 -1131 2705 -1047
rect 2735 -1131 2802 -1047
rect 2832 -1131 2884 -1001
rect 3851 -1047 3901 -1003
rect 2949 -1131 3001 -1047
rect 3031 -1131 3085 -1047
rect 3115 -1131 3167 -1047
rect 3235 -1131 3340 -1047
rect 3370 -1059 3420 -1047
rect 3579 -1059 3697 -1047
rect 3370 -1131 3435 -1059
rect 3465 -1131 3531 -1059
rect 3561 -1131 3697 -1059
rect 3727 -1131 3769 -1047
rect 3799 -1131 3901 -1047
rect 3931 -1059 3985 -1003
rect 4155 -1059 4205 -1047
rect 3931 -1131 4000 -1059
rect 4030 -1131 4109 -1059
rect 4139 -1131 4205 -1059
rect 4235 -1131 4354 -1047
rect 4384 -1131 4445 -1047
rect 4475 -1131 4527 -1047
rect 4581 -1131 4633 -1001
rect 4663 -1131 4715 -1001
rect 4866 -1047 4918 -1001
rect 4769 -1131 4821 -1047
rect 4851 -1131 4918 -1047
rect 4948 -1131 5000 -1001
rect 5967 -1047 6017 -1003
rect 5065 -1131 5117 -1047
rect 5147 -1131 5201 -1047
rect 5231 -1131 5283 -1047
rect 5351 -1131 5456 -1047
rect 5486 -1059 5536 -1047
rect 5695 -1059 5813 -1047
rect 5486 -1131 5551 -1059
rect 5581 -1131 5647 -1059
rect 5677 -1131 5813 -1059
rect 5843 -1131 5885 -1047
rect 5915 -1131 6017 -1047
rect 6047 -1059 6101 -1003
rect 6271 -1059 6321 -1047
rect 6047 -1131 6116 -1059
rect 6146 -1131 6225 -1059
rect 6255 -1131 6321 -1059
rect 6351 -1131 6470 -1047
rect 6500 -1131 6561 -1047
rect 6591 -1131 6643 -1047
rect 6697 -1131 6749 -1001
rect 6779 -1131 6831 -1001
rect 6982 -1047 7034 -1001
rect 6885 -1131 6937 -1047
rect 6967 -1131 7034 -1047
rect 7064 -1131 7116 -1001
<< locali >>
rect 232 -792 432 -788
rect 232 -936 238 -792
rect 426 -936 432 -792
rect 7084 -816 7230 -806
rect 232 -940 432 -936
rect 736 -982 894 -854
rect 2852 -858 3010 -854
rect 2852 -972 2854 -858
rect 2986 -972 3010 -858
rect 4968 -860 5126 -854
rect 2852 -982 3010 -972
rect 4968 -974 4970 -860
rect 5102 -974 5126 -860
rect 7084 -930 7086 -816
rect 7218 -930 7230 -816
rect 7084 -940 7230 -930
rect 4968 -982 5126 -974
<< viali >>
rect 238 -936 426 -792
rect 536 -960 598 -856
rect 1102 -892 1142 -852
rect 2854 -972 2986 -858
rect 3218 -892 3258 -852
rect 4970 -974 5102 -860
rect 5336 -892 5376 -852
rect 7086 -930 7218 -816
<< metal1 >>
rect 232 -792 432 -748
rect 232 -936 238 -792
rect 426 -936 432 -792
rect 232 -948 432 -936
rect 522 -816 528 -716
rect 616 -816 622 -716
rect 522 -856 622 -816
rect 7074 -724 7230 -716
rect 7074 -846 7084 -724
rect 522 -960 536 -856
rect 598 -960 622 -856
rect 1090 -852 1256 -846
rect 1090 -892 1102 -852
rect 1142 -858 1256 -852
rect 1470 -858 1974 -846
rect 2092 -858 3000 -846
rect 1142 -886 2854 -858
rect 1142 -892 1256 -886
rect 1090 -898 1256 -892
rect 1380 -898 1974 -886
rect 2370 -898 2854 -886
rect 522 -976 622 -960
rect 2204 -928 2334 -920
rect 2204 -1044 2210 -928
rect 2326 -1044 2334 -928
rect 2842 -972 2854 -898
rect 2986 -898 3000 -858
rect 3206 -852 3372 -846
rect 3206 -892 3218 -852
rect 3258 -858 3372 -852
rect 3586 -858 4090 -846
rect 4208 -858 5114 -846
rect 3258 -860 5114 -858
rect 3258 -886 4970 -860
rect 3258 -892 3372 -886
rect 3206 -898 3372 -892
rect 3496 -898 4090 -886
rect 4486 -898 4970 -886
rect 2986 -972 2998 -898
rect 2842 -982 2998 -972
rect 4318 -926 4448 -920
rect 2204 -1050 2334 -1044
rect 4318 -1042 4326 -926
rect 4442 -1042 4448 -926
rect 4958 -974 4970 -898
rect 5102 -974 5114 -860
rect 5324 -852 5490 -846
rect 5324 -892 5336 -852
rect 5376 -858 5490 -852
rect 5700 -858 6204 -846
rect 6322 -858 7084 -846
rect 5376 -886 7084 -858
rect 5376 -892 5490 -886
rect 5324 -898 5490 -892
rect 5610 -898 6204 -886
rect 6602 -898 7084 -886
rect 4958 -980 5114 -974
rect 6434 -928 6564 -922
rect 4318 -1050 4448 -1042
rect 6434 -1044 6442 -928
rect 6558 -1044 6564 -928
rect 7074 -930 7084 -898
rect 7222 -930 7230 -724
rect 7074 -940 7230 -930
rect 6434 -1052 6564 -1044
<< via1 >>
rect 528 -816 616 -716
rect 7084 -816 7222 -724
rect 2210 -1044 2326 -928
rect 4326 -1042 4442 -926
rect 6442 -1044 6558 -928
rect 7084 -930 7086 -816
rect 7086 -930 7218 -816
rect 7218 -930 7222 -816
<< metal2 >>
rect 522 -816 528 -716
rect 616 -724 7230 -716
rect 616 -816 7084 -724
rect 2194 -926 2344 -910
rect 4308 -926 4458 -910
rect 6426 -926 6576 -912
rect 714 -928 4326 -926
rect 232 -1004 432 -976
rect 714 -1004 2210 -928
rect 232 -1044 2210 -1004
rect 2326 -1042 4326 -928
rect 4442 -928 6576 -926
rect 4442 -1042 6442 -928
rect 2326 -1044 6442 -1042
rect 6558 -1044 6576 -928
rect 7074 -930 7084 -816
rect 7222 -740 7230 -724
rect 7222 -930 7274 -740
rect 7074 -940 7274 -930
rect 232 -1046 6576 -1044
rect 232 -1136 832 -1046
rect 2194 -1060 2344 -1046
rect 4308 -1060 4458 -1046
rect 6426 -1062 6576 -1046
rect 232 -1176 432 -1136
use sky130_fd_sc_hd__and2_0  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712867472
transform 1 0 346 0 1 -1178
box -38 -48 498 592
use sky130_fd_sc_hd__dfrbp_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712867472
transform 1 0 806 0 1 -1178
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  x3
timestamp 1712867472
transform 1 0 2922 0 1 -1178
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  x4
timestamp 1712867472
transform 1 0 5038 0 1 -1178
box -38 -48 2154 592
<< labels >>
flabel space 346 -1226 7154 -1195 0 FreeSans 800 0 0 0 dvss
port 19 nsew
flabel space 3721 -682 3779 -586 0 FreeSans 800 0 0 0 dvdd
port 18 nsew
flabel metal2 7074 -940 7274 -740 0 FreeSans 800 0 0 0 doneb
port 14 nsew
flabel metal2 232 -1176 432 -976 0 FreeSans 800 0 0 0 ena
port 4 nsew
flabel space 6773 -1081 6839 -1047 0 FreeSans 800 0 0 0 done
port 5 nsew
flabel metal1 232 -948 432 -748 0 FreeSans 800 0 0 0 clkin
port 3 nsew
<< end >>
