magic
tech sky130A
magscale 1 2
timestamp 1713025933
<< nwell >>
rect -2398 -683 2398 683
<< pmos >>
rect -2202 64 -1802 464
rect -1630 64 -1230 464
rect -1058 64 -658 464
rect -486 64 -86 464
rect 86 64 486 464
rect 658 64 1058 464
rect 1230 64 1630 464
rect 1802 64 2202 464
rect -2202 -464 -1802 -64
rect -1630 -464 -1230 -64
rect -1058 -464 -658 -64
rect -486 -464 -86 -64
rect 86 -464 486 -64
rect 658 -464 1058 -64
rect 1230 -464 1630 -64
rect 1802 -464 2202 -64
<< pdiff >>
rect -2260 452 -2202 464
rect -2260 76 -2248 452
rect -2214 76 -2202 452
rect -2260 64 -2202 76
rect -1802 452 -1744 464
rect -1802 76 -1790 452
rect -1756 76 -1744 452
rect -1802 64 -1744 76
rect -1688 452 -1630 464
rect -1688 76 -1676 452
rect -1642 76 -1630 452
rect -1688 64 -1630 76
rect -1230 452 -1172 464
rect -1230 76 -1218 452
rect -1184 76 -1172 452
rect -1230 64 -1172 76
rect -1116 452 -1058 464
rect -1116 76 -1104 452
rect -1070 76 -1058 452
rect -1116 64 -1058 76
rect -658 452 -600 464
rect -658 76 -646 452
rect -612 76 -600 452
rect -658 64 -600 76
rect -544 452 -486 464
rect -544 76 -532 452
rect -498 76 -486 452
rect -544 64 -486 76
rect -86 452 -28 464
rect -86 76 -74 452
rect -40 76 -28 452
rect -86 64 -28 76
rect 28 452 86 464
rect 28 76 40 452
rect 74 76 86 452
rect 28 64 86 76
rect 486 452 544 464
rect 486 76 498 452
rect 532 76 544 452
rect 486 64 544 76
rect 600 452 658 464
rect 600 76 612 452
rect 646 76 658 452
rect 600 64 658 76
rect 1058 452 1116 464
rect 1058 76 1070 452
rect 1104 76 1116 452
rect 1058 64 1116 76
rect 1172 452 1230 464
rect 1172 76 1184 452
rect 1218 76 1230 452
rect 1172 64 1230 76
rect 1630 452 1688 464
rect 1630 76 1642 452
rect 1676 76 1688 452
rect 1630 64 1688 76
rect 1744 452 1802 464
rect 1744 76 1756 452
rect 1790 76 1802 452
rect 1744 64 1802 76
rect 2202 452 2260 464
rect 2202 76 2214 452
rect 2248 76 2260 452
rect 2202 64 2260 76
rect -2260 -76 -2202 -64
rect -2260 -452 -2248 -76
rect -2214 -452 -2202 -76
rect -2260 -464 -2202 -452
rect -1802 -76 -1744 -64
rect -1802 -452 -1790 -76
rect -1756 -452 -1744 -76
rect -1802 -464 -1744 -452
rect -1688 -76 -1630 -64
rect -1688 -452 -1676 -76
rect -1642 -452 -1630 -76
rect -1688 -464 -1630 -452
rect -1230 -76 -1172 -64
rect -1230 -452 -1218 -76
rect -1184 -452 -1172 -76
rect -1230 -464 -1172 -452
rect -1116 -76 -1058 -64
rect -1116 -452 -1104 -76
rect -1070 -452 -1058 -76
rect -1116 -464 -1058 -452
rect -658 -76 -600 -64
rect -658 -452 -646 -76
rect -612 -452 -600 -76
rect -658 -464 -600 -452
rect -544 -76 -486 -64
rect -544 -452 -532 -76
rect -498 -452 -486 -76
rect -544 -464 -486 -452
rect -86 -76 -28 -64
rect -86 -452 -74 -76
rect -40 -452 -28 -76
rect -86 -464 -28 -452
rect 28 -76 86 -64
rect 28 -452 40 -76
rect 74 -452 86 -76
rect 28 -464 86 -452
rect 486 -76 544 -64
rect 486 -452 498 -76
rect 532 -452 544 -76
rect 486 -464 544 -452
rect 600 -76 658 -64
rect 600 -452 612 -76
rect 646 -452 658 -76
rect 600 -464 658 -452
rect 1058 -76 1116 -64
rect 1058 -452 1070 -76
rect 1104 -452 1116 -76
rect 1058 -464 1116 -452
rect 1172 -76 1230 -64
rect 1172 -452 1184 -76
rect 1218 -452 1230 -76
rect 1172 -464 1230 -452
rect 1630 -76 1688 -64
rect 1630 -452 1642 -76
rect 1676 -452 1688 -76
rect 1630 -464 1688 -452
rect 1744 -76 1802 -64
rect 1744 -452 1756 -76
rect 1790 -452 1802 -76
rect 1744 -464 1802 -452
rect 2202 -76 2260 -64
rect 2202 -452 2214 -76
rect 2248 -452 2260 -76
rect 2202 -464 2260 -452
<< pdiffc >>
rect -2248 76 -2214 452
rect -1790 76 -1756 452
rect -1676 76 -1642 452
rect -1218 76 -1184 452
rect -1104 76 -1070 452
rect -646 76 -612 452
rect -532 76 -498 452
rect -74 76 -40 452
rect 40 76 74 452
rect 498 76 532 452
rect 612 76 646 452
rect 1070 76 1104 452
rect 1184 76 1218 452
rect 1642 76 1676 452
rect 1756 76 1790 452
rect 2214 76 2248 452
rect -2248 -452 -2214 -76
rect -1790 -452 -1756 -76
rect -1676 -452 -1642 -76
rect -1218 -452 -1184 -76
rect -1104 -452 -1070 -76
rect -646 -452 -612 -76
rect -532 -452 -498 -76
rect -74 -452 -40 -76
rect 40 -452 74 -76
rect 498 -452 532 -76
rect 612 -452 646 -76
rect 1070 -452 1104 -76
rect 1184 -452 1218 -76
rect 1642 -452 1676 -76
rect 1756 -452 1790 -76
rect 2214 -452 2248 -76
<< nsubdiff >>
rect -2362 613 -2266 647
rect 2266 613 2362 647
rect -2362 551 -2328 613
rect 2328 551 2362 613
rect -2362 -613 -2328 -551
rect 2328 -613 2362 -551
rect -2362 -647 -2266 -613
rect 2266 -647 2362 -613
<< nsubdiffcont >>
rect -2266 613 2266 647
rect -2362 -551 -2328 551
rect 2328 -551 2362 551
rect -2266 -647 2266 -613
<< poly >>
rect -2202 545 -1802 561
rect -2202 511 -2186 545
rect -1818 511 -1802 545
rect -2202 464 -1802 511
rect -1630 545 -1230 561
rect -1630 511 -1614 545
rect -1246 511 -1230 545
rect -1630 464 -1230 511
rect -1058 545 -658 561
rect -1058 511 -1042 545
rect -674 511 -658 545
rect -1058 464 -658 511
rect -486 545 -86 561
rect -486 511 -470 545
rect -102 511 -86 545
rect -486 464 -86 511
rect 86 545 486 561
rect 86 511 102 545
rect 470 511 486 545
rect 86 464 486 511
rect 658 545 1058 561
rect 658 511 674 545
rect 1042 511 1058 545
rect 658 464 1058 511
rect 1230 545 1630 561
rect 1230 511 1246 545
rect 1614 511 1630 545
rect 1230 464 1630 511
rect 1802 545 2202 561
rect 1802 511 1818 545
rect 2186 511 2202 545
rect 1802 464 2202 511
rect -2202 17 -1802 64
rect -2202 -17 -2186 17
rect -1818 -17 -1802 17
rect -2202 -64 -1802 -17
rect -1630 17 -1230 64
rect -1630 -17 -1614 17
rect -1246 -17 -1230 17
rect -1630 -64 -1230 -17
rect -1058 17 -658 64
rect -1058 -17 -1042 17
rect -674 -17 -658 17
rect -1058 -64 -658 -17
rect -486 17 -86 64
rect -486 -17 -470 17
rect -102 -17 -86 17
rect -486 -64 -86 -17
rect 86 17 486 64
rect 86 -17 102 17
rect 470 -17 486 17
rect 86 -64 486 -17
rect 658 17 1058 64
rect 658 -17 674 17
rect 1042 -17 1058 17
rect 658 -64 1058 -17
rect 1230 17 1630 64
rect 1230 -17 1246 17
rect 1614 -17 1630 17
rect 1230 -64 1630 -17
rect 1802 17 2202 64
rect 1802 -17 1818 17
rect 2186 -17 2202 17
rect 1802 -64 2202 -17
rect -2202 -511 -1802 -464
rect -2202 -545 -2186 -511
rect -1818 -545 -1802 -511
rect -2202 -561 -1802 -545
rect -1630 -511 -1230 -464
rect -1630 -545 -1614 -511
rect -1246 -545 -1230 -511
rect -1630 -561 -1230 -545
rect -1058 -511 -658 -464
rect -1058 -545 -1042 -511
rect -674 -545 -658 -511
rect -1058 -561 -658 -545
rect -486 -511 -86 -464
rect -486 -545 -470 -511
rect -102 -545 -86 -511
rect -486 -561 -86 -545
rect 86 -511 486 -464
rect 86 -545 102 -511
rect 470 -545 486 -511
rect 86 -561 486 -545
rect 658 -511 1058 -464
rect 658 -545 674 -511
rect 1042 -545 1058 -511
rect 658 -561 1058 -545
rect 1230 -511 1630 -464
rect 1230 -545 1246 -511
rect 1614 -545 1630 -511
rect 1230 -561 1630 -545
rect 1802 -511 2202 -464
rect 1802 -545 1818 -511
rect 2186 -545 2202 -511
rect 1802 -561 2202 -545
<< polycont >>
rect -2186 511 -1818 545
rect -1614 511 -1246 545
rect -1042 511 -674 545
rect -470 511 -102 545
rect 102 511 470 545
rect 674 511 1042 545
rect 1246 511 1614 545
rect 1818 511 2186 545
rect -2186 -17 -1818 17
rect -1614 -17 -1246 17
rect -1042 -17 -674 17
rect -470 -17 -102 17
rect 102 -17 470 17
rect 674 -17 1042 17
rect 1246 -17 1614 17
rect 1818 -17 2186 17
rect -2186 -545 -1818 -511
rect -1614 -545 -1246 -511
rect -1042 -545 -674 -511
rect -470 -545 -102 -511
rect 102 -545 470 -511
rect 674 -545 1042 -511
rect 1246 -545 1614 -511
rect 1818 -545 2186 -511
<< locali >>
rect -2362 613 -2266 647
rect 2266 613 2362 647
rect -2362 551 -2328 613
rect 2328 551 2362 613
rect -2202 511 -2186 545
rect -1818 511 -1802 545
rect -1630 511 -1614 545
rect -1246 511 -1230 545
rect -1058 511 -1042 545
rect -674 511 -658 545
rect -486 511 -470 545
rect -102 511 -86 545
rect 86 511 102 545
rect 470 511 486 545
rect 658 511 674 545
rect 1042 511 1058 545
rect 1230 511 1246 545
rect 1614 511 1630 545
rect 1802 511 1818 545
rect 2186 511 2202 545
rect -2248 452 -2214 468
rect -2248 60 -2214 76
rect -1790 452 -1756 468
rect -1790 60 -1756 76
rect -1676 452 -1642 468
rect -1676 60 -1642 76
rect -1218 452 -1184 468
rect -1218 60 -1184 76
rect -1104 452 -1070 468
rect -1104 60 -1070 76
rect -646 452 -612 468
rect -646 60 -612 76
rect -532 452 -498 468
rect -532 60 -498 76
rect -74 452 -40 468
rect -74 60 -40 76
rect 40 452 74 468
rect 40 60 74 76
rect 498 452 532 468
rect 498 60 532 76
rect 612 452 646 468
rect 612 60 646 76
rect 1070 452 1104 468
rect 1070 60 1104 76
rect 1184 452 1218 468
rect 1184 60 1218 76
rect 1642 452 1676 468
rect 1642 60 1676 76
rect 1756 452 1790 468
rect 1756 60 1790 76
rect 2214 452 2248 468
rect 2214 60 2248 76
rect -2202 -17 -2186 17
rect -1818 -17 -1802 17
rect -1630 -17 -1614 17
rect -1246 -17 -1230 17
rect -1058 -17 -1042 17
rect -674 -17 -658 17
rect -486 -17 -470 17
rect -102 -17 -86 17
rect 86 -17 102 17
rect 470 -17 486 17
rect 658 -17 674 17
rect 1042 -17 1058 17
rect 1230 -17 1246 17
rect 1614 -17 1630 17
rect 1802 -17 1818 17
rect 2186 -17 2202 17
rect -2248 -76 -2214 -60
rect -2248 -468 -2214 -452
rect -1790 -76 -1756 -60
rect -1790 -468 -1756 -452
rect -1676 -76 -1642 -60
rect -1676 -468 -1642 -452
rect -1218 -76 -1184 -60
rect -1218 -468 -1184 -452
rect -1104 -76 -1070 -60
rect -1104 -468 -1070 -452
rect -646 -76 -612 -60
rect -646 -468 -612 -452
rect -532 -76 -498 -60
rect -532 -468 -498 -452
rect -74 -76 -40 -60
rect -74 -468 -40 -452
rect 40 -76 74 -60
rect 40 -468 74 -452
rect 498 -76 532 -60
rect 498 -468 532 -452
rect 612 -76 646 -60
rect 612 -468 646 -452
rect 1070 -76 1104 -60
rect 1070 -468 1104 -452
rect 1184 -76 1218 -60
rect 1184 -468 1218 -452
rect 1642 -76 1676 -60
rect 1642 -468 1676 -452
rect 1756 -76 1790 -60
rect 1756 -468 1790 -452
rect 2214 -76 2248 -60
rect 2214 -468 2248 -452
rect -2202 -545 -2186 -511
rect -1818 -545 -1802 -511
rect -1630 -545 -1614 -511
rect -1246 -545 -1230 -511
rect -1058 -545 -1042 -511
rect -674 -545 -658 -511
rect -486 -545 -470 -511
rect -102 -545 -86 -511
rect 86 -545 102 -511
rect 470 -545 486 -511
rect 658 -545 674 -511
rect 1042 -545 1058 -511
rect 1230 -545 1246 -511
rect 1614 -545 1630 -511
rect 1802 -545 1818 -511
rect 2186 -545 2202 -511
rect -2362 -613 -2328 -551
rect 2328 -613 2362 -551
rect -2362 -647 -2266 -613
rect 2266 -647 2362 -613
<< viali >>
rect -2149 511 -1855 545
rect -1577 511 -1283 545
rect -1005 511 -711 545
rect -433 511 -139 545
rect 139 511 433 545
rect 711 511 1005 545
rect 1283 511 1577 545
rect 1855 511 2149 545
rect -2248 76 -2214 452
rect -1790 76 -1756 452
rect -1676 76 -1642 452
rect -1218 76 -1184 452
rect -1104 76 -1070 452
rect -646 76 -612 452
rect -532 76 -498 452
rect -74 76 -40 452
rect 40 76 74 452
rect 498 76 532 452
rect 612 76 646 452
rect 1070 76 1104 452
rect 1184 76 1218 452
rect 1642 76 1676 452
rect 1756 76 1790 452
rect 2214 76 2248 452
rect -2149 -17 -1855 17
rect -1577 -17 -1283 17
rect -1005 -17 -711 17
rect -433 -17 -139 17
rect 139 -17 433 17
rect 711 -17 1005 17
rect 1283 -17 1577 17
rect 1855 -17 2149 17
rect -2248 -452 -2214 -76
rect -1790 -452 -1756 -76
rect -1676 -452 -1642 -76
rect -1218 -452 -1184 -76
rect -1104 -452 -1070 -76
rect -646 -452 -612 -76
rect -532 -452 -498 -76
rect -74 -452 -40 -76
rect 40 -452 74 -76
rect 498 -452 532 -76
rect 612 -452 646 -76
rect 1070 -452 1104 -76
rect 1184 -452 1218 -76
rect 1642 -452 1676 -76
rect 1756 -452 1790 -76
rect 2214 -452 2248 -76
rect -2149 -545 -1855 -511
rect -1577 -545 -1283 -511
rect -1005 -545 -711 -511
rect -433 -545 -139 -511
rect 139 -545 433 -511
rect 711 -545 1005 -511
rect 1283 -545 1577 -511
rect 1855 -545 2149 -511
<< metal1 >>
rect -2161 545 -1843 551
rect -2161 511 -2149 545
rect -1855 511 -1843 545
rect -2161 505 -1843 511
rect -1589 545 -1271 551
rect -1589 511 -1577 545
rect -1283 511 -1271 545
rect -1589 505 -1271 511
rect -1017 545 -699 551
rect -1017 511 -1005 545
rect -711 511 -699 545
rect -1017 505 -699 511
rect -445 545 -127 551
rect -445 511 -433 545
rect -139 511 -127 545
rect -445 505 -127 511
rect 127 545 445 551
rect 127 511 139 545
rect 433 511 445 545
rect 127 505 445 511
rect 699 545 1017 551
rect 699 511 711 545
rect 1005 511 1017 545
rect 699 505 1017 511
rect 1271 545 1589 551
rect 1271 511 1283 545
rect 1577 511 1589 545
rect 1271 505 1589 511
rect 1843 545 2161 551
rect 1843 511 1855 545
rect 2149 511 2161 545
rect 1843 505 2161 511
rect -2254 452 -2208 464
rect -2254 76 -2248 452
rect -2214 76 -2208 452
rect -2254 64 -2208 76
rect -1796 452 -1750 464
rect -1796 76 -1790 452
rect -1756 76 -1750 452
rect -1796 64 -1750 76
rect -1682 452 -1636 464
rect -1682 76 -1676 452
rect -1642 76 -1636 452
rect -1682 64 -1636 76
rect -1224 452 -1178 464
rect -1224 76 -1218 452
rect -1184 76 -1178 452
rect -1224 64 -1178 76
rect -1110 452 -1064 464
rect -1110 76 -1104 452
rect -1070 76 -1064 452
rect -1110 64 -1064 76
rect -652 452 -606 464
rect -652 76 -646 452
rect -612 76 -606 452
rect -652 64 -606 76
rect -538 452 -492 464
rect -538 76 -532 452
rect -498 76 -492 452
rect -538 64 -492 76
rect -80 452 -34 464
rect -80 76 -74 452
rect -40 76 -34 452
rect -80 64 -34 76
rect 34 452 80 464
rect 34 76 40 452
rect 74 76 80 452
rect 34 64 80 76
rect 492 452 538 464
rect 492 76 498 452
rect 532 76 538 452
rect 492 64 538 76
rect 606 452 652 464
rect 606 76 612 452
rect 646 76 652 452
rect 606 64 652 76
rect 1064 452 1110 464
rect 1064 76 1070 452
rect 1104 76 1110 452
rect 1064 64 1110 76
rect 1178 452 1224 464
rect 1178 76 1184 452
rect 1218 76 1224 452
rect 1178 64 1224 76
rect 1636 452 1682 464
rect 1636 76 1642 452
rect 1676 76 1682 452
rect 1636 64 1682 76
rect 1750 452 1796 464
rect 1750 76 1756 452
rect 1790 76 1796 452
rect 1750 64 1796 76
rect 2208 452 2254 464
rect 2208 76 2214 452
rect 2248 76 2254 452
rect 2208 64 2254 76
rect -2161 17 -1843 23
rect -2161 -17 -2149 17
rect -1855 -17 -1843 17
rect -2161 -23 -1843 -17
rect -1589 17 -1271 23
rect -1589 -17 -1577 17
rect -1283 -17 -1271 17
rect -1589 -23 -1271 -17
rect -1017 17 -699 23
rect -1017 -17 -1005 17
rect -711 -17 -699 17
rect -1017 -23 -699 -17
rect -445 17 -127 23
rect -445 -17 -433 17
rect -139 -17 -127 17
rect -445 -23 -127 -17
rect 127 17 445 23
rect 127 -17 139 17
rect 433 -17 445 17
rect 127 -23 445 -17
rect 699 17 1017 23
rect 699 -17 711 17
rect 1005 -17 1017 17
rect 699 -23 1017 -17
rect 1271 17 1589 23
rect 1271 -17 1283 17
rect 1577 -17 1589 17
rect 1271 -23 1589 -17
rect 1843 17 2161 23
rect 1843 -17 1855 17
rect 2149 -17 2161 17
rect 1843 -23 2161 -17
rect -2254 -76 -2208 -64
rect -2254 -452 -2248 -76
rect -2214 -452 -2208 -76
rect -2254 -464 -2208 -452
rect -1796 -76 -1750 -64
rect -1796 -452 -1790 -76
rect -1756 -452 -1750 -76
rect -1796 -464 -1750 -452
rect -1682 -76 -1636 -64
rect -1682 -452 -1676 -76
rect -1642 -452 -1636 -76
rect -1682 -464 -1636 -452
rect -1224 -76 -1178 -64
rect -1224 -452 -1218 -76
rect -1184 -452 -1178 -76
rect -1224 -464 -1178 -452
rect -1110 -76 -1064 -64
rect -1110 -452 -1104 -76
rect -1070 -452 -1064 -76
rect -1110 -464 -1064 -452
rect -652 -76 -606 -64
rect -652 -452 -646 -76
rect -612 -452 -606 -76
rect -652 -464 -606 -452
rect -538 -76 -492 -64
rect -538 -452 -532 -76
rect -498 -452 -492 -76
rect -538 -464 -492 -452
rect -80 -76 -34 -64
rect -80 -452 -74 -76
rect -40 -452 -34 -76
rect -80 -464 -34 -452
rect 34 -76 80 -64
rect 34 -452 40 -76
rect 74 -452 80 -76
rect 34 -464 80 -452
rect 492 -76 538 -64
rect 492 -452 498 -76
rect 532 -452 538 -76
rect 492 -464 538 -452
rect 606 -76 652 -64
rect 606 -452 612 -76
rect 646 -452 652 -76
rect 606 -464 652 -452
rect 1064 -76 1110 -64
rect 1064 -452 1070 -76
rect 1104 -452 1110 -76
rect 1064 -464 1110 -452
rect 1178 -76 1224 -64
rect 1178 -452 1184 -76
rect 1218 -452 1224 -76
rect 1178 -464 1224 -452
rect 1636 -76 1682 -64
rect 1636 -452 1642 -76
rect 1676 -452 1682 -76
rect 1636 -464 1682 -452
rect 1750 -76 1796 -64
rect 1750 -452 1756 -76
rect 1790 -452 1796 -76
rect 1750 -464 1796 -452
rect 2208 -76 2254 -64
rect 2208 -452 2214 -76
rect 2248 -452 2254 -76
rect 2208 -464 2254 -452
rect -2161 -511 -1843 -505
rect -2161 -545 -2149 -511
rect -1855 -545 -1843 -511
rect -2161 -551 -1843 -545
rect -1589 -511 -1271 -505
rect -1589 -545 -1577 -511
rect -1283 -545 -1271 -511
rect -1589 -551 -1271 -545
rect -1017 -511 -699 -505
rect -1017 -545 -1005 -511
rect -711 -545 -699 -511
rect -1017 -551 -699 -545
rect -445 -511 -127 -505
rect -445 -545 -433 -511
rect -139 -545 -127 -511
rect -445 -551 -127 -545
rect 127 -511 445 -505
rect 127 -545 139 -511
rect 433 -545 445 -511
rect 127 -551 445 -545
rect 699 -511 1017 -505
rect 699 -545 711 -511
rect 1005 -545 1017 -511
rect 699 -551 1017 -545
rect 1271 -511 1589 -505
rect 1271 -545 1283 -511
rect 1577 -545 1589 -511
rect 1271 -551 1589 -545
rect 1843 -511 2161 -505
rect 1843 -545 1855 -511
rect 2149 -545 2161 -511
rect 1843 -551 2161 -545
<< properties >>
string FIXED_BBOX -2345 -630 2345 630
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 2 m 2 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
