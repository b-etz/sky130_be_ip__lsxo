magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< pwell >>
rect -201 -260582 201 260582
<< psubdiff >>
rect -165 260512 -69 260546
rect 69 260512 165 260546
rect -165 260450 -131 260512
rect 131 260450 165 260512
rect -165 -260512 -131 -260450
rect 131 -260512 165 -260450
rect -165 -260546 -69 -260512
rect 69 -260546 165 -260512
<< psubdiffcont >>
rect -69 260512 69 260546
rect -165 -260450 -131 260450
rect 131 -260450 165 260450
rect -69 -260546 69 -260512
<< xpolycontact >>
rect -35 259984 35 260416
rect -35 -260416 35 -259984
<< xpolyres >>
rect -35 -259984 35 259984
<< locali >>
rect -165 260512 -69 260546
rect 69 260512 165 260546
rect -165 260450 -131 260512
rect 131 260450 165 260512
rect -165 -260512 -131 -260450
rect 131 -260512 165 -260450
rect -165 -260546 -69 -260512
rect 69 -260546 165 -260512
<< viali >>
rect -19 260001 19 260398
rect -19 -260398 19 -260001
<< metal1 >>
rect -25 260398 25 260410
rect -25 260001 -19 260398
rect 19 260001 25 260398
rect -25 259989 25 260001
rect -25 -260001 25 -259989
rect -25 -260398 -19 -260001
rect 19 -260398 25 -260001
rect -25 -260410 25 -260398
<< properties >>
string FIXED_BBOX -148 -260529 148 260529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 2600.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 14.858meg dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
