magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< pwell >>
rect -2193 -4582 2193 4582
<< psubdiff >>
rect -2157 4512 -2061 4546
rect 2061 4512 2157 4546
rect -2157 4450 -2123 4512
rect 2123 4450 2157 4512
rect -2157 -4512 -2123 -4450
rect 2123 -4512 2157 -4450
rect -2157 -4546 -2061 -4512
rect 2061 -4546 2157 -4512
<< psubdiffcont >>
rect -2061 4512 2061 4546
rect -2157 -4450 -2123 4450
rect 2123 -4450 2157 4450
rect -2061 -4546 2061 -4512
<< xpolycontact >>
rect -2027 3984 -1957 4416
rect -2027 -4416 -1957 -3984
rect -1861 3984 -1791 4416
rect -1861 -4416 -1791 -3984
rect -1695 3984 -1625 4416
rect -1695 -4416 -1625 -3984
rect -1529 3984 -1459 4416
rect -1529 -4416 -1459 -3984
rect -1363 3984 -1293 4416
rect -1363 -4416 -1293 -3984
rect -1197 3984 -1127 4416
rect -1197 -4416 -1127 -3984
rect -1031 3984 -961 4416
rect -1031 -4416 -961 -3984
rect -865 3984 -795 4416
rect -865 -4416 -795 -3984
rect -699 3984 -629 4416
rect -699 -4416 -629 -3984
rect -533 3984 -463 4416
rect -533 -4416 -463 -3984
rect -367 3984 -297 4416
rect -367 -4416 -297 -3984
rect -201 3984 -131 4416
rect -201 -4416 -131 -3984
rect -35 3984 35 4416
rect -35 -4416 35 -3984
rect 131 3984 201 4416
rect 131 -4416 201 -3984
rect 297 3984 367 4416
rect 297 -4416 367 -3984
rect 463 3984 533 4416
rect 463 -4416 533 -3984
rect 629 3984 699 4416
rect 629 -4416 699 -3984
rect 795 3984 865 4416
rect 795 -4416 865 -3984
rect 961 3984 1031 4416
rect 961 -4416 1031 -3984
rect 1127 3984 1197 4416
rect 1127 -4416 1197 -3984
rect 1293 3984 1363 4416
rect 1293 -4416 1363 -3984
rect 1459 3984 1529 4416
rect 1459 -4416 1529 -3984
rect 1625 3984 1695 4416
rect 1625 -4416 1695 -3984
rect 1791 3984 1861 4416
rect 1791 -4416 1861 -3984
rect 1957 3984 2027 4416
rect 1957 -4416 2027 -3984
<< xpolyres >>
rect -2027 -3984 -1957 3984
rect -1861 -3984 -1791 3984
rect -1695 -3984 -1625 3984
rect -1529 -3984 -1459 3984
rect -1363 -3984 -1293 3984
rect -1197 -3984 -1127 3984
rect -1031 -3984 -961 3984
rect -865 -3984 -795 3984
rect -699 -3984 -629 3984
rect -533 -3984 -463 3984
rect -367 -3984 -297 3984
rect -201 -3984 -131 3984
rect -35 -3984 35 3984
rect 131 -3984 201 3984
rect 297 -3984 367 3984
rect 463 -3984 533 3984
rect 629 -3984 699 3984
rect 795 -3984 865 3984
rect 961 -3984 1031 3984
rect 1127 -3984 1197 3984
rect 1293 -3984 1363 3984
rect 1459 -3984 1529 3984
rect 1625 -3984 1695 3984
rect 1791 -3984 1861 3984
rect 1957 -3984 2027 3984
<< locali >>
rect -2157 4512 -2061 4546
rect 2061 4512 2157 4546
rect -2157 4450 -2123 4512
rect 2123 4450 2157 4512
rect -2157 -4512 -2123 -4450
rect 2123 -4512 2157 -4450
rect -2157 -4546 -2061 -4512
rect 2061 -4546 2157 -4512
<< viali >>
rect -2011 4001 -1973 4398
rect -1845 4001 -1807 4398
rect -1679 4001 -1641 4398
rect -1513 4001 -1475 4398
rect -1347 4001 -1309 4398
rect -1181 4001 -1143 4398
rect -1015 4001 -977 4398
rect -849 4001 -811 4398
rect -683 4001 -645 4398
rect -517 4001 -479 4398
rect -351 4001 -313 4398
rect -185 4001 -147 4398
rect -19 4001 19 4398
rect 147 4001 185 4398
rect 313 4001 351 4398
rect 479 4001 517 4398
rect 645 4001 683 4398
rect 811 4001 849 4398
rect 977 4001 1015 4398
rect 1143 4001 1181 4398
rect 1309 4001 1347 4398
rect 1475 4001 1513 4398
rect 1641 4001 1679 4398
rect 1807 4001 1845 4398
rect 1973 4001 2011 4398
rect -2011 -4398 -1973 -4001
rect -1845 -4398 -1807 -4001
rect -1679 -4398 -1641 -4001
rect -1513 -4398 -1475 -4001
rect -1347 -4398 -1309 -4001
rect -1181 -4398 -1143 -4001
rect -1015 -4398 -977 -4001
rect -849 -4398 -811 -4001
rect -683 -4398 -645 -4001
rect -517 -4398 -479 -4001
rect -351 -4398 -313 -4001
rect -185 -4398 -147 -4001
rect -19 -4398 19 -4001
rect 147 -4398 185 -4001
rect 313 -4398 351 -4001
rect 479 -4398 517 -4001
rect 645 -4398 683 -4001
rect 811 -4398 849 -4001
rect 977 -4398 1015 -4001
rect 1143 -4398 1181 -4001
rect 1309 -4398 1347 -4001
rect 1475 -4398 1513 -4001
rect 1641 -4398 1679 -4001
rect 1807 -4398 1845 -4001
rect 1973 -4398 2011 -4001
<< metal1 >>
rect -2017 4398 -1967 4410
rect -2017 4001 -2011 4398
rect -1973 4001 -1967 4398
rect -2017 3989 -1967 4001
rect -1851 4398 -1801 4410
rect -1851 4001 -1845 4398
rect -1807 4001 -1801 4398
rect -1851 3989 -1801 4001
rect -1685 4398 -1635 4410
rect -1685 4001 -1679 4398
rect -1641 4001 -1635 4398
rect -1685 3989 -1635 4001
rect -1519 4398 -1469 4410
rect -1519 4001 -1513 4398
rect -1475 4001 -1469 4398
rect -1519 3989 -1469 4001
rect -1353 4398 -1303 4410
rect -1353 4001 -1347 4398
rect -1309 4001 -1303 4398
rect -1353 3989 -1303 4001
rect -1187 4398 -1137 4410
rect -1187 4001 -1181 4398
rect -1143 4001 -1137 4398
rect -1187 3989 -1137 4001
rect -1021 4398 -971 4410
rect -1021 4001 -1015 4398
rect -977 4001 -971 4398
rect -1021 3989 -971 4001
rect -855 4398 -805 4410
rect -855 4001 -849 4398
rect -811 4001 -805 4398
rect -855 3989 -805 4001
rect -689 4398 -639 4410
rect -689 4001 -683 4398
rect -645 4001 -639 4398
rect -689 3989 -639 4001
rect -523 4398 -473 4410
rect -523 4001 -517 4398
rect -479 4001 -473 4398
rect -523 3989 -473 4001
rect -357 4398 -307 4410
rect -357 4001 -351 4398
rect -313 4001 -307 4398
rect -357 3989 -307 4001
rect -191 4398 -141 4410
rect -191 4001 -185 4398
rect -147 4001 -141 4398
rect -191 3989 -141 4001
rect -25 4398 25 4410
rect -25 4001 -19 4398
rect 19 4001 25 4398
rect -25 3989 25 4001
rect 141 4398 191 4410
rect 141 4001 147 4398
rect 185 4001 191 4398
rect 141 3989 191 4001
rect 307 4398 357 4410
rect 307 4001 313 4398
rect 351 4001 357 4398
rect 307 3989 357 4001
rect 473 4398 523 4410
rect 473 4001 479 4398
rect 517 4001 523 4398
rect 473 3989 523 4001
rect 639 4398 689 4410
rect 639 4001 645 4398
rect 683 4001 689 4398
rect 639 3989 689 4001
rect 805 4398 855 4410
rect 805 4001 811 4398
rect 849 4001 855 4398
rect 805 3989 855 4001
rect 971 4398 1021 4410
rect 971 4001 977 4398
rect 1015 4001 1021 4398
rect 971 3989 1021 4001
rect 1137 4398 1187 4410
rect 1137 4001 1143 4398
rect 1181 4001 1187 4398
rect 1137 3989 1187 4001
rect 1303 4398 1353 4410
rect 1303 4001 1309 4398
rect 1347 4001 1353 4398
rect 1303 3989 1353 4001
rect 1469 4398 1519 4410
rect 1469 4001 1475 4398
rect 1513 4001 1519 4398
rect 1469 3989 1519 4001
rect 1635 4398 1685 4410
rect 1635 4001 1641 4398
rect 1679 4001 1685 4398
rect 1635 3989 1685 4001
rect 1801 4398 1851 4410
rect 1801 4001 1807 4398
rect 1845 4001 1851 4398
rect 1801 3989 1851 4001
rect 1967 4398 2017 4410
rect 1967 4001 1973 4398
rect 2011 4001 2017 4398
rect 1967 3989 2017 4001
rect -2017 -4001 -1967 -3989
rect -2017 -4398 -2011 -4001
rect -1973 -4398 -1967 -4001
rect -2017 -4410 -1967 -4398
rect -1851 -4001 -1801 -3989
rect -1851 -4398 -1845 -4001
rect -1807 -4398 -1801 -4001
rect -1851 -4410 -1801 -4398
rect -1685 -4001 -1635 -3989
rect -1685 -4398 -1679 -4001
rect -1641 -4398 -1635 -4001
rect -1685 -4410 -1635 -4398
rect -1519 -4001 -1469 -3989
rect -1519 -4398 -1513 -4001
rect -1475 -4398 -1469 -4001
rect -1519 -4410 -1469 -4398
rect -1353 -4001 -1303 -3989
rect -1353 -4398 -1347 -4001
rect -1309 -4398 -1303 -4001
rect -1353 -4410 -1303 -4398
rect -1187 -4001 -1137 -3989
rect -1187 -4398 -1181 -4001
rect -1143 -4398 -1137 -4001
rect -1187 -4410 -1137 -4398
rect -1021 -4001 -971 -3989
rect -1021 -4398 -1015 -4001
rect -977 -4398 -971 -4001
rect -1021 -4410 -971 -4398
rect -855 -4001 -805 -3989
rect -855 -4398 -849 -4001
rect -811 -4398 -805 -4001
rect -855 -4410 -805 -4398
rect -689 -4001 -639 -3989
rect -689 -4398 -683 -4001
rect -645 -4398 -639 -4001
rect -689 -4410 -639 -4398
rect -523 -4001 -473 -3989
rect -523 -4398 -517 -4001
rect -479 -4398 -473 -4001
rect -523 -4410 -473 -4398
rect -357 -4001 -307 -3989
rect -357 -4398 -351 -4001
rect -313 -4398 -307 -4001
rect -357 -4410 -307 -4398
rect -191 -4001 -141 -3989
rect -191 -4398 -185 -4001
rect -147 -4398 -141 -4001
rect -191 -4410 -141 -4398
rect -25 -4001 25 -3989
rect -25 -4398 -19 -4001
rect 19 -4398 25 -4001
rect -25 -4410 25 -4398
rect 141 -4001 191 -3989
rect 141 -4398 147 -4001
rect 185 -4398 191 -4001
rect 141 -4410 191 -4398
rect 307 -4001 357 -3989
rect 307 -4398 313 -4001
rect 351 -4398 357 -4001
rect 307 -4410 357 -4398
rect 473 -4001 523 -3989
rect 473 -4398 479 -4001
rect 517 -4398 523 -4001
rect 473 -4410 523 -4398
rect 639 -4001 689 -3989
rect 639 -4398 645 -4001
rect 683 -4398 689 -4001
rect 639 -4410 689 -4398
rect 805 -4001 855 -3989
rect 805 -4398 811 -4001
rect 849 -4398 855 -4001
rect 805 -4410 855 -4398
rect 971 -4001 1021 -3989
rect 971 -4398 977 -4001
rect 1015 -4398 1021 -4001
rect 971 -4410 1021 -4398
rect 1137 -4001 1187 -3989
rect 1137 -4398 1143 -4001
rect 1181 -4398 1187 -4001
rect 1137 -4410 1187 -4398
rect 1303 -4001 1353 -3989
rect 1303 -4398 1309 -4001
rect 1347 -4398 1353 -4001
rect 1303 -4410 1353 -4398
rect 1469 -4001 1519 -3989
rect 1469 -4398 1475 -4001
rect 1513 -4398 1519 -4001
rect 1469 -4410 1519 -4398
rect 1635 -4001 1685 -3989
rect 1635 -4398 1641 -4001
rect 1679 -4398 1685 -4001
rect 1635 -4410 1685 -4398
rect 1801 -4001 1851 -3989
rect 1801 -4398 1807 -4001
rect 1845 -4398 1851 -4001
rect 1801 -4410 1851 -4398
rect 1967 -4001 2017 -3989
rect 1967 -4398 1973 -4001
rect 2011 -4398 2017 -4001
rect 1967 -4410 2017 -4398
<< properties >>
string FIXED_BBOX -2140 -4529 2140 4529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 40.0 m 1 nx 25 wmin 0.350 lmin 0.50 rho 2000 val 229.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
