magic
tech sky130A
magscale 1 2
timestamp 1713210209
<< pwell >>
rect -1083 -610 1083 610
<< nmos >>
rect -887 -400 -487 400
rect -429 -400 -29 400
rect 29 -400 429 400
rect 487 -400 887 400
<< ndiff >>
rect -945 388 -887 400
rect -945 -388 -933 388
rect -899 -388 -887 388
rect -945 -400 -887 -388
rect -487 388 -429 400
rect -487 -388 -475 388
rect -441 -388 -429 388
rect -487 -400 -429 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 429 388 487 400
rect 429 -388 441 388
rect 475 -388 487 388
rect 429 -400 487 -388
rect 887 388 945 400
rect 887 -388 899 388
rect 933 -388 945 388
rect 887 -400 945 -388
<< ndiffc >>
rect -933 -388 -899 388
rect -475 -388 -441 388
rect -17 -388 17 388
rect 441 -388 475 388
rect 899 -388 933 388
<< psubdiff >>
rect -1047 540 -951 574
rect 951 540 1047 574
rect -1047 478 -1013 540
rect 1013 478 1047 540
rect -1047 -540 -1013 -478
rect 1013 -540 1047 -478
rect -1047 -574 -951 -540
rect 951 -574 1047 -540
<< psubdiffcont >>
rect -951 540 951 574
rect -1047 -478 -1013 478
rect 1013 -478 1047 478
rect -951 -574 951 -540
<< poly >>
rect -887 472 -487 488
rect -887 438 -871 472
rect -503 438 -487 472
rect -887 400 -487 438
rect -429 472 -29 488
rect -429 438 -413 472
rect -45 438 -29 472
rect -429 400 -29 438
rect 29 472 429 488
rect 29 438 45 472
rect 413 438 429 472
rect 29 400 429 438
rect 487 472 887 488
rect 487 438 503 472
rect 871 438 887 472
rect 487 400 887 438
rect -887 -438 -487 -400
rect -887 -472 -871 -438
rect -503 -472 -487 -438
rect -887 -488 -487 -472
rect -429 -438 -29 -400
rect -429 -472 -413 -438
rect -45 -472 -29 -438
rect -429 -488 -29 -472
rect 29 -438 429 -400
rect 29 -472 45 -438
rect 413 -472 429 -438
rect 29 -488 429 -472
rect 487 -438 887 -400
rect 487 -472 503 -438
rect 871 -472 887 -438
rect 487 -488 887 -472
<< polycont >>
rect -871 438 -503 472
rect -413 438 -45 472
rect 45 438 413 472
rect 503 438 871 472
rect -871 -472 -503 -438
rect -413 -472 -45 -438
rect 45 -472 413 -438
rect 503 -472 871 -438
<< locali >>
rect -1047 540 -951 574
rect 951 540 1047 574
rect -1047 478 -1013 540
rect 1013 478 1047 540
rect -887 438 -871 472
rect -503 438 -487 472
rect -429 438 -413 472
rect -45 438 -29 472
rect 29 438 45 472
rect 413 438 429 472
rect 487 438 503 472
rect 871 438 887 472
rect -933 388 -899 404
rect -933 -404 -899 -388
rect -475 388 -441 404
rect -475 -404 -441 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 441 388 475 404
rect 441 -404 475 -388
rect 899 388 933 404
rect 899 -404 933 -388
rect -887 -472 -871 -438
rect -503 -472 -487 -438
rect -429 -472 -413 -438
rect -45 -472 -29 -438
rect 29 -472 45 -438
rect 413 -472 429 -438
rect 487 -472 503 -438
rect 871 -472 887 -438
rect -1047 -540 -1013 -478
rect 1013 -540 1047 -478
rect -1047 -574 -951 -540
rect 951 -574 1047 -540
<< viali >>
rect -834 438 -540 472
rect -376 438 -82 472
rect 82 438 376 472
rect 540 438 834 472
rect -834 -472 -540 -438
rect -376 -472 -82 -438
rect 82 -472 376 -438
rect 540 -472 834 -438
<< metal1 >>
rect -846 472 -528 478
rect -846 438 -834 472
rect -540 438 -528 472
rect -846 432 -528 438
rect -388 472 -70 478
rect -388 438 -376 472
rect -82 438 -70 472
rect -388 432 -70 438
rect 70 472 388 478
rect 70 438 82 472
rect 376 438 388 472
rect 70 432 388 438
rect 528 472 846 478
rect 528 438 540 472
rect 834 438 846 472
rect 528 432 846 438
rect -846 -438 -528 -432
rect -846 -472 -834 -438
rect -540 -472 -528 -438
rect -846 -478 -528 -472
rect -388 -438 -70 -432
rect -388 -472 -376 -438
rect -82 -472 -70 -438
rect -388 -478 -70 -472
rect 70 -438 388 -432
rect 70 -472 82 -438
rect 376 -472 388 -438
rect 70 -478 388 -472
rect 528 -438 846 -432
rect 528 -472 540 -438
rect 834 -472 846 -438
rect 528 -478 846 -472
<< properties >>
string FIXED_BBOX -1030 -557 1030 557
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 2 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
