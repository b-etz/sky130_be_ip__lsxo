magic
tech sky130A
magscale 1 2
timestamp 1713192904
<< pwell >>
rect -1584 -1113 1584 1113
<< mvnmos >>
rect -1356 55 -956 855
rect -778 55 -378 855
rect -200 55 200 855
rect 378 55 778 855
rect 956 55 1356 855
rect -1356 -855 -956 -55
rect -778 -855 -378 -55
rect -200 -855 200 -55
rect 378 -855 778 -55
rect 956 -855 1356 -55
<< mvndiff >>
rect -1414 843 -1356 855
rect -1414 67 -1402 843
rect -1368 67 -1356 843
rect -1414 55 -1356 67
rect -956 843 -898 855
rect -956 67 -944 843
rect -910 67 -898 843
rect -956 55 -898 67
rect -836 843 -778 855
rect -836 67 -824 843
rect -790 67 -778 843
rect -836 55 -778 67
rect -378 843 -320 855
rect -378 67 -366 843
rect -332 67 -320 843
rect -378 55 -320 67
rect -258 843 -200 855
rect -258 67 -246 843
rect -212 67 -200 843
rect -258 55 -200 67
rect 200 843 258 855
rect 200 67 212 843
rect 246 67 258 843
rect 200 55 258 67
rect 320 843 378 855
rect 320 67 332 843
rect 366 67 378 843
rect 320 55 378 67
rect 778 843 836 855
rect 778 67 790 843
rect 824 67 836 843
rect 778 55 836 67
rect 898 843 956 855
rect 898 67 910 843
rect 944 67 956 843
rect 898 55 956 67
rect 1356 843 1414 855
rect 1356 67 1368 843
rect 1402 67 1414 843
rect 1356 55 1414 67
rect -1414 -67 -1356 -55
rect -1414 -843 -1402 -67
rect -1368 -843 -1356 -67
rect -1414 -855 -1356 -843
rect -956 -67 -898 -55
rect -956 -843 -944 -67
rect -910 -843 -898 -67
rect -956 -855 -898 -843
rect -836 -67 -778 -55
rect -836 -843 -824 -67
rect -790 -843 -778 -67
rect -836 -855 -778 -843
rect -378 -67 -320 -55
rect -378 -843 -366 -67
rect -332 -843 -320 -67
rect -378 -855 -320 -843
rect -258 -67 -200 -55
rect -258 -843 -246 -67
rect -212 -843 -200 -67
rect -258 -855 -200 -843
rect 200 -67 258 -55
rect 200 -843 212 -67
rect 246 -843 258 -67
rect 200 -855 258 -843
rect 320 -67 378 -55
rect 320 -843 332 -67
rect 366 -843 378 -67
rect 320 -855 378 -843
rect 778 -67 836 -55
rect 778 -843 790 -67
rect 824 -843 836 -67
rect 778 -855 836 -843
rect 898 -67 956 -55
rect 898 -843 910 -67
rect 944 -843 956 -67
rect 898 -855 956 -843
rect 1356 -67 1414 -55
rect 1356 -843 1368 -67
rect 1402 -843 1414 -67
rect 1356 -855 1414 -843
<< mvndiffc >>
rect -1402 67 -1368 843
rect -944 67 -910 843
rect -824 67 -790 843
rect -366 67 -332 843
rect -246 67 -212 843
rect 212 67 246 843
rect 332 67 366 843
rect 790 67 824 843
rect 910 67 944 843
rect 1368 67 1402 843
rect -1402 -843 -1368 -67
rect -944 -843 -910 -67
rect -824 -843 -790 -67
rect -366 -843 -332 -67
rect -246 -843 -212 -67
rect 212 -843 246 -67
rect 332 -843 366 -67
rect 790 -843 824 -67
rect 910 -843 944 -67
rect 1368 -843 1402 -67
<< mvpsubdiff >>
rect -1548 1065 1548 1077
rect -1548 1031 -1440 1065
rect 1440 1031 1548 1065
rect -1548 1019 1548 1031
rect -1548 969 -1490 1019
rect -1548 -969 -1536 969
rect -1502 -969 -1490 969
rect 1490 969 1548 1019
rect -1548 -1019 -1490 -969
rect 1490 -969 1502 969
rect 1536 -969 1548 969
rect 1490 -1019 1548 -969
rect -1548 -1031 1548 -1019
rect -1548 -1065 -1440 -1031
rect 1440 -1065 1548 -1031
rect -1548 -1077 1548 -1065
<< mvpsubdiffcont >>
rect -1440 1031 1440 1065
rect -1536 -969 -1502 969
rect 1502 -969 1536 969
rect -1440 -1065 1440 -1031
<< poly >>
rect -1356 927 -956 943
rect -1356 893 -1340 927
rect -972 893 -956 927
rect -1356 855 -956 893
rect -778 927 -378 943
rect -778 893 -762 927
rect -394 893 -378 927
rect -778 855 -378 893
rect -200 927 200 943
rect -200 893 -184 927
rect 184 893 200 927
rect -200 855 200 893
rect 378 927 778 943
rect 378 893 394 927
rect 762 893 778 927
rect 378 855 778 893
rect 956 927 1356 943
rect 956 893 972 927
rect 1340 893 1356 927
rect 956 855 1356 893
rect -1356 17 -956 55
rect -1356 -17 -1340 17
rect -972 -17 -956 17
rect -1356 -55 -956 -17
rect -778 17 -378 55
rect -778 -17 -762 17
rect -394 -17 -378 17
rect -778 -55 -378 -17
rect -200 17 200 55
rect -200 -17 -184 17
rect 184 -17 200 17
rect -200 -55 200 -17
rect 378 17 778 55
rect 378 -17 394 17
rect 762 -17 778 17
rect 378 -55 778 -17
rect 956 17 1356 55
rect 956 -17 972 17
rect 1340 -17 1356 17
rect 956 -55 1356 -17
rect -1356 -893 -956 -855
rect -1356 -927 -1340 -893
rect -972 -927 -956 -893
rect -1356 -943 -956 -927
rect -778 -893 -378 -855
rect -778 -927 -762 -893
rect -394 -927 -378 -893
rect -778 -943 -378 -927
rect -200 -893 200 -855
rect -200 -927 -184 -893
rect 184 -927 200 -893
rect -200 -943 200 -927
rect 378 -893 778 -855
rect 378 -927 394 -893
rect 762 -927 778 -893
rect 378 -943 778 -927
rect 956 -893 1356 -855
rect 956 -927 972 -893
rect 1340 -927 1356 -893
rect 956 -943 1356 -927
<< polycont >>
rect -1340 893 -972 927
rect -762 893 -394 927
rect -184 893 184 927
rect 394 893 762 927
rect 972 893 1340 927
rect -1340 -17 -972 17
rect -762 -17 -394 17
rect -184 -17 184 17
rect 394 -17 762 17
rect 972 -17 1340 17
rect -1340 -927 -972 -893
rect -762 -927 -394 -893
rect -184 -927 184 -893
rect 394 -927 762 -893
rect 972 -927 1340 -893
<< locali >>
rect -1536 1031 -1440 1065
rect 1440 1031 1536 1065
rect -1536 969 -1502 1031
rect 1502 969 1536 1031
rect -1356 893 -1340 927
rect -972 893 -956 927
rect -778 893 -762 927
rect -394 893 -378 927
rect -200 893 -184 927
rect 184 893 200 927
rect 378 893 394 927
rect 762 893 778 927
rect 956 893 972 927
rect 1340 893 1356 927
rect -1402 843 -1368 859
rect -1402 51 -1368 67
rect -944 843 -910 859
rect -944 51 -910 67
rect -824 843 -790 859
rect -824 51 -790 67
rect -366 843 -332 859
rect -366 51 -332 67
rect -246 843 -212 859
rect -246 51 -212 67
rect 212 843 246 859
rect 212 51 246 67
rect 332 843 366 859
rect 332 51 366 67
rect 790 843 824 859
rect 790 51 824 67
rect 910 843 944 859
rect 910 51 944 67
rect 1368 843 1402 859
rect 1368 51 1402 67
rect -1356 -17 -1340 17
rect -972 -17 -956 17
rect -778 -17 -762 17
rect -394 -17 -378 17
rect -200 -17 -184 17
rect 184 -17 200 17
rect 378 -17 394 17
rect 762 -17 778 17
rect 956 -17 972 17
rect 1340 -17 1356 17
rect -1402 -67 -1368 -51
rect -1402 -859 -1368 -843
rect -944 -67 -910 -51
rect -944 -859 -910 -843
rect -824 -67 -790 -51
rect -824 -859 -790 -843
rect -366 -67 -332 -51
rect -366 -859 -332 -843
rect -246 -67 -212 -51
rect -246 -859 -212 -843
rect 212 -67 246 -51
rect 212 -859 246 -843
rect 332 -67 366 -51
rect 332 -859 366 -843
rect 790 -67 824 -51
rect 790 -859 824 -843
rect 910 -67 944 -51
rect 910 -859 944 -843
rect 1368 -67 1402 -51
rect 1368 -859 1402 -843
rect -1356 -927 -1340 -893
rect -972 -927 -956 -893
rect -778 -927 -762 -893
rect -394 -927 -378 -893
rect -200 -927 -184 -893
rect 184 -927 200 -893
rect 378 -927 394 -893
rect 762 -927 778 -893
rect 956 -927 972 -893
rect 1340 -927 1356 -893
rect -1536 -1031 -1502 -969
rect 1502 -1031 1536 -969
rect -1536 -1065 -1440 -1031
rect 1440 -1065 1536 -1031
<< viali >>
rect -1303 893 -1009 927
rect -725 893 -431 927
rect -147 893 147 927
rect 431 893 725 927
rect 1009 893 1303 927
rect -1303 -17 -1009 17
rect -725 -17 -431 17
rect -147 -17 147 17
rect 431 -17 725 17
rect 1009 -17 1303 17
rect -1303 -927 -1009 -893
rect -725 -927 -431 -893
rect -147 -927 147 -893
rect 431 -927 725 -893
rect 1009 -927 1303 -893
<< metal1 >>
rect -1315 927 -997 933
rect -1315 893 -1303 927
rect -1009 893 -997 927
rect -1315 887 -997 893
rect -737 927 -419 933
rect -737 893 -725 927
rect -431 893 -419 927
rect -737 887 -419 893
rect -159 927 159 933
rect -159 893 -147 927
rect 147 893 159 927
rect -159 887 159 893
rect 419 927 737 933
rect 419 893 431 927
rect 725 893 737 927
rect 419 887 737 893
rect 997 927 1315 933
rect 997 893 1009 927
rect 1303 893 1315 927
rect 997 887 1315 893
rect -1315 17 -997 23
rect -1315 -17 -1303 17
rect -1009 -17 -997 17
rect -1315 -23 -997 -17
rect -737 17 -419 23
rect -737 -17 -725 17
rect -431 -17 -419 17
rect -737 -23 -419 -17
rect -159 17 159 23
rect -159 -17 -147 17
rect 147 -17 159 17
rect -159 -23 159 -17
rect 419 17 737 23
rect 419 -17 431 17
rect 725 -17 737 17
rect 419 -23 737 -17
rect 997 17 1315 23
rect 997 -17 1009 17
rect 1303 -17 1315 17
rect 997 -23 1315 -17
rect -1315 -893 -997 -887
rect -1315 -927 -1303 -893
rect -1009 -927 -997 -893
rect -1315 -933 -997 -927
rect -737 -893 -419 -887
rect -737 -927 -725 -893
rect -431 -927 -419 -893
rect -737 -933 -419 -927
rect -159 -893 159 -887
rect -159 -927 -147 -893
rect 147 -927 159 -893
rect -159 -933 159 -927
rect 419 -893 737 -887
rect 419 -927 431 -893
rect 725 -927 737 -893
rect 419 -933 737 -927
rect 997 -893 1315 -887
rect 997 -927 1009 -893
rect 1303 -927 1315 -893
rect 997 -933 1315 -927
<< properties >>
string FIXED_BBOX -1519 -1048 1519 1048
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4 l 2 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
