magic
tech sky130A
magscale 1 2
timestamp 1712250795
<< pwell >>
rect -948 -2082 948 2082
<< psubdiff >>
rect -912 2012 -816 2046
rect 816 2012 912 2046
rect -912 1950 -878 2012
rect 878 1950 912 2012
rect -912 -2012 -878 -1950
rect 878 -2012 912 -1950
rect -912 -2046 -816 -2012
rect 816 -2046 912 -2012
<< psubdiffcont >>
rect -816 2012 816 2046
rect -912 -1950 -878 1950
rect 878 -1950 912 1950
rect -816 -2046 816 -2012
<< xpolycontact >>
rect -782 1484 -712 1916
rect -782 -1916 -712 -1484
rect -616 1484 -546 1916
rect -616 -1916 -546 -1484
rect -450 1484 -380 1916
rect -450 -1916 -380 -1484
rect -284 1484 -214 1916
rect -284 -1916 -214 -1484
rect -118 1484 -48 1916
rect -118 -1916 -48 -1484
rect 48 1484 118 1916
rect 48 -1916 118 -1484
rect 214 1484 284 1916
rect 214 -1916 284 -1484
rect 380 1484 450 1916
rect 380 -1916 450 -1484
rect 546 1484 616 1916
rect 546 -1916 616 -1484
rect 712 1484 782 1916
rect 712 -1916 782 -1484
<< xpolyres >>
rect -782 -1484 -712 1484
rect -616 -1484 -546 1484
rect -450 -1484 -380 1484
rect -284 -1484 -214 1484
rect -118 -1484 -48 1484
rect 48 -1484 118 1484
rect 214 -1484 284 1484
rect 380 -1484 450 1484
rect 546 -1484 616 1484
rect 712 -1484 782 1484
<< locali >>
rect -912 2012 -816 2046
rect 816 2012 912 2046
rect -912 1950 -878 2012
rect 878 1950 912 2012
rect -912 -2012 -878 -1950
rect 878 -2012 912 -1950
rect -912 -2046 -816 -2012
rect 816 -2046 912 -2012
<< viali >>
rect -766 1501 -728 1898
rect -600 1501 -562 1898
rect -434 1501 -396 1898
rect -268 1501 -230 1898
rect -102 1501 -64 1898
rect 64 1501 102 1898
rect 230 1501 268 1898
rect 396 1501 434 1898
rect 562 1501 600 1898
rect 728 1501 766 1898
rect -766 -1898 -728 -1501
rect -600 -1898 -562 -1501
rect -434 -1898 -396 -1501
rect -268 -1898 -230 -1501
rect -102 -1898 -64 -1501
rect 64 -1898 102 -1501
rect 230 -1898 268 -1501
rect 396 -1898 434 -1501
rect 562 -1898 600 -1501
rect 728 -1898 766 -1501
<< metal1 >>
rect -772 1898 -722 1910
rect -772 1501 -766 1898
rect -728 1501 -722 1898
rect -772 1489 -722 1501
rect -606 1898 -556 1910
rect -606 1501 -600 1898
rect -562 1501 -556 1898
rect -606 1489 -556 1501
rect -440 1898 -390 1910
rect -440 1501 -434 1898
rect -396 1501 -390 1898
rect -440 1489 -390 1501
rect -274 1898 -224 1910
rect -274 1501 -268 1898
rect -230 1501 -224 1898
rect -274 1489 -224 1501
rect -108 1898 -58 1910
rect -108 1501 -102 1898
rect -64 1501 -58 1898
rect -108 1489 -58 1501
rect 58 1898 108 1910
rect 58 1501 64 1898
rect 102 1501 108 1898
rect 58 1489 108 1501
rect 224 1898 274 1910
rect 224 1501 230 1898
rect 268 1501 274 1898
rect 224 1489 274 1501
rect 390 1898 440 1910
rect 390 1501 396 1898
rect 434 1501 440 1898
rect 390 1489 440 1501
rect 556 1898 606 1910
rect 556 1501 562 1898
rect 600 1501 606 1898
rect 556 1489 606 1501
rect 722 1898 772 1910
rect 722 1501 728 1898
rect 766 1501 772 1898
rect 722 1489 772 1501
rect -772 -1501 -722 -1489
rect -772 -1898 -766 -1501
rect -728 -1898 -722 -1501
rect -772 -1910 -722 -1898
rect -606 -1501 -556 -1489
rect -606 -1898 -600 -1501
rect -562 -1898 -556 -1501
rect -606 -1910 -556 -1898
rect -440 -1501 -390 -1489
rect -440 -1898 -434 -1501
rect -396 -1898 -390 -1501
rect -440 -1910 -390 -1898
rect -274 -1501 -224 -1489
rect -274 -1898 -268 -1501
rect -230 -1898 -224 -1501
rect -274 -1910 -224 -1898
rect -108 -1501 -58 -1489
rect -108 -1898 -102 -1501
rect -64 -1898 -58 -1501
rect -108 -1910 -58 -1898
rect 58 -1501 108 -1489
rect 58 -1898 64 -1501
rect 102 -1898 108 -1501
rect 58 -1910 108 -1898
rect 224 -1501 274 -1489
rect 224 -1898 230 -1501
rect 268 -1898 274 -1501
rect 224 -1910 274 -1898
rect 390 -1501 440 -1489
rect 390 -1898 396 -1501
rect 434 -1898 440 -1501
rect 390 -1910 440 -1898
rect 556 -1501 606 -1489
rect 556 -1898 562 -1501
rect 600 -1898 606 -1501
rect 556 -1910 606 -1898
rect 722 -1501 772 -1489
rect 722 -1898 728 -1501
rect 766 -1898 772 -1501
rect 722 -1910 772 -1898
<< properties >>
string FIXED_BBOX -895 -2029 895 2029
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 15 m 1 nx 10 wmin 0.350 lmin 0.50 rho 2000 val 86.789k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
