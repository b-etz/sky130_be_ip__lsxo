magic
tech sky130A
magscale 1 2
timestamp 1712511904
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 0 1 2982 -1 0 -616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x2
timestamp 1707688321
transform 0 1 9098 -1 0 -780
box -38 -48 314 592
use level_shift  x3
timestamp 1712511643
transform 0 1 4250 -1 0 -1190
box 652 -1950 5670 -128
use level_shift  x4
timestamp 1712511643
transform 0 -1 4086 -1 0 -1188
box 652 -1950 5670 -128
use bias_gen  x5
timestamp 1712250795
transform 1 0 1962 0 1 -15524
box -450 -14480 16732 3256
use dout_amp  x6
timestamp 1712087189
transform 1 0 20214 0 1 -2274
box -1220 -12900 16982 200
use ripl_dly_clk_buf  x7
timestamp 1712087189
transform 1 0 38260 0 1 -6068
box 872 -3046 9184 598
use sky130_fd_pr__cap_mim_m3_1_KAF84V  XC1
timestamp 1712073300
transform -1 0 17850 0 -1 -24526
box -886 -3440 886 3440
use sky130_fd_pr__cap_mim_m3_1_4HJTN9  XC2
timestamp 1712437813
transform 1 0 33062 0 1 -21822
box -7716 -4640 7716 4640
use sky130_fd_pr__cap_mim_m3_1_4DMTN9  XC3
timestamp 1712250795
transform 1 0 12064 0 1 -6736
box -2492 -2320 2492 2320
use sky130_fd_pr__cap_mim_m3_1_4HHTN9  XC4
timestamp 1712073300
transform 0 -1 42836 1 0 -10682
box -1186 -4640 1186 4640
use sky130_fd_pr__nfet_g5v0d10v5_MHWJF7  XM1
timestamp 1712250795
transform 1 0 20755 0 1 -24504
box -989 -658 989 658
use sky130_fd_pr__pfet_g5v0d10v5_28EAA9  XM2
timestamp 1712250795
transform 0 1 20849 -1 0 -21271
box -2519 -697 2519 697
use sky130_fd_pr__nfet_01v8_AHZR5K  XM3
timestamp 1712071977
transform 1 0 39782 0 1 -9680
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_HZ6WG7  XM4
timestamp 1712071977
transform 1 0 46948 0 1 -11363
box -296 -285 296 285
use sky130_fd_pr__nfet_g5v0d10v5_ZPGQJT  XM5
timestamp 1712087189
transform 1 0 2288 0 1 -8894
box -594 -658 594 658
use sky130_fd_pr__pfet_g5v0d10v5_KLKQZ5  XM6
timestamp 1712087189
transform 1 0 4274 0 1 -8937
box -624 -697 624 697
use sky130_fd_pr__pfet_01v8_3H68VM  XM7
timestamp 1712071977
transform 1 0 46810 0 1 -10257
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_XPHWY6  XM8
timestamp 1712087189
transform 1 0 16278 0 1 -1749
box -562 -1137 562 1137
use sky130_fd_pr__pfet_g5v0d10v5_KL3SY6  XM9
timestamp 1712071977
transform 0 1 19719 -1 0 -1200
box -308 -697 308 697
use sky130_fd_pr__nfet_01v8_Y5BWKS  XM11
timestamp 1712087189
transform 1 0 16360 0 1 -4521
box -562 -1119 562 1119
use sky130_fd_pr__res_xhigh_po_0p35_27M88N  XR2
timestamp 1712437813
transform 0 1 12474 -1 0 -27691
box -2359 -10982 2359 10982
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 dvdd
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 dvss
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 ibias
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 ena
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 standby
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 dout
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 xin
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 xout
port 9 nsew
<< end >>
