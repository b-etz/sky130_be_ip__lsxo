* PEX produced on Wed Apr 17 10:14:11 EDT 2024 using /home/brady/sources/osic-multitool-src/iic-pex.sh with m=3 and s=1
* NGSPICE file created from sky130_be_ip__lsxo.ext - technology: sky130A

.subckt sky130_be_ip__lsxo ibias dout xout xin ena avss avdd standby dvss dvdd
X0 a_16620_n1869.t2 a_15705_n2241.t2 a_16273_n2273.t2 dvss.t177 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1 a_20376_n2791.t0 x7.stby_done_b.t2 dvdd.t18 dvdd.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_21036_n1869.t2 a_19955_n2241.t2 a_20689_n2273.t2 dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3 a_10620_n8338.t0 a_24220_n8172.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X4 a_16795_n2817.t0 a_16620_n2791.t4 a_16974_n2791.t0 dvss.t66 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5 dvdd.t5 ena_ip.t2 x3.in_b.t0 dvdd.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X6 dvdd.t46 a_21036_n1869.t4 a_21211_n1943.t0 dvdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_18828_n2791.t1 a_17913_n2791.t2 a_18481_n2549.t1 dvss.t72 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X8 a_2130_n19848.t0 a_24530_n20014.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X9 vbreg.t5 icnode.t0 a_11526_n12394.t1 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X10 x7.x2.x2.CLK.t1 a_15000_n2791.t3 dvss.t78 dvss.t77 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X11 a_18168_n1881.t1 x7.x1.Qb2.t2 dvss.t99 dvss.t98 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X12 tail.t9 vbp.t1 dvdd_ip.t33 dvdd_ip.t23 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X13 a_16317_n2791.t0 a_16273_n2549.t4 a_16151_n2791.t0 dvss.t90 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X14 dvss.t164 standby_b.t0 dvss_ip dvss.t163 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X15 a_9120_n9346.t4 a_24220_n9832.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X16 a_16795_n1943.t1 a_16620_n1869.t4 a_16974_n1881.t0 dvss.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X17 x7.ena_done_b.t0 a_21775_n2247.t2 dvdd.t166 dvdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X18 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X19 a_20121_n2241.t0 a_19955_n2241.t3 dvdd.t71 dvdd.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_2130_n21176.t1 a_24530_n21342.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X21 ibias_ip.t10 standby_33.t3 ibias.t1 ibias.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X22 xout.t22 vbreg.t9 avdd_ip.t28 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X23 inv_m1.t1 inv_in.t1 dvdd_ip.t42 dvdd_ip.t41 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X24 a_2132_n15590.t0 a_18932_n15756.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X25 dout_ip.t3 inv_m2.t2 dvdd_ip.t4 dvdd_ip.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X26 a_20733_n2791.t1 a_20689_n2549.t4 a_20567_n2791.t0 dvss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X27 inv_in.t2 xin_buf.t3 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X28 x7.x1.x2.CLK.t1 a_15000_n1881.t3 dvss.t20 dvss.t19 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X29 avdd_ip.t29 avss_ip sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X30 a_16317_n1881.t1 a_16273_n2273.t4 a_16151_n1869.t0 dvss.t45 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X31 x7.stby_done_b.t1 a_21775_n2791.t2 dvss.t210 dvss.t209 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X32 a_14009_n2701.t1 x7.clk_disable.t2 dvss.t84 dvss.t83 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.07665 ps=0.785 w=0.42 l=0.15
X33 dvss.t31 standby_ip.t2 x4.in_b dvss.t30 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X34 dvss.t42 a_2971_n1521.t2 ena_ip.t0 dvss.t41 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X35 dvss.t166 standby_b.t1 a_16317_n2791.t1 dvss.t165 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X36 avdd_ip.t30 avss_ip sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X37 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X38 dvss.t193 x7.ena_done_b.t2 a_14035_n1997.t1 dvss.t33 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X39 x7.stby_done_b.t0 a_21775_n2791.t3 dvdd.t59 dvdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X40 a_2132_n17582.t1 a_18932_n17416.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X41 inv_m1.t0 inv_in.t3 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X42 avss.t26 avdd.t14 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X43 a_10620_n9666.t0 a_24220_n9832.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X44 a_20733_n1881.t0 a_20689_n2273.t4 a_20567_n1869.t0 dvss.t131 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X45 dvdd.t110 x7.x2.x2.CLK.t2 a_15539_n2791.t0 dvdd.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X46 a_16782_n2425.t1 a_15705_n2791.t2 a_16620_n2791.t0 dvdd.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X47 dvdd_ip.t53 inv_m1.t2 inv_m2.t1 dvdd_ip.t35 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X48 a_4857_n1521.t0 standby.t0 dvdd.t38 dvdd.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X49 avdd_ip.t4 x3.out_b.t3 avdd.t16 avdd.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X50 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X51 a_20121_n2791.t1 a_19955_n2791.t2 dvss.t213 dvss.t212 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X52 dvss.t4 ena_ip.t3 a_16317_n1881.t0 dvss.t3 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X53 x7.x1.Qb2.t0 a_19567_n2247.t2 dvss.t74 dvss.t73 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X54 dvss.t190 ena.t0 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X55 dvdd.t139 a_19003_n2817.t3 a_19567_n2791.t0 dvdd.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X56 avss_ip vg1.t1 vg1.t2 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X57 a_21145_n1869.t0 a_19955_n2241.t4 a_21036_n1869.t3 dvss.t95 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X58 avdd_ip.t21 vbreg.t10 avdd_ip.t20 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X59 a_21211_n2817.t2 standby_b.t2 dvdd.t106 dvdd.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X60 avss_ip xin.t6 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=23.6118 ps=175.6 w=4 l=0.5
X61 a_19003_n2817.t2 a_18828_n2791.t4 a_19182_n2791.t1 dvss.t124 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X62 a_15000_n1881.t1 dout_ip.t4 dvdd.t114 dvdd.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
X63 a_2132_n17250.t1 a_18932_n17416.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X64 a_20121_n2241.t1 a_19955_n2241.t5 dvss.t97 dvss.t96 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X65 dvss_ip ibias_ip.t11 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=5.8 ps=45.8 w=2 l=2
X66 a_10620_n9666.t1 a_24220_n9500.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X67 a_18359_n1869.t0 a_17913_n2241.t2 a_18263_n1869.t2 dvss.t182 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X68 xout.t21 vbreg.t11 avdd_ip.t27 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X69 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=75
X70 vbreg.t8 vg2.t5 vrb.t4 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X71 a_18525_n2791.t0 a_18481_n2549.t4 a_18359_n2791.t0 dvss.t23 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X72 a_2130_n20844.t1 a_24530_n21010.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X73 a_15083_n2791.t1 dout_ip.t5 a_15000_n2791.t1 dvss.t102 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X74 a_21036_n1869.t0 a_20121_n2241.t2 a_20689_n2273.t1 dvss.t44 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X75 dvss_ip standby_b.t3 dvss.t76 dvss.t75 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X76 a_2132_n15590.t1 a_18932_n15424.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X77 a_14285_n2079.t1 x7.ena_done_b.t3 a_14285_n2281.t3 dvdd.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X78 a_19003_n1943.t2 a_18828_n1869.t4 a_19182_n1881.t1 dvss.t69 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X79 vn.t6 xin.t7 vn.t5 dvdd_ip.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X80 avss.t7 standby_b.t4 standby_33.t2 avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X81 a_10620_n7674.t1 a_24220_n7840.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X82 ibias_ip.t9 ibias_ip.t8 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X83 avdd.t5 x3.out_b.t4 avdd_ip.t0 avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X84 a_15960_n2791.t1 x7.x2.Qb1.t2 dvdd.t140 dvdd.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X85 a_2130_n19516.t0 a_24530_n19682.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X86 xin.t8 avdd_ip.t5 sky130_fd_pr__diode_pd2nw_05v5 perim=1.8e+06 area=2.025e+11
X87 a_20579_n2247.t1 ena_ip.t4 dvdd.t167 dvdd.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X88 dvdd.t83 a_2971_n1521.t3 ena_ip.t1 dvdd.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X89 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X90 a_15083_n1881.t1 dout_ip.t6 a_15000_n1881.t2 dvss.t171 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X91 a_18525_n1881.t1 a_18481_n2273.t4 a_18359_n1869.t1 dvss.t154 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X92 a_18168_n2791.t1 x7.x2.Qb2.t2 dvdd.t23 dvdd.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X93 dvss.t65 standby_b.t5 a_18525_n2791.t1 dvss.t64 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X94 xin_buf.t1 xout.t23 tail.t11 dvdd_ip.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X95 a_16273_n2549.t0 a_16055_n2791.t4 dvdd.t89 dvdd.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X96 dvss.t123 x7.stby_done_b.t3 a_15083_n2791.t0 dvss.t122 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X97 xout.t2 xin.t9 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X98 x7.x1.x4.Q.t1 a_21211_n1943.t3 dvss.t113 dvss.t112 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X99 dvdd.t16 x7.stby_done_b.t4 a_15000_n2791.t0 dvdd.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X100 a_14009_n2404.t2 standby_ip.t3 a_14285_n2079.t2 dvdd.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X101 dvss_ip standby_b.t6 dvss.t158 dvss.t157 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X102 avdd_ip.t26 vbreg.t12 xout.t20 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X103 tail.t8 vbp.t2 dvdd_ip.t32 dvdd_ip.t13 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X104 a_2130_n20844.t0 a_24530_n20678.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X105 a_16729_n1869.t1 a_15539_n2241.t2 a_16620_n1869.t3 dvss.t194 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X106 avss_ip vg2.t3 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X107 dvdd_ip.t31 vbp.t3 dvdd_ip.t30 dvdd_ip.t10 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X108 a_16273_n2273.t3 a_16055_n1869.t4 dvdd.t162 dvdd.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X109 a_2132_n15258.t0 a_18932_n15424.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X110 a_18990_n2425.t1 a_17913_n2791.t3 a_18828_n2791.t2 dvdd.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X111 a_14285_n2281.t0 x7.stby_done_b.t5 dvdd.t14 dvdd.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X112 avdd_ip.t25 vbreg.t13 avdd_ip.t24 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X113 dvss.t201 ena_ip.t5 a_18525_n1881.t0 dvss.t200 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X114 dvdd.t124 a_21211_n1943.t4 a_21775_n2247.t0 dvdd.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X115 dvss.t144 x7.ena_done_b.t4 a_15083_n1881.t0 dvss.t143 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X116 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X117 a_16795_n1943.t2 ena_ip.t6 dvdd.t127 dvdd.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X118 dvss.t108 standby.t1 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X119 dvss.t160 standby_b.t7 dvss_ip dvss.t159 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X120 a_2130_n19516.t1 a_24530_n19350.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X121 dvdd.t87 a_14009_n2404.t4 x7.clk_disable.t0 dvdd.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X122 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X123 dvdd_ip.t47 standby_ip.t4 dvdd.t116 dvdd.t115 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X124 a_16163_n2247.t0 ena_ip.t7 dvdd.t128 dvdd.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X125 a_2132_n16918.t0 a_18932_n17084.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X126 dvdd.t135 x7.x2.Qb2.t3 a_19955_n2791.t1 dvdd.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X127 a_19003_n1943.t0 ena_ip.t8 dvdd.t130 dvdd.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X128 inv_in.t4 xin_buf.t3 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X129 a_10620_n9334.t1 a_24220_n9500.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X130 dvss.t53 a_21211_n2817.t3 a_21775_n2791.t1 dvss.t52 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X131 a_3134_n13324.t0 vrb.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=75
X132 dvdd_ip.t48 standby_ip.t5 dvdd.t118 dvdd.t117 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X133 a_16974_n2791.t1 standby_b.t8 dvss.t92 dvss.t91 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X134 x7.x1.x2.Q.t1 a_16795_n1943.t3 dvss.t38 dvss.t37 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X135 a_2132_n17582.t0 a_18932_n17748.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X136 dvdd.t173 x7.x1.x2.CLK.t2 a_15539_n2241.t0 dvdd.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X137 dvdd_ip.t29 vbp.t4 tail.t7 dvdd_ip.t8 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X138 a_19182_n2791.t0 standby_b.t9 dvss.t94 dvss.t93 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X139 dvss.t105 a_19003_n2817.t4 a_18937_n2791.t0 dvss.t104 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X140 avss_ip avss_ip avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X141 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X142 dout_ip.t1 inv_m2.t3 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X143 a_15705_n2791.t0 a_15539_n2791.t2 dvdd.t56 dvdd.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X144 avdd.t6 x3.out_b.t5 x3.out.t2 avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X145 dvdd.t29 a_16795_n2817.t3 a_16782_n2425.t0 dvdd.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X146 dvss.t138 a_21211_n1943.t5 a_21775_n2247.t1 dvss.t137 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X147 xout.t10 xin.t10 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X148 avss_ip avss_ip avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X149 a_16974_n1881.t1 ena_ip.t9 dvss.t130 dvss.t129 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X150 dvdd.t66 a_16795_n1943.t4 a_17359_n2247.t0 dvdd.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X151 xin.t0 a_24530_n22338.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X152 avss_ip x3.out.t3 avss.t9 avss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X153 dvss.t86 x7.clk_disable.t3 dout_filt.t0 dvss.t85 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X154 a_16055_n2791.t1 a_15539_n2791.t3 a_15960_n2791.t0 dvss.t134 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X155 dvdd.t36 standby_ip.t6 dvdd_ip.t34 dvdd.t35 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X156 standby_33.t0 x4.out_b.t3 avdd.t1 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X157 a_16055_n1869.t2 a_15705_n2241.t3 a_15960_n1881.t3 dvdd.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X158 dvdd_ip.t28 vbp.t5 tail.t6 dvdd_ip.t19 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X159 a_20471_n2791.t2 a_20121_n2791.t2 a_20376_n2791.t2 dvdd.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X160 avss_ip xout.t24 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
**devattr s=257843176,88584 d=257843176,88584
X161 tail.t5 vbp.t6 dvdd_ip.t27 dvdd_ip.t17 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X162 dvdd.t136 a_19003_n2817.t5 a_18990_n2425.t0 dvdd.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X163 a_10620_n9334.t0 a_24220_n9168.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X164 a_19182_n1881.t0 ena_ip.t10 dvss.t150 dvss.t149 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X165 avdd_ip.t23 vbreg.t14 xout.t19 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X166 avss_ip xin.t11 xout.t6 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X167 xin_buf.t0 xout.t25 xin_buf.t0 dvdd_ip.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0 ps=0 w=4 l=2
X168 a_3134_n13324.t1 avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=75
X169 a_21036_n2791.t1 a_19955_n2791.t3 a_20689_n2549.t3 dvdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X170 dvss.t49 a_19003_n1943.t3 a_18937_n1869.t1 dvss.t48 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X171 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X172 a_18937_n2791.t1 a_17747_n2791.t2 a_18828_n2791.t0 dvss.t87 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X173 dvss.t63 a_16795_n2817.t4 a_17359_n2791.t1 dvss.t62 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X174 a_16273_n2273.t0 a_16055_n1869.t5 dvss.t51 dvss.t50 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X175 dvdd.t12 a_16620_n1869.t5 a_16795_n1943.t0 dvdd.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X176 x7.x1.x2.Q.t0 a_16795_n1943.t5 dvdd.t151 dvdd.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X177 a_2130_n20512.t1 a_24530_n20678.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X178 avss_ip xin.t12 xout.t8 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X179 dvdd.t9 a_21036_n2791.t4 a_21211_n2817.t1 dvdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X180 x4.out_b.t2 standby_ip.t7 avss.t23 avss.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X181 a_18481_n2549.t0 a_18263_n2791.t4 dvdd.t77 dvdd.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X182 dvss_ip inv_m1.t3 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=7.9025 ps=61.46 w=0.5 l=1
X183 ibias_ip.t7 ibias_ip.t6 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X184 dvss.t181 x7.x2.x2.CLK.t3 a_15539_n2791.t1 dvss.t180 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X185 xout.t7 xin.t13 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X186 a_2132_n14926.t1 a_18932_n15092.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X187 dvdd.t52 x7.clk_disable.t4 a_14357_n2743.t0 dvdd.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.005 as=0.0672 ps=0.85 w=0.64 l=0.15
X188 vn.t4 vn.t2 vn.t3 dvss_ip sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X189 a_20567_n2791.t1 a_20121_n2791.t3 a_20471_n2791.t3 dvss.t189 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X190 dvdd.t143 standby_ip.t8 dvdd_ip.t50 dvdd.t142 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X191 dvss_ip dout_filt.t3 dout.t0 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=1
X192 a_20471_n1869.t0 a_19955_n2241.t6 a_20376_n1881.t0 dvss.t211 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X193 a_18481_n2273.t1 a_18263_n1869.t4 dvdd.t125 dvdd.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X194 avss.t19 x3.out.t4 avss_ip avss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X195 dvss.t169 a_16795_n1943.t6 a_17359_n2247.t1 dvss.t168 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X196 x7.x1.Qb1.t0 a_17359_n2247.t2 dvdd.t1 dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X197 dvdd_ip.t26 vbp.t7 tail.t4 dvdd_ip.t15 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X198 avss.t27 avdd.t13 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X199 x7.x2.x2.Q.t0 a_16795_n2817.t5 dvdd.t99 dvdd.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X200 a_14035_n2743.t1 dout_ip.t7 dout_filt.t1 dvss.t83 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X201 dvss.t208 x7.x1.x2.CLK.t3 a_15539_n2241.t1 dvss.t207 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X202 dout_ip.t0 inv_m2.t4 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X203 xin_buf.t4 vn.t8 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X204 avdd_ip.t22 vbreg.t15 vg1.t3 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X205 a_2130_n19848.t1 a_24530_n19682.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X206 vrb.t3 vg2.t6 vbreg.t0 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X207 a_18828_n1869.t1 a_17913_n2241.t3 a_18481_n2273.t0 dvss.t148 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X208 x7.x2.Qb1.t1 a_17359_n2791.t2 dvss.t142 dvss.t141 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X209 a_2130_n20512.t0 a_24530_n20346.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X210 dvdd.t67 a_20689_n2273.t5 a_20579_n2247.t0 dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X211 x7.x1.x2.CLK.t0 a_15000_n1881.t4 dvdd.t34 dvdd.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X212 dvdd_ip.t51 standby_ip.t9 dvdd.t145 dvdd.t144 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X213 a_2132_n14926.t0 a_18932_n14760.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X214 x7.x2.Qb1.t0 a_17359_n2791.t3 dvdd.t91 dvdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X215 x7.x1.x3.Q.t1 a_19003_n1943.t4 dvss.t119 dvss.t118 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X216 xout.t4 xin.t14 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X217 avdd.t8 x3.out_b.t6 avdd_ip.t1 avdd.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X218 a_16273_n2549.t2 a_16055_n2791.t5 dvss.t140 dvss.t139 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X219 a_16151_n2791.t1 a_15705_n2791.t3 a_16055_n2791.t3 dvss.t34 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X220 vg1.t4 xin.t5 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X221 avss_ip xin.t15 xout.t1 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X222 dvss_ip inv_m1.t4 inv_m2.t0 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X223 a_2130_n19184.t0 a_24530_n19018.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X224 dvdd_ip.t25 vbp.t8 dvdd_ip.t24 dvdd_ip.t23 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X225 inv_in.t5 xin_buf.t3 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X226 dvdd.t153 a_4857_n1521.t2 standby_ip.t1 dvdd.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X227 a_14035_n1997.t0 ena_ip.t11 a_14009_n2404.t1 dvss.t33 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X228 a_17913_n2791.t1 a_17747_n2791.t3 dvdd.t168 dvdd.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X229 a_4857_n1521.t1 standby.t2 dvss.t109 dvss.t106 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X230 a_10620_n9002.t0 a_24220_n9168.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X231 a_18263_n2791.t0 a_17747_n2791.t4 a_18168_n2791.t0 dvss.t58 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X232 a_14009_n2404.t0 standby_b.t10 a_14035_n2281.t1 dvss.t33 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X233 a_16620_n1869.t0 a_15539_n2241.t3 a_16273_n2273.t1 dvdd.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X234 a_18263_n1869.t1 a_17913_n2241.t4 a_18168_n1881.t2 dvdd.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X235 a_10620_n9002.t1 a_24220_n8836.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X236 dvdd.t112 x7.x1.Qb2.t3 a_19955_n2241.t0 dvdd.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X237 a_2130_n20180.t1 a_24530_n20346.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X238 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X239 x3.out_b.t0 x3.out.t5 avdd.t3 avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X240 xout.t5 xin.t16 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X241 avdd.t17 standby_33.t4 x4.out_b.t0 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
X242 a_20579_n2247.t2 a_19955_n2241.t7 a_20471_n1869.t1 dvdd.t174 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X243 dvdd.t85 a_16273_n2273.t5 a_16163_n2247.t1 dvdd.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X244 a_15000_n2791.t2 dout_ip.t8 dvdd.t133 dvdd.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
X245 dvdd.t40 a_18828_n1869.t5 a_19003_n1943.t1 dvdd.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X246 a_2130_n22172.t1 a_24530_n22006.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X247 avss_ip xin.t17 xout.t0 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X248 avdd_ip.t31 avss_ip sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X249 a_15705_n2241.t1 a_15539_n2241.t4 dvdd.t161 dvdd.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X250 a_2130_n21840.t0 a_24530_n22006.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X251 avdd_ip.t19 vbreg.t16 xout.t18 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X252 dvdd.t123 x7.x2.Qb1.t3 a_17747_n2791.t0 dvdd.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X253 a_2132_n16586.t1 a_18932_n16420.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X254 avss_ip xin.t18 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X255 a_10620_n8670.t1 a_24220_n8836.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X256 xin_buf.t2 vn.t9 xin_buf.t2 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0 ps=0 w=4 l=2
X257 x7.x1.Qb2.t1 a_19567_n2247.t3 dvdd.t158 dvdd.t146 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X258 a_2132_n17250.t0 a_18932_n17084.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X259 a_14009_n2701.t0 x7.clk_disable.t5 dvdd.t54 dvdd.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.10855 ps=1.005 w=0.42 l=0.15
X260 dvss.t68 x7.x2.Qb2.t4 a_19955_n2791.t0 dvss.t67 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X261 dvss.t203 standby_ip.t10 x7.clkin dvss.t202 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X262 dvss_ip ibias_ip.t12 vbp dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X263 inv_in.t6 xin_buf.t3 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X264 a_22601_n15524.t1 vbreg.t17 a_22601_n15524.t0 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X265 a_20579_n2425.t0 standby_b.t11 dvdd.t48 dvdd.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X266 a_16163_n2247.t2 a_15539_n2241.t5 a_16055_n1869.t0 dvdd.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X267 avss_ip xin.t19 xout.t9 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X268 x7.x2.Qb2.t1 a_19567_n2791.t2 dvss.t199 dvss.t198 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X269 vbreg.t4 vg1.t5 vbreg.t3 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X270 vg1.t6 xin.t4 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X271 avss_ip x3.out.t6 avss.t15 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X272 x3.in_b.t1 ena_ip.t12 dvss.t162 dvss.t161 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X273 x7.x2.Qb2.t0 a_19567_n2791.t3 dvdd.t147 dvdd.t146 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X274 dvss.t179 x7.x1.Qb2.t4 a_19955_n2241.t1 dvss.t178 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X275 a_15705_n2791.t1 a_15539_n2791.t4 dvss.t136 dvss.t135 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X276 standby_33.t1 standby_b.t12 avss.t5 avss.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X277 vbreg.t1 vg2.t7 vrb.t2 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X278 tail.t10 xin.t20 vn.t7 dvdd_ip.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X279 dout_ip.t2 inv_m2.t5 dvdd_ip.t1 dvdd_ip.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X280 dvdd.t175 dvss.t170 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X281 dvdd.t138 a_21211_n1943.t6 a_21198_n2247.t1 dvdd.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X282 a_2130_n20180.t0 a_24530_n20014.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X283 dvdd_ip.t22 vbp.t9 dvdd_ip.t21 dvdd_ip.t5 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X284 a_20376_n2791.t1 x7.stby_done_b.t6 dvss.t152 dvss.t151 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X285 a_18828_n1869.t3 a_17747_n2241.t2 a_18481_n2273.t3 dvdd.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X286 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X287 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X288 a_16795_n2817.t2 standby_b.t13 dvdd.t129 dvdd.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X289 a_2132_n14594.t0 a_18932_n14428.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X290 a_15705_n2241.t0 a_15539_n2241.t6 dvss.t101 dvss.t100 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X291 x3.out.t1 x3.in_b.t2 avss.t3 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X292 a_16163_n2425.t1 standby_b.t14 dvdd.t73 dvdd.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X293 inv_in.t7 xin_buf.t3 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X294 a_2132_n15258.t1 a_18932_n15092.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X295 a_19003_n2817.t0 standby_b.t15 dvdd.t75 dvdd.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X296 dvdd.t163 a_18481_n2273.t5 a_18371_n2247.t1 dvdd.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X297 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X298 a_20376_n1881.t2 x7.ena_done_b.t5 dvss.t146 dvss.t145 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X299 dvdd_ip.t37 inv_m1.t5 dvdd_ip.t36 dvdd_ip.t35 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=1
X300 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X301 dvss.t184 standby_b.t16 dvss_ip dvss.t183 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X302 vg1.t7 xin.t3 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X303 a_2130_n19184.t1 a_24530_n19350.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X304 a_10620_n8670.t0 a_24220_n8504.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X305 a_17913_n2241.t1 a_17747_n2241.t3 dvdd.t165 dvdd.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X306 x7.x2.x4.Q.t1 a_21211_n2817.t4 dvss.t29 dvss.t28 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X307 dvss_ip ibias_ip.t4 ibias_ip.t5 dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X308 a_21198_n2247.t0 a_20121_n2241.t3 a_21036_n1869.t1 dvdd.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X309 a_20689_n2273.t0 a_20471_n1869.t4 dvss.t40 dvss.t39 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X310 x7.x1.x4.Q.t0 a_21211_n1943.t7 dvdd.t103 dvdd.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X311 xout.t12 vbreg.t18 xout.t11 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X312 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X313 a_2132_n16918.t1 a_18932_n16752.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X314 avss_ip vg2.t2 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X315 a_16055_n2791.t2 a_15705_n2791.t4 a_15960_n2791.t3 dvdd.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X316 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=75
X317 avss.t1 x3.in_b.t3 x3.out.t0 avss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X318 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X319 dvss_ip standby_b.t17 dvss.t186 dvss.t185 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X320 a_18371_n2247.t0 ena_ip.t13 dvdd.t149 dvdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X321 a_2130_n21508.t1 a_24530_n21674.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X322 a_18371_n2247.t2 a_17747_n2241.t4 a_18263_n1869.t0 dvdd.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X323 vbreg.t7 vbreg.t6 avdd_ip.t18 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X324 a_16620_n2791.t3 a_15705_n2791.t5 a_16273_n2549.t3 dvss.t167 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X325 x7.x2.x4.Q.t0 a_21211_n2817.t5 dvdd.t148 dvdd.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X326 dvdd.t101 a_16620_n2791.t5 a_16795_n2817.t1 dvdd.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X327 dvss_ip standby_b.t18 dvss.t173 dvss.t172 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X328 a_2130_n22172.t0 a_24530_n22338.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X329 a_10620_n8338.t1 a_24220_n8504.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X330 dvdd.t172 x7.x1.Qb1.t2 a_17747_n2241.t0 dvdd.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X331 dvdd.t170 standby_ip.t11 dvdd_ip.t55 dvdd.t169 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X332 inv_in.t8 xin_buf.t3 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X333 a_2132_n16586.t0 a_18932_n16752.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X334 a_17913_n2791.t0 a_17747_n2791.t5 dvss.t12 dvss.t11 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X335 a_16055_n1869.t1 a_15539_n2241.t7 a_15960_n1881.t2 dvss.t18 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X336 x7.x2.x2.Q.t1 a_16795_n2817.t6 dvss.t57 dvss.t56 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X337 avdd_ip.t32 avss_ip sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X338 x7.ena_done_b.t1 a_21775_n2247.t3 dvss.t121 dvss.t120 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X339 avss_ip vg2.t1 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X340 avss_ip avss_ip avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X341 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X342 a_20689_n2549.t1 a_20471_n2791.t4 dvss.t6 dvss.t5 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X343 dvss.t175 standby_b.t19 dvss_ip dvss.t174 sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X344 dvdd.t121 a_19003_n1943.t5 a_19567_n2247.t1 dvdd.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X345 dvdd_ip.t46 a_9120_n9346.t2 a_9120_n9346.t3 dvdd_ip.t45 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X346 dvdd.t32 a_21211_n2817.t6 a_21775_n2791.t0 dvdd.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X347 a_20376_n1881.t1 x7.ena_done_b.t6 dvdd.t61 dvdd.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X348 a_18937_n1869.t0 a_17747_n2241.t5 a_18828_n1869.t2 dvss.t103 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X349 avss_ip xin.t21 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
**devattr s=257843176,88584 d=257843176,88584
X350 dvdd_ip.t20 vbp.t10 tail.t3 dvdd_ip.t19 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X351 a_21211_n2817.t0 a_21036_n2791.t5 a_21390_n2791.t1 dvss.t7 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X352 tail.t2 vbp.t11 dvdd_ip.t18 dvdd_ip.t17 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X353 a_17913_n2241.t0 a_17747_n2241.t6 dvss.t22 dvss.t21 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X354 dvdd.t3 a_20689_n2549.t5 a_20579_n2425.t2 dvdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X355 dvdd_ip.t39 standby_ip.t12 dvdd.t50 dvdd.t49 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X356 a_20567_n1869.t1 a_20121_n2241.t4 a_20471_n1869.t2 dvss.t147 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X357 dvdd.t176 dvss.t114 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X358 dvss.t25 a_19003_n2817.t6 a_19567_n2791.t1 dvss.t24 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X359 a_18481_n2273.t2 a_18263_n1869.t5 dvss.t196 dvss.t195 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X360 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X361 dvss_ip vn.t0 vn.t1 dvss_ip sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X362 a_2130_n18852.t0 a_24530_n19018.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X363 dvss.t55 x7.x2.Qb1.t4 a_17747_n2791.t1 dvss.t54 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X364 dvdd.t177 dvss.t115 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X365 avss.t28 avdd.t12 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X366 avss.t21 standby_ip.t13 x4.out_b.t1 avss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X367 icnode.t1 vg2.t8 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X368 avdd_ip.t17 vbreg.t19 xout.t17 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X369 a_21211_n1943.t1 a_21036_n1869.t5 a_21390_n1881.t0 dvss.t32 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X370 a_15960_n2791.t2 x7.x2.Qb1.t5 dvss.t80 dvss.t79 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X371 a_11526_n12394.t0 icnode.t0 a_8268_n12482.t1 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X372 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X373 dvss.t47 a_19003_n1943.t6 a_19567_n2247.t0 dvss.t46 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X374 xout.t16 vbreg.t20 avdd_ip.t16 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X375 dvss.t107 a_4857_n1521.t3 standby_ip.t0 dvss.t106 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X376 a_14009_n2404.t3 standby_ip.t14 dvss.t59 dvss.t33 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X377 inv_in.t9 xin_buf.t3 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X378 dvdd_ip.t16 vbp.t0 vbp dvdd_ip.t15 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X379 a_2132_n14594.t1 a_18932_n14760.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X380 a_16620_n2791.t2 a_15539_n2791.t5 a_16273_n2549.t1 dvdd.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X381 dvss.t89 x7.x1.Qb1.t3 a_17747_n2241.t1 dvss.t88 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X382 a_18263_n2791.t2 a_17913_n2791.t4 a_18168_n2791.t3 dvdd.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X383 dvdd.t90 a_16795_n2817.t7 a_17359_n2791.t0 dvdd.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X384 a_2971_n1521.t1 ena.t1 dvss.t192 dvss.t191 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X385 dvss.t126 standby_b.t20 a_20733_n2791.t0 dvss.t125 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X386 a_15960_n1881.t0 x7.x1.Qb1.t4 dvss.t27 dvss.t26 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X387 a_14035_n2281.t0 x7.stby_done_b.t7 dvss.t153 dvss.t33 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X388 a_20579_n2425.t1 a_19955_n2791.t4 a_20471_n2791.t0 dvdd.t174 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X389 a_21145_n2791.t0 a_19955_n2791.t5 a_21036_n2791.t0 dvss.t10 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X390 dvdd.t100 a_16273_n2549.t5 a_16163_n2425.t0 dvdd.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X391 a_16151_n1869.t1 a_15705_n2241.t4 a_16055_n1869.t3 dvss.t176 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X392 a_2130_n18852.t1 xout.t3 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X393 dvdd.t97 a_18828_n2791.t5 a_19003_n2817.t1 dvdd.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X394 a_16782_n2247.t1 a_15705_n2241.t5 a_16620_n1869.t1 dvdd.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X395 x3.out_b.t2 ena_ip.t14 avss.t13 avss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
X396 dvss.t197 a_14009_n2404.t5 x7.clk_disable.t1 dvss.t33 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X397 avss.t29 avdd.t11 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X398 dvdd.t95 standby_ip.t15 dvdd_ip.t44 dvdd.t94 sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X399 a_18481_n2549.t2 a_18263_n2791.t5 dvss.t206 dvss.t205 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X400 a_18359_n2791.t1 a_17913_n2791.t5 a_18263_n2791.t3 dvss.t17 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X401 avdd_ip.t2 x3.out_b.t7 avdd.t10 avdd.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X402 a_18263_n1869.t3 a_17747_n2241.t7 a_18168_n1881.t3 dvss.t204 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X403 dvss.t111 ena_ip.t15 a_20733_n1881.t1 dvss.t110 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X404 x7.x2.x3.Q.t1 a_19003_n2817.t7 dvss.t82 dvss.t81 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X405 xout.t15 vbreg.t21 avdd_ip.t15 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X406 avss_ip avss_ip avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X407 x7.x1.x3.Q.t0 a_19003_n1943.t7 dvdd.t45 dvdd.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X408 a_21036_n2791.t3 a_20121_n2791.t4 a_20689_n2549.t2 dvss.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X409 dvss.t128 standby_b.t21 dvss_ip dvss.t127 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X410 avdd_ip.t33 icnode.t0 sky130_fd_pr__cap_mim_m3_1 l=20 w=20
X411 a_21211_n1943.t2 ena_ip.t16 dvdd.t159 dvdd.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X412 inv_in.t10 xin_buf.t3 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X413 inv_in.t11 xin_buf.t3 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X414 a_10620_n8006.t0 a_24220_n8172.t1 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X415 avdd_ip.t14 vbreg.t22 xout.t14 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X416 a_2130_n21840.t1 a_24530_n21674.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X417 inv_in.t12 xin_buf.t3 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X418 a_10620_n8006.t1 a_24220_n7840.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X419 avdd.t19 x3.out_b.t8 avdd_ip.t6 avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X420 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X421 avss.t11 ena_ip.t17 x3.out_b.t1 avss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X422 a_2132_n16254.t1 a_18932_n16420.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X423 a_16163_n2425.t2 a_15539_n2791.t6 a_16055_n2791.t0 dvdd.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X424 tail.t1 vbp.t12 dvdd_ip.t14 dvdd_ip.t13 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X425 a_8268_n12482.t1 a_8268_n12482.t0 avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X426 x7.x2.x3.Q.t0 a_19003_n2817.t8 dvdd.t108 dvdd.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X427 dvss.t117 a_14009_n2701.t2 a_14035_n2743.t0 dvss.t83 sky130_fd_pr__nfet_01v8 ad=0.07665 pd=0.785 as=0.0441 ps=0.63 w=0.42 l=0.15
X428 x7.x2.x2.CLK.t0 a_15000_n2791.t4 dvdd.t107 dvdd.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X429 dvdd_ip.t12 vbp.t13 dvdd_ip.t11 dvdd_ip.t10 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X430 a_21390_n2791.t0 standby_b.t22 dvss.t14 dvss.t13 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X431 dvss.t133 a_21211_n2817.t7 a_21145_n2791.t1 dvss.t132 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X432 vg1.t8 xin.t2 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X433 dvss_ip standby_b.t23 dvss.t16 dvss.t15 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X434 inv_in.t13 xin_buf.t3 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X435 a_16729_n2791.t1 a_15539_n2791.t7 a_16620_n2791.t1 dvss.t43 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X436 a_9120_n9346.t1 a_9120_n9346.t0 dvss_ip dvss_ip sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X437 a_2130_n21176.t0 a_24530_n21010.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X438 a_2132_n17914.t0 vg1.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X439 a_15960_n1881.t1 x7.x1.Qb1.t5 dvdd.t42 dvdd.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X440 a_20121_n2791.t0 a_19955_n2791.t6 dvdd.t21 dvdd.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X441 dvdd.t171 a_21211_n2817.t8 a_21198_n2425.t0 dvdd.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X442 a_14357_n2743.t1 dout_ip.t9 dout_filt.t2 dvdd.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1664 ps=1.8 w=0.64 l=0.15
X443 a_2971_n1521.t0 ena.t2 dvdd.t157 dvdd.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X444 a_21390_n1881.t1 ena_ip.t18 dvss.t188 dvss.t187 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X445 x4.in_b standby_ip.t16 dvdd.t79 dvdd.t78 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X446 dvss_ip ibias_ip.t2 ibias_ip.t3 dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X447 avss_ip x3.out.t7 avss.t25 avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X448 a_18828_n2791.t3 a_17747_n2791.t6 a_18481_n2549.t3 dvdd.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X449 a_18168_n1881.t0 x7.x1.Qb2.t5 dvdd.t154 dvdd.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X450 dvdd.t178 dvss.t116 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X451 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X452 dvss.t71 a_21211_n1943.t8 a_21145_n1869.t1 dvss.t70 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X453 a_14285_n2281.t2 ena_ip.t19 a_14285_n2079.t0 dvdd.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X454 avdd_ip.t13 vbreg.t23 avdd_ip.t12 avdd_ip.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X455 a_2132_n16254.t0 a_18932_n16088.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X456 a_20689_n2549.t0 a_20471_n2791.t5 dvdd.t7 dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X457 dvdd.t62 x7.ena_done_b.t7 a_15000_n1881.t0 dvdd.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X458 dvdd.t25 standby_b.t24 a_14285_n2281.t1 dvdd.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X459 dvdd.t64 a_18481_n2549.t5 a_18371_n2425.t0 dvdd.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X460 dvdd_ip.t9 vbp.t14 tail.t0 dvdd_ip.t8 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X461 xout.t13 vbreg.t24 avdd_ip.t10 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X462 a_18990_n2247.t0 a_17913_n2241.t5 a_18828_n1869.t0 dvdd.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X463 a_20689_n2273.t3 a_20471_n1869.t5 dvdd.t96 dvdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X464 dvss_ip ibias_ip.t13 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X465 vg1.t9 xin.t1 sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X466 avss.t17 x3.out.t8 avss_ip avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X467 avss_ip avss_ip avss_ip avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X468 a_2132_n17914.t1 a_18932_n17748.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X469 a_2132_n14262.t1 a_18932_n14428.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X470 a_21198_n2425.t1 a_20121_n2791.t5 a_21036_n2791.t2 dvdd.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X471 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X472 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X473 dvss.t61 a_16795_n2817.t8 a_16729_n2791.t0 dvss.t60 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X474 inv_in.t14 xin_buf.t3 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X475 dvdd_ip.t7 vbp.t15 dvdd_ip.t6 dvdd_ip.t5 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=2
X476 dvdd_ip.t40 standby_ip.t17 dvdd.t81 dvdd.t80 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X477 avss_ip vg2.t0 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X478 a_2132_n15922.t0 a_18932_n16088.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X479 a_18371_n2425.t1 standby_b.t25 dvdd.t27 dvdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X480 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X481 a_18371_n2425.t2 a_17747_n2791.t7 a_18263_n2791.t1 dvdd.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X482 ibias_ip.t1 ibias_ip.t0 dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X483 dvss.t36 a_16795_n1943.t7 a_16729_n1869.t0 dvss.t35 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X484 dout.t1 dout_filt.t4 dvdd_ip.t3 dvdd_ip.t2 sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X485 a_2132_n14262.t0 vg2.t4 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
X486 dvdd.t60 a_16795_n1943.t8 a_16782_n2247.t0 dvdd.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X487 avdd_ip.t9 vbreg.t25 avdd_ip.t8 avdd_ip.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=2
X488 xout.t26 avdd_ip.t3 sky130_fd_pr__diode_pd2nw_05v5 perim=1.8e+06 area=2.025e+11
X489 a_20471_n2791.t1 a_19955_n2791.t7 a_20376_n2791.t3 dvss.t214 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X490 x7.x1.Qb1.t1 a_17359_n2247.t3 dvss.t2 dvss.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X491 a_20471_n1869.t3 a_20121_n2241.t5 a_20376_n1881.t3 dvdd.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X492 dvdd.t93 standby_ip.t18 dvdd_ip.t43 dvdd.t92 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X493 a_2130_n21508.t0 a_24530_n21342.t0 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=110
X494 a_10620_n7674.t0 inv_in.t0 dvss_ip sky130_fd_pr__res_xhigh_po_0p35 l=66
X495 dvdd.t69 a_19003_n1943.t8 a_18990_n2247.t1 dvdd.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X496 dvdd_ip.t56 dvss_ip sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X497 a_18168_n2791.t2 x7.x2.Qb2.t5 dvss.t156 dvss.t155 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X498 vrb.t1 vg2.t9 vbreg.t2 avss_ip sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X499 a_2132_n15922.t1 a_18932_n15756.t1 avss_ip sky130_fd_pr__res_xhigh_po_0p35 l=82
R0 a_15705_n2241.t1 a_15705_n2241.n3 370.026
R1 a_15705_n2241.n0 a_15705_n2241.t2 351.356
R2 a_15705_n2241.n1 a_15705_n2241.t4 334.717
R3 a_15705_n2241.n3 a_15705_n2241.t0 325.971
R4 a_15705_n2241.n1 a_15705_n2241.t3 309.935
R5 a_15705_n2241.n0 a_15705_n2241.t5 305.683
R6 a_15705_n2241.n2 a_15705_n2241.n0 16.879
R7 a_15705_n2241.n3 a_15705_n2241.n2 10.8867
R8 a_15705_n2241.n2 a_15705_n2241.n1 9.3005
R9 a_16273_n2273.n3 a_16273_n2273.n2 647.119
R10 a_16273_n2273.n1 a_16273_n2273.t4 350.253
R11 a_16273_n2273.n2 a_16273_n2273.n0 260.339
R12 a_16273_n2273.n2 a_16273_n2273.n1 246.119
R13 a_16273_n2273.n1 a_16273_n2273.t5 189.588
R14 a_16273_n2273.n3 a_16273_n2273.t1 89.1195
R15 a_16273_n2273.n0 a_16273_n2273.t2 63.3338
R16 a_16273_n2273.t3 a_16273_n2273.n3 41.0422
R17 a_16273_n2273.n0 a_16273_n2273.t0 31.9797
R18 a_16620_n1869.n3 a_16620_n1869.n2 636.953
R19 a_16620_n1869.n1 a_16620_n1869.t4 366.856
R20 a_16620_n1869.n2 a_16620_n1869.n0 300.2
R21 a_16620_n1869.n2 a_16620_n1869.n1 225.036
R22 a_16620_n1869.n1 a_16620_n1869.t5 174.056
R23 a_16620_n1869.n0 a_16620_n1869.t2 70.0005
R24 a_16620_n1869.t0 a_16620_n1869.n3 68.0124
R25 a_16620_n1869.n3 a_16620_n1869.t1 63.3219
R26 a_16620_n1869.n0 a_16620_n1869.t3 61.6672
R27 dvss.n623 dvss.n622 844724
R28 dvss.n146 dvss.n145 148018
R29 dvss.n650 dvss.n17 121073
R30 dvss.n144 dvss.n44 20785.4
R31 dvss.n145 dvss.n144 13161.6
R32 dvss.n43 dvss.n42 10590.5
R33 dvss.n142 dvss.n40 8607.23
R34 dvss.n562 dvss.n546 8366.71
R35 dvss.n546 dvss.n92 8366.71
R36 dvss.n544 dvss.n92 8366.71
R37 dvss.n562 dvss.n544 8366.71
R38 dvss.n613 dvss.n612 5881.35
R39 dvss.n88 dvss.n40 5784.65
R40 dvss.n624 dvss.n31 5227.07
R41 dvss.n32 dvss.n31 5083.5
R42 dvss.n612 dvss.n44 4954.5
R43 dvss.n229 dvss.n227 4604.94
R44 dvss.n603 dvss.n44 4392.82
R45 dvss.n101 dvss.n93 4247.09
R46 dvss.n541 dvss.n93 4247.09
R47 dvss.n101 dvss.n94 4247.09
R48 dvss.n541 dvss.n94 4247.09
R49 dvss.n213 dvss.n206 4247.09
R50 dvss.n218 dvss.n206 4247.09
R51 dvss.n213 dvss.n207 4247.09
R52 dvss.n218 dvss.n207 4247.09
R53 dvss.n623 dvss.n32 3898.89
R54 dvss.n622 dvss.n621 3764.56
R55 dvss.n625 dvss.n624 3697.38
R56 dvss.n227 dvss.n90 3234.36
R57 dvss.n29 dvss.n15 2798.56
R58 dvss.n653 dvss.n15 2798.56
R59 dvss.n29 dvss.n16 2798.56
R60 dvss.n653 dvss.n16 2798.56
R61 dvss.n589 dvss.n55 2798.56
R62 dvss.n56 dvss.n55 2798.56
R63 dvss.n589 dvss.n60 2798.56
R64 dvss.n60 dvss.n56 2798.56
R65 dvss.n543 dvss.n542 2575.49
R66 dvss.n624 dvss.n623 2562.64
R67 dvss.n613 dvss.n43 2543.9
R68 dvss.n233 dvss.n83 2397.52
R69 dvss.n303 dvss.n302 2387.64
R70 dvss.n436 dvss.n146 2316.35
R71 dvss.n143 dvss.n142 2162.81
R72 dvss.n566 dvss.n90 2000.34
R73 dvss.n649 dvss.n18 1686.66
R74 dvss.n304 dvss.n303 1680.95
R75 dvss.n630 dvss.n626 1407.97
R76 dvss.n636 dvss.n626 1407.97
R77 dvss.n636 dvss.n627 1407.97
R78 dvss.n586 dvss.n62 1407.97
R79 dvss.n70 dvss.n62 1407.97
R80 dvss.n586 dvss.n63 1407.97
R81 dvss.n70 dvss.n63 1407.97
R82 dvss.n34 dvss.n32 1313.59
R83 dvss.n681 dvss.n0 1212.38
R84 dvss.n588 dvss.n61 1202.51
R85 dvss.n220 dvss.n7 1198.25
R86 dvss.n302 dvss.n301 1198.25
R87 dvss.n289 dvss.n235 1198.25
R88 dvss.n518 dvss.n109 1198.25
R89 dvss.n478 dvss.n126 1198.25
R90 dvss.n438 dvss.n437 1198.25
R91 dvss.n435 dvss.n434 1198.25
R92 dvss.n209 dvss.n164 1198.25
R93 dvss.n210 dvss.n181 1198.25
R94 dvss.n315 dvss.n200 1198.25
R95 dvss.n305 dvss.n304 1198.25
R96 dvss.n639 dvss.n638 1198.25
R97 dvss.n73 dvss.n72 1198.25
R98 dvss.n651 dvss.n650 1184.03
R99 dvss.n681 dvss.n680 1175.19
R100 dvss.n615 dvss.n35 1127.15
R101 dvss.n42 dvss.n41 1064.88
R102 dvss.t145 dvss.t96 935.78
R103 dvss.t98 dvss.t21 935.78
R104 dvss.t26 dvss.t100 935.78
R105 dvss.n574 dvss.n85 927.908
R106 dvss.n145 dvss.n49 900.194
R107 dvss.n620 dvss.n35 884.347
R108 dvss.n554 dvss.n553 784.03
R109 dvss.n561 dvss.n560 783.962
R110 dvss.n553 dvss.n552 783.75
R111 dvss.n561 dvss.n551 783.683
R112 dvss.n235 dvss.t19 748.625
R113 dvss.n614 dvss.n613 720.655
R114 dvss.t212 dvss.t151 717.851
R115 dvss.t11 dvss.t155 717.851
R116 dvss.t137 dvss.t112 689.909
R117 dvss.t112 dvss.t32 689.909
R118 dvss.t46 dvss.t118 689.909
R119 dvss.t118 dvss.t69 689.909
R120 dvss.t37 dvss.t168 689.909
R121 dvss.t9 dvss.t37 689.909
R122 dvss.n211 dvss.t135 655.918
R123 dvss.n652 dvss.n651 639.12
R124 dvss.n598 dvss.n597 626.816
R125 dvss.n30 dvss.t161 618.75
R126 dvss.n652 dvss.t161 618.75
R127 dvss.t131 dvss.t147 609.174
R128 dvss.t154 dvss.t182 609.174
R129 dvss.t176 dvss.t45 609.174
R130 dvss.n84 dvss.n81 585
R131 dvss.n84 dvss.n61 585
R132 dvss.n605 dvss.n604 585
R133 dvss.n604 dvss.n603 585
R134 dvss.n229 dvss.n107 585
R135 dvss.n229 dvss.n228 585
R136 dvss.n230 dvss.n83 585
R137 dvss.n91 dvss.n83 585
R138 dvss.n571 dvss.n570 585
R139 dvss.n572 dvss.n571 585
R140 dvss.n569 dvss.n88 585
R141 dvss.n88 dvss.n86 585
R142 dvss.t77 dvss.n200 574.28
R143 dvss.n437 dvss.t120 554.129
R144 dvss.n126 dvss.t73 554.129
R145 dvss.t1 dvss.n109 554.129
R146 dvss.t187 dvss.t70 546.789
R147 dvss.t149 dvss.t48 546.789
R148 dvss.t35 dvss.t129 546.789
R149 dvss.t28 dvss.t52 529.24
R150 dvss.t7 dvss.t28 529.24
R151 dvss.t81 dvss.t24 529.24
R152 dvss.t124 dvss.t81 529.24
R153 dvss.t56 dvss.t62 529.24
R154 dvss.t66 dvss.t56 529.24
R155 dvss.t39 dvss.t110 484.404
R156 dvss.t195 dvss.t200 484.404
R157 dvss.t3 dvss.t50 484.404
R158 dvss.t189 dvss.t0 467.307
R159 dvss.t17 dvss.t23 467.307
R160 dvss.t34 dvss.t90 467.307
R161 dvss.n615 dvss.n39 467.033
R162 dvss.t19 dvss.t143 447.707
R163 dvss.n303 dvss.n220 426.382
R164 dvss.n435 dvss.t209 425.08
R165 dvss.t198 dvss.n209 425.08
R166 dvss.t141 dvss.n210 425.08
R167 dvss.t132 dvss.t13 419.45
R168 dvss.t104 dvss.t93 419.45
R169 dvss.t60 dvss.t91 419.45
R170 dvss.n638 dvss.n637 419.18
R171 dvss.n597 dvss.n50 404.022
R172 dvss.t95 dvss.t44 400
R173 dvss.t103 dvss.t148 400
R174 dvss.t177 dvss.t194 400
R175 dvss.n630 dvss.n629 390.825
R176 dvss.t125 dvss.t5 371.594
R177 dvss.t64 dvss.t205 371.594
R178 dvss.t165 dvss.t139 371.594
R179 dvss.n651 dvss.t41 366.435
R180 dvss.t44 dvss.t39 363.303
R181 dvss.t148 dvss.t195 363.303
R182 dvss.t50 dvss.t177 363.303
R183 dvss.t120 dvss.t137 355.964
R184 dvss.t73 dvss.t46 355.964
R185 dvss.t168 dvss.t1 355.964
R186 dvss.t70 dvss.t95 352.295
R187 dvss.t147 dvss.t211 352.295
R188 dvss.t48 dvss.t103 352.295
R189 dvss.t182 dvss.t204 352.295
R190 dvss.t194 dvss.t35 352.295
R191 dvss.t211 dvss.t145 348.625
R192 dvss.t204 dvss.t98 348.625
R193 dvss.t18 dvss.t26 348.625
R194 dvss.n637 dvss.n625 344.228
R195 dvss.t122 dvss.t77 343.442
R196 dvss.n233 dvss.n229 335.039
R197 dvss.t32 dvss.t187 333.945
R198 dvss.t69 dvss.t149 333.945
R199 dvss.t129 dvss.t9 333.945
R200 dvss.n85 dvss.n84 331.606
R201 dvss.n228 dvss.t18 326.606
R202 dvss.n615 dvss.n40 310.599
R203 dvss.n41 dvss.n35 308.933
R204 dvss.n437 dvss.n436 308.257
R205 dvss.t96 dvss.t178 308.257
R206 dvss.t21 dvss.t88 308.257
R207 dvss.n638 dvss 308.139
R208 dvss.n283 dvss.t27 307.536
R209 dvss.n512 dvss.t99 307.536
R210 dvss.n472 dvss.t146 307.536
R211 dvss.n161 dvss.t152 307.536
R212 dvss.n178 dvss.t156 307.536
R213 dvss.n321 dvss.t80 307.536
R214 dvss.t8 dvss.t10 306.846
R215 dvss.t72 dvss.t87 306.846
R216 dvss.t167 dvss.t43 306.846
R217 dvss.n70 dvss.n69 292.5
R218 dvss.n71 dvss.n70 292.5
R219 dvss.n68 dvss.n63 292.5
R220 dvss.t108 dvss.n63 292.5
R221 dvss.n586 dvss.n585 292.5
R222 dvss.n587 dvss.n586 292.5
R223 dvss.n64 dvss.n62 292.5
R224 dvss.t108 dvss.n62 292.5
R225 dvss.n633 dvss.n627 292.5
R226 dvss.n636 dvss.n635 292.5
R227 dvss.n637 dvss.n636 292.5
R228 dvss.n628 dvss.n626 292.5
R229 dvss.t190 dvss.n626 292.5
R230 dvss.n631 dvss.n630 292.5
R231 dvss.t171 dvss 289.909
R232 dvss.t5 dvss.t8 278.695
R233 dvss.t205 dvss.t72 278.695
R234 dvss.t139 dvss.t167 278.695
R235 dvss.n217 dvss.n215 276.286
R236 dvss dvss.n126 275.229
R237 dvss dvss.n109 275.229
R238 dvss.n235 dvss 275.229
R239 dvss.n302 dvss 275.229
R240 dvss.t202 dvss.n0 273.678
R241 dvss.n542 dvss.t202 273.678
R242 dvss.t52 dvss.t209 273.065
R243 dvss.t24 dvss.t198 273.065
R244 dvss.t62 dvss.t141 273.065
R245 dvss.t10 dvss.t132 270.25
R246 dvss.t214 dvss.t189 270.25
R247 dvss.t87 dvss.t104 270.25
R248 dvss.t58 dvss.t17 270.25
R249 dvss.t43 dvss.t60 270.25
R250 dvss.t151 dvss.t214 267.435
R251 dvss.t155 dvss.t58 267.435
R252 dvss.t134 dvss.t79 267.435
R253 dvss.t110 dvss.t131 264.221
R254 dvss.t200 dvss.t154 264.221
R255 dvss.t45 dvss.t3 264.221
R256 dvss.t143 dvss.t171 264.221
R257 dvss.n611 dvss.n45 258.5
R258 dvss.t13 dvss.t7 256.175
R259 dvss.t93 dvss.t124 256.175
R260 dvss.t91 dvss.t66 256.175
R261 dvss.n543 dvss.t174 255.168
R262 dvss.n256 dvss.t38 246.817
R263 dvss.n485 dvss.t119 246.817
R264 dvss.n445 dvss.t113 246.817
R265 dvss.n151 dvss.t29 246.817
R266 dvss.n386 dvss.t82 246.817
R267 dvss.n347 dvss.t57 246.817
R268 dvss.t191 dvss.t41 244.291
R269 dvss.t178 dvss 238.532
R270 dvss.t88 dvss 238.532
R271 dvss dvss.t207 238.532
R272 dvss.n436 dvss.n435 236.469
R273 dvss.t67 dvss.t212 236.469
R274 dvss.t54 dvss.t11 236.469
R275 dvss.t135 dvss.t180 236.469
R276 dvss.n61 dvss.n42 236.023
R277 dvss.n588 dvss.n587 230.855
R278 dvss.n325 dvss.t86 229.185
R279 dvss.n522 dvss.n521 227.357
R280 dvss.n97 dvss.t203 219.8
R281 dvss.n540 dvss.n95 217.329
R282 dvss.n215 dvss.n214 217.225
R283 dvss.n249 dvss.n248 214.742
R284 dvss.n123 dvss.n122 214.742
R285 dvss.n140 dvss.n139 214.742
R286 dvss.n150 dvss.n149 214.742
R287 dvss.n392 dvss.n166 214.742
R288 dvss.n353 dvss.n183 214.742
R289 dvss.n571 dvss.n87 213.325
R290 dvss.n209 dvss 211.132
R291 dvss.n210 dvss 211.132
R292 dvss dvss.n200 211.132
R293 dvss.n304 dvss 211.132
R294 dvss.n263 dvss.n245 209.254
R295 dvss.n492 dvss.n119 209.254
R296 dvss.n452 dvss.n136 209.254
R297 dvss.n154 dvss.n153 209.254
R298 dvss.n172 dvss.n171 209.254
R299 dvss.n189 dvss.n188 209.254
R300 dvss.t174 dvss.t185 208.894
R301 dvss.t185 dvss.t159 208.894
R302 dvss.t159 dvss.t15 208.894
R303 dvss.t15 dvss.t127 208.894
R304 dvss.t75 dvss.t163 208.894
R305 dvss.t163 dvss.t172 208.894
R306 dvss.t183 dvss.t157 208.894
R307 dvss.n526 dvss.n525 203.619
R308 dvss.t0 dvss.t125 202.688
R309 dvss.t23 dvss.t64 202.688
R310 dvss.t90 dvss.t165 202.688
R311 dvss.t102 dvss.t122 202.688
R312 dvss.n666 dvss.n6 202.067
R313 dvss.n604 dvss.n45 202.048
R314 dvss.n3 dvss.n2 200.516
R315 dvss.n237 dvss.n236 199.739
R316 dvss.n271 dvss.n270 199.739
R317 dvss.n111 dvss.n110 199.739
R318 dvss.n500 dvss.n499 199.739
R319 dvss.n128 dvss.n127 199.739
R320 dvss.n460 dvss.n459 199.739
R321 dvss.n412 dvss.n158 199.739
R322 dvss.n399 dvss.n163 199.739
R323 dvss.n373 dvss.n175 199.739
R324 dvss.n360 dvss.n180 199.739
R325 dvss.n334 dvss.n192 199.739
R326 dvss.n199 dvss.n198 199.739
R327 dvss.n24 dvss.n23 199.739
R328 dvss.n75 dvss.n74 199.739
R329 dvss.n540 dvss.n539 198.024
R330 dvss.n587 dvss.t30 187.785
R331 dvss.n295 dvss.n294 185
R332 dvss.n205 dvss.n204 185
R333 dvss.n679 dvss.n678 185
R334 dvss dvss.t67 182.982
R335 dvss dvss.t54 182.982
R336 dvss.n28 dvss.n12 181.835
R337 dvss.n28 dvss.n27 181.835
R338 dvss.n58 dvss.n57 181.835
R339 dvss.n59 dvss.n58 181.835
R340 dvss.n629 dvss.n627 174.962
R341 dvss.n212 dvss.t134 166.091
R342 dvss.n234 dvss.t100 161.469
R343 dvss.n31 dvss.n30 155.325
R344 dvss.n219 dvss.t102 154.831
R345 dvss.n95 dvss.n93 148.029
R346 dvss.t207 dvss.n234 146.79
R347 dvss.n218 dvss.n217 146.25
R348 dvss.n219 dvss.n218 146.25
R349 dvss.n214 dvss.n213 146.25
R350 dvss.n213 dvss.n212 146.25
R351 dvss.n96 dvss.n94 146.25
R352 dvss.n94 dvss.t202 146.25
R353 dvss.n93 dvss.t202 146.25
R354 dvss.n102 dvss.n95 143.809
R355 dvss.n577 dvss.n81 143.196
R356 dvss.t106 dvss 141.269
R357 dvss.t180 dvss.t85 140.756
R358 dvss dvss.t83 140.144
R359 dvss.n545 dvss.n86 129.567
R360 dvss.n574 dvss.n83 128.583
R361 dvss.n217 dvss.n216 127.487
R362 dvss.n72 dvss.n33 122.319
R363 dvss.t157 dvss.n572 120.312
R364 dvss.n58 dvss.n56 117.001
R365 dvss.n56 dvss.n33 117.001
R366 dvss.n60 dvss.n59 117.001
R367 dvss.t30 dvss.n60 117.001
R368 dvss.n590 dvss.n589 117.001
R369 dvss.n589 dvss.n588 117.001
R370 dvss.n57 dvss.n55 117.001
R371 dvss.t30 dvss.n55 117.001
R372 dvss.n654 dvss.n653 117.001
R373 dvss.n653 dvss.n652 117.001
R374 dvss.n16 dvss.n12 117.001
R375 dvss.t161 dvss.n16 117.001
R376 dvss.n29 dvss.n28 117.001
R377 dvss.n30 dvss.n29 117.001
R378 dvss.n27 dvss.n15 117.001
R379 dvss.t161 dvss.n15 117.001
R380 dvss.n573 dvss.t172 113.703
R381 dvss.n232 dvss.n231 108.201
R382 dvss.n622 dvss.n33 105.091
R383 dvss.n212 dvss.t34 104.159
R384 dvss.n654 dvss.n13 102.025
R385 dvss.n655 dvss.n654 102.025
R386 dvss.n590 dvss.n52 102.025
R387 dvss.n590 dvss.n54 102.025
R388 dvss.n648 dvss.n19 101.874
R389 dvss.t127 dvss.n91 101.803
R390 dvss.n245 dvss.t130 100.001
R391 dvss.n119 dvss.t150 100.001
R392 dvss.n136 dvss.t188 100.001
R393 dvss.n153 dvss.t14 100.001
R394 dvss.n171 dvss.t94 100.001
R395 dvss.n188 dvss.t92 100.001
R396 dvss.n599 dvss.n598 98.4337
R397 dvss.n573 dvss.t183 95.1928
R398 dvss.n631 dvss.n628 91.4829
R399 dvss.n69 dvss.n64 91.4829
R400 dvss.n545 dvss.n43 85.938
R401 dvss.n53 dvss.t31 83.7183
R402 dvss.n646 dvss.t162 83.7183
R403 dvss.n142 dvss.n45 81.509
R404 dvss.n629 dvss.t190 81.1932
R405 dvss dvss.t191 80.5052
R406 dvss.n655 dvss.n12 79.8123
R407 dvss.n27 dvss.n13 79.8123
R408 dvss.n59 dvss.n52 79.8123
R409 dvss.n57 dvss.n54 79.8123
R410 dvss.n617 dvss.n616 73.2369
R411 dvss.n616 dvss.n615 73.1255
R412 dvss.n615 dvss.n614 73.1255
R413 dvss.n294 dvss.t20 72.8576
R414 dvss.n270 dvss.t4 72.8576
R415 dvss.n499 dvss.t201 72.8576
R416 dvss.n459 dvss.t111 72.8576
R417 dvss.n204 dvss.t78 72.8576
R418 dvss.n158 dvss.t126 72.8576
R419 dvss.n175 dvss.t65 72.8576
R420 dvss.n192 dvss.t166 72.8576
R421 dvss.n41 dvss.n39 72.01
R422 dvss.n521 dvss.n107 71.4371
R423 dvss.n245 dvss.t36 70.0005
R424 dvss.n119 dvss.t49 70.0005
R425 dvss.n136 dvss.t71 70.0005
R426 dvss.n153 dvss.t133 70.0005
R427 dvss.n171 dvss.t105 70.0005
R428 dvss.n188 dvss.t61 70.0005
R429 dvss.n69 dvss.n68 69.6045
R430 dvss.n635 dvss.n628 69.0306
R431 dvss dvss.t108 68.912
R432 dvss.n208 dvss.n196 68.8106
R433 dvss dvss.n219 67.5629
R434 dvss.n585 dvss.n64 66.3131
R435 dvss.n632 dvss.n631 65.475
R436 dvss.n527 dvss.n526 64.5768
R437 dvss.n564 dvss.t75 63.462
R438 dvss.t79 dvss.n211 61.9327
R439 dvss.n270 dvss.t51 60.5809
R440 dvss.n499 dvss.t196 60.5809
R441 dvss.n459 dvss.t40 60.5809
R442 dvss.n158 dvss.t6 60.5809
R443 dvss.n175 dvss.t206 60.5809
R444 dvss.n192 dvss.t140 60.5809
R445 dvss.n294 dvss.t144 58.5719
R446 dvss.n204 dvss.t123 58.5719
R447 dvss.n619 dvss.n617 57.4606
R448 dvss.n599 dvss.n49 57.2559
R449 dvss.n248 dvss.t169 57.1434
R450 dvss.n122 dvss.t47 57.1434
R451 dvss.n139 dvss.t138 57.1434
R452 dvss.n149 dvss.t53 57.1434
R453 dvss.n166 dvss.t25 57.1434
R454 dvss.n183 dvss.t63 57.1434
R455 dvss.n614 dvss.n42 54.0496
R456 dvss.n678 dvss.t117 52.8576
R457 dvss.n678 dvss.t84 51.4291
R458 dvss.n576 dvss.n575 45.2502
R459 dvss.n85 dvss.n39 44.978
R460 dvss.t85 dvss 42.227
R461 dvss.n216 dvss.n207 41.7862
R462 dvss.t85 dvss.n207 41.7862
R463 dvss.n215 dvss.n206 41.7862
R464 dvss.t85 dvss.n206 41.7862
R465 dvss.n541 dvss.n540 41.7862
R466 dvss.n542 dvss.n541 41.7862
R467 dvss.n102 dvss.n101 41.7862
R468 dvss.n101 dvss.n0 41.7862
R469 dvss.n554 dvss.n546 41.7862
R470 dvss.n546 dvss.n545 41.7862
R471 dvss.n552 dvss.n544 41.7862
R472 dvss.n544 dvss.n543 41.7862
R473 dvss.n231 dvss.n230 40.2432
R474 dvss.n677 dvss.n676 40.0735
R475 dvss.n236 dvss.t101 38.5719
R476 dvss.n236 dvss.t208 38.5719
R477 dvss.n110 dvss.t22 38.5719
R478 dvss.n110 dvss.t89 38.5719
R479 dvss.n127 dvss.t97 38.5719
R480 dvss.n127 dvss.t179 38.5719
R481 dvss.n163 dvss.t213 38.5719
R482 dvss.n163 dvss.t68 38.5719
R483 dvss.n180 dvss.t12 38.5719
R484 dvss.n180 dvss.t55 38.5719
R485 dvss.n198 dvss.t136 38.5719
R486 dvss.n198 dvss.t181 38.5719
R487 dvss.n634 dvss.n633 37.6894
R488 dvss.n584 dvss.n65 37.4862
R489 dvss.n611 dvss.n40 36.1883
R490 dvss.t108 dvss.t30 36.179
R491 dvss.n72 dvss.n71 36.179
R492 dvss.n6 dvss.t193 36.0005
R493 dvss.n565 dvss.n563 35.6976
R494 dvss.n537 dvss.n536 35.5421
R495 dvss.n670 dvss.n5 34.6358
R496 dvss.n671 dvss.n670 34.6358
R497 dvss.n672 dvss.n671 34.6358
R498 dvss.n300 dvss.n225 34.6358
R499 dvss.n293 dvss.n226 34.6358
R500 dvss.n276 dvss.n241 34.6358
R501 dvss.n277 dvss.n276 34.6358
R502 dvss.n278 dvss.n277 34.6358
R503 dvss.n278 dvss.n239 34.6358
R504 dvss.n282 dvss.n239 34.6358
R505 dvss.n264 dvss.n243 34.6358
R506 dvss.n268 dvss.n243 34.6358
R507 dvss.n269 dvss.n268 34.6358
R508 dvss.n272 dvss.n269 34.6358
R509 dvss.n251 dvss.n108 34.6358
R510 dvss.n255 dvss.n254 34.6358
R511 dvss.n257 dvss.n255 34.6358
R512 dvss.n261 dvss.n246 34.6358
R513 dvss.n262 dvss.n261 34.6358
R514 dvss.n505 dvss.n115 34.6358
R515 dvss.n506 dvss.n505 34.6358
R516 dvss.n507 dvss.n506 34.6358
R517 dvss.n507 dvss.n113 34.6358
R518 dvss.n511 dvss.n113 34.6358
R519 dvss.n493 dvss.n117 34.6358
R520 dvss.n497 dvss.n117 34.6358
R521 dvss.n498 dvss.n497 34.6358
R522 dvss.n501 dvss.n498 34.6358
R523 dvss.n480 dvss.n479 34.6358
R524 dvss.n484 dvss.n483 34.6358
R525 dvss.n486 dvss.n484 34.6358
R526 dvss.n490 dvss.n120 34.6358
R527 dvss.n491 dvss.n490 34.6358
R528 dvss.n465 dvss.n132 34.6358
R529 dvss.n466 dvss.n465 34.6358
R530 dvss.n467 dvss.n466 34.6358
R531 dvss.n467 dvss.n130 34.6358
R532 dvss.n471 dvss.n130 34.6358
R533 dvss.n453 dvss.n134 34.6358
R534 dvss.n457 dvss.n134 34.6358
R535 dvss.n458 dvss.n457 34.6358
R536 dvss.n461 dvss.n458 34.6358
R537 dvss.n440 dvss.n439 34.6358
R538 dvss.n444 dvss.n443 34.6358
R539 dvss.n446 dvss.n444 34.6358
R540 dvss.n450 dvss.n137 34.6358
R541 dvss.n451 dvss.n450 34.6358
R542 dvss.n433 dvss.n147 34.6358
R543 dvss.n429 dvss.n428 34.6358
R544 dvss.n428 dvss.n427 34.6358
R545 dvss.n424 dvss.n423 34.6358
R546 dvss.n423 dvss.n422 34.6358
R547 dvss.n419 dvss.n418 34.6358
R548 dvss.n418 dvss.n417 34.6358
R549 dvss.n417 dvss.n156 34.6358
R550 dvss.n413 dvss.n156 34.6358
R551 dvss.n411 dvss.n410 34.6358
R552 dvss.n410 dvss.n159 34.6358
R553 dvss.n406 dvss.n159 34.6358
R554 dvss.n406 dvss.n405 34.6358
R555 dvss.n405 dvss.n404 34.6358
R556 dvss.n394 dvss.n393 34.6358
R557 dvss.n391 dvss.n167 34.6358
R558 dvss.n387 dvss.n167 34.6358
R559 dvss.n385 dvss.n384 34.6358
R560 dvss.n384 dvss.n169 34.6358
R561 dvss.n380 dvss.n379 34.6358
R562 dvss.n379 dvss.n378 34.6358
R563 dvss.n378 dvss.n173 34.6358
R564 dvss.n374 dvss.n173 34.6358
R565 dvss.n372 dvss.n371 34.6358
R566 dvss.n371 dvss.n176 34.6358
R567 dvss.n367 dvss.n176 34.6358
R568 dvss.n367 dvss.n366 34.6358
R569 dvss.n366 dvss.n365 34.6358
R570 dvss.n355 dvss.n354 34.6358
R571 dvss.n352 dvss.n184 34.6358
R572 dvss.n348 dvss.n184 34.6358
R573 dvss.n346 dvss.n345 34.6358
R574 dvss.n345 dvss.n186 34.6358
R575 dvss.n341 dvss.n340 34.6358
R576 dvss.n340 dvss.n190 34.6358
R577 dvss.n336 dvss.n190 34.6358
R578 dvss.n336 dvss.n335 34.6358
R579 dvss.n333 dvss.n193 34.6358
R580 dvss.n329 dvss.n193 34.6358
R581 dvss.n329 dvss.n328 34.6358
R582 dvss.n328 dvss.n195 34.6358
R583 dvss.n322 dvss.n195 34.6358
R584 dvss.n314 dvss.n202 34.6358
R585 dvss.n309 dvss.n308 34.6358
R586 dvss.n23 dvss.t192 33.462
R587 dvss.n23 dvss.t42 33.462
R588 dvss.n74 dvss.t109 33.462
R589 dvss.n74 dvss.t107 33.462
R590 dvss.n2 dvss.t197 33.2313
R591 dvss.n24 dvss.n21 31.5123
R592 dvss.n254 dvss.n249 31.2476
R593 dvss.n483 dvss.n123 31.2476
R594 dvss.n443 dvss.n140 31.2476
R595 dvss.n429 dvss.n150 31.2476
R596 dvss.n392 dvss.n391 31.2476
R597 dvss.n353 dvss.n352 31.2476
R598 dvss.t33 dvss.t83 30.4092
R599 dvss dvss.n681 30.4092
R600 dvss.n616 dvss.n37 30.2484
R601 dvss.n284 dvss.n283 29.7417
R602 dvss.n513 dvss.n512 29.7417
R603 dvss.n473 dvss.n472 29.7417
R604 dvss.n400 dvss.n161 29.7417
R605 dvss.n361 dvss.n178 29.7417
R606 dvss.n321 dvss.n320 29.7417
R607 dvss.n80 dvss.n37 28.5338
R608 dvss.n538 dvss.n99 28.3255
R609 dvss.n527 dvss.n100 27.9866
R610 dvss.n256 dvss.n246 27.8593
R611 dvss.n485 dvss.n120 27.8593
R612 dvss.n445 dvss.n137 27.8593
R613 dvss.n424 dvss.n151 27.8593
R614 dvss.n386 dvss.n385 27.8593
R615 dvss.n347 dvss.n346 27.8593
R616 dvss.n676 dvss.n3 25.977
R617 dvss.n228 dvss.t176 25.6886
R618 dvss.n248 dvss.t2 25.4291
R619 dvss.n122 dvss.t74 25.4291
R620 dvss.n139 dvss.t121 25.4291
R621 dvss.n149 dvss.t210 25.4291
R622 dvss.n166 dvss.t199 25.4291
R623 dvss.n183 dvss.t142 25.4291
R624 dvss.n2 dvss.t153 24.9236
R625 dvss.n6 dvss.t59 24.9236
R626 dvss.n562 dvss.n561 24.3755
R627 dvss.n563 dvss.n562 24.3755
R628 dvss.n553 dvss.n92 24.3755
R629 dvss.n563 dvss.n92 24.3755
R630 dvss.n296 dvss.n225 23.7737
R631 dvss.n310 dvss.n309 23.7737
R632 dvss.n665 dvss.n7 23.7181
R633 dvss.n301 dvss.n300 23.7181
R634 dvss.n289 dvss.n226 23.7181
R635 dvss.n289 dvss.n288 23.7181
R636 dvss.n518 dvss.n108 23.7181
R637 dvss.n518 dvss.n517 23.7181
R638 dvss.n479 dvss.n478 23.7181
R639 dvss.n478 dvss.n477 23.7181
R640 dvss.n439 dvss.n438 23.7181
R641 dvss.n434 dvss.n433 23.7181
R642 dvss.n398 dvss.n164 23.7181
R643 dvss.n394 dvss.n164 23.7181
R644 dvss.n359 dvss.n181 23.7181
R645 dvss.n355 dvss.n181 23.7181
R646 dvss.n316 dvss.n315 23.7181
R647 dvss.n315 dvss.n314 23.7181
R648 dvss.n308 dvss.n305 23.7181
R649 dvss.n639 dvss.n26 23.7181
R650 dvss.n76 dvss.n73 23.7181
R651 dvss.n666 dvss.n5 22.9652
R652 dvss.n284 dvss.n237 22.9652
R653 dvss.n513 dvss.n111 22.9652
R654 dvss.n473 dvss.n128 22.9652
R655 dvss.n400 dvss.n399 22.9652
R656 dvss.n361 dvss.n360 22.9652
R657 dvss.n320 dvss.n199 22.9652
R658 dvss.n537 dvss.n533 22.1054
R659 dvss.n232 dvss.n107 21.7695
R660 dvss.n98 dvss.n97 21.753
R661 dvss.n666 dvss.n665 21.4593
R662 dvss.n288 dvss.n237 21.4593
R663 dvss.n517 dvss.n111 21.4593
R664 dvss.n477 dvss.n128 21.4593
R665 dvss.n399 dvss.n398 21.4593
R666 dvss.n360 dvss.n359 21.4593
R667 dvss.n316 dvss.n199 21.4593
R668 dvss.n680 dvss.n679 21.4265
R669 dvss.n552 dvss.t175 21.1687
R670 dvss.n554 dvss.t158 21.1687
R671 dvss.n220 dvss.t33 21.1543
R672 dvss.n295 dvss.n293 20.9718
R673 dvss.n205 dvss.n202 20.9718
R674 dvss.n576 dvss.n37 20.1009
R675 dvss.n617 dvss.n36 20.0732
R676 dvss.n528 dvss.n527 18.7867
R677 dvss.n559 dvss.n555 18.4515
R678 dvss.n558 dvss.n556 18.4515
R679 dvss.n549 dvss.n548 18.4515
R680 dvss.n550 dvss.n547 18.4515
R681 dvss.n672 dvss.n3 18.4476
R682 dvss.n263 dvss.n262 17.6946
R683 dvss.n492 dvss.n491 17.6946
R684 dvss.n452 dvss.n451 17.6946
R685 dvss.n422 dvss.n154 17.6946
R686 dvss.n172 dvss.n169 17.6946
R687 dvss.n189 dvss.n186 17.6946
R688 dvss.t190 dvss.n625 16.6567
R689 dvss dvss.n24 15.0593
R690 dvss dvss.n75 15.0593
R691 dvss.n283 dvss.n282 14.6829
R692 dvss.n512 dvss.n511 14.6829
R693 dvss.n472 dvss.n471 14.6829
R694 dvss.n404 dvss.n161 14.6829
R695 dvss.n365 dvss.n178 14.6829
R696 dvss.n322 dvss.n321 14.6829
R697 dvss.n594 dvss.n593 14.3573
R698 dvss.n570 dvss.n568 13.8612
R699 dvss.n71 dvss.t106 13.7828
R700 dvss.n99 dvss.n98 13.2836
R701 dvss.n606 dvss.n47 13.0628
R702 dvss.n610 dvss.n609 12.2414
R703 dvss.n97 dvss.n95 11.7338
R704 dvss.n581 dvss.n54 10.5081
R705 dvss.n597 dvss.n596 10.2484
R706 dvss.n592 dvss.n52 10.2179
R707 dvss.n656 dvss.n655 10.1264
R708 dvss.n649 dvss.n648 9.79535
R709 dvss.n582 dvss.n79 9.76662
R710 dvss.n596 dvss.n38 9.49353
R711 dvss.n80 dvss.n79 9.30109
R712 dvss.n306 dvss.n305 9.3005
R713 dvss.n324 dvss.n195 9.3005
R714 dvss.n323 dvss.n322 9.3005
R715 dvss.n321 dvss.n197 9.3005
R716 dvss.n320 dvss.n319 9.3005
R717 dvss.n318 dvss.n199 9.3005
R718 dvss.n317 dvss.n316 9.3005
R719 dvss.n315 dvss.n201 9.3005
R720 dvss.n314 dvss.n313 9.3005
R721 dvss.n312 dvss.n202 9.3005
R722 dvss.n311 dvss.n310 9.3005
R723 dvss.n309 dvss.n203 9.3005
R724 dvss.n308 dvss.n307 9.3005
R725 dvss.n434 dvss.n105 9.3005
R726 dvss.n433 dvss.n432 9.3005
R727 dvss.n431 dvss.n147 9.3005
R728 dvss.n430 dvss.n429 9.3005
R729 dvss.n428 dvss.n148 9.3005
R730 dvss.n427 dvss.n426 9.3005
R731 dvss.n425 dvss.n424 9.3005
R732 dvss.n423 dvss.n152 9.3005
R733 dvss.n422 dvss.n421 9.3005
R734 dvss.n420 dvss.n419 9.3005
R735 dvss.n418 dvss.n155 9.3005
R736 dvss.n417 dvss.n416 9.3005
R737 dvss.n415 dvss.n156 9.3005
R738 dvss.n414 dvss.n413 9.3005
R739 dvss.n411 dvss.n157 9.3005
R740 dvss.n410 dvss.n409 9.3005
R741 dvss.n408 dvss.n159 9.3005
R742 dvss.n407 dvss.n406 9.3005
R743 dvss.n405 dvss.n160 9.3005
R744 dvss.n404 dvss.n403 9.3005
R745 dvss.n402 dvss.n161 9.3005
R746 dvss.n401 dvss.n400 9.3005
R747 dvss.n399 dvss.n162 9.3005
R748 dvss.n398 dvss.n397 9.3005
R749 dvss.n396 dvss.n164 9.3005
R750 dvss.n395 dvss.n394 9.3005
R751 dvss.n393 dvss.n165 9.3005
R752 dvss.n391 dvss.n390 9.3005
R753 dvss.n389 dvss.n167 9.3005
R754 dvss.n388 dvss.n387 9.3005
R755 dvss.n385 dvss.n168 9.3005
R756 dvss.n384 dvss.n383 9.3005
R757 dvss.n382 dvss.n169 9.3005
R758 dvss.n381 dvss.n380 9.3005
R759 dvss.n379 dvss.n170 9.3005
R760 dvss.n378 dvss.n377 9.3005
R761 dvss.n376 dvss.n173 9.3005
R762 dvss.n375 dvss.n374 9.3005
R763 dvss.n372 dvss.n174 9.3005
R764 dvss.n371 dvss.n370 9.3005
R765 dvss.n369 dvss.n176 9.3005
R766 dvss.n368 dvss.n367 9.3005
R767 dvss.n366 dvss.n177 9.3005
R768 dvss.n365 dvss.n364 9.3005
R769 dvss.n363 dvss.n178 9.3005
R770 dvss.n362 dvss.n361 9.3005
R771 dvss.n360 dvss.n179 9.3005
R772 dvss.n359 dvss.n358 9.3005
R773 dvss.n357 dvss.n181 9.3005
R774 dvss.n356 dvss.n355 9.3005
R775 dvss.n354 dvss.n182 9.3005
R776 dvss.n352 dvss.n351 9.3005
R777 dvss.n350 dvss.n184 9.3005
R778 dvss.n349 dvss.n348 9.3005
R779 dvss.n346 dvss.n185 9.3005
R780 dvss.n345 dvss.n344 9.3005
R781 dvss.n343 dvss.n186 9.3005
R782 dvss.n342 dvss.n341 9.3005
R783 dvss.n340 dvss.n339 9.3005
R784 dvss.n338 dvss.n190 9.3005
R785 dvss.n337 dvss.n336 9.3005
R786 dvss.n335 dvss.n191 9.3005
R787 dvss.n333 dvss.n332 9.3005
R788 dvss.n331 dvss.n193 9.3005
R789 dvss.n330 dvss.n329 9.3005
R790 dvss.n328 dvss.n327 9.3005
R791 dvss.n438 dvss.n106 9.3005
R792 dvss.n439 dvss.n141 9.3005
R793 dvss.n441 dvss.n440 9.3005
R794 dvss.n443 dvss.n442 9.3005
R795 dvss.n444 dvss.n138 9.3005
R796 dvss.n447 dvss.n446 9.3005
R797 dvss.n448 dvss.n137 9.3005
R798 dvss.n450 dvss.n449 9.3005
R799 dvss.n451 dvss.n135 9.3005
R800 dvss.n454 dvss.n453 9.3005
R801 dvss.n455 dvss.n134 9.3005
R802 dvss.n457 dvss.n456 9.3005
R803 dvss.n458 dvss.n133 9.3005
R804 dvss.n462 dvss.n461 9.3005
R805 dvss.n463 dvss.n132 9.3005
R806 dvss.n465 dvss.n464 9.3005
R807 dvss.n466 dvss.n131 9.3005
R808 dvss.n468 dvss.n467 9.3005
R809 dvss.n469 dvss.n130 9.3005
R810 dvss.n471 dvss.n470 9.3005
R811 dvss.n472 dvss.n129 9.3005
R812 dvss.n474 dvss.n473 9.3005
R813 dvss.n475 dvss.n128 9.3005
R814 dvss.n477 dvss.n476 9.3005
R815 dvss.n478 dvss.n125 9.3005
R816 dvss.n479 dvss.n124 9.3005
R817 dvss.n481 dvss.n480 9.3005
R818 dvss.n483 dvss.n482 9.3005
R819 dvss.n484 dvss.n121 9.3005
R820 dvss.n487 dvss.n486 9.3005
R821 dvss.n488 dvss.n120 9.3005
R822 dvss.n490 dvss.n489 9.3005
R823 dvss.n491 dvss.n118 9.3005
R824 dvss.n494 dvss.n493 9.3005
R825 dvss.n495 dvss.n117 9.3005
R826 dvss.n497 dvss.n496 9.3005
R827 dvss.n498 dvss.n116 9.3005
R828 dvss.n502 dvss.n501 9.3005
R829 dvss.n503 dvss.n115 9.3005
R830 dvss.n505 dvss.n504 9.3005
R831 dvss.n506 dvss.n114 9.3005
R832 dvss.n508 dvss.n507 9.3005
R833 dvss.n509 dvss.n113 9.3005
R834 dvss.n511 dvss.n510 9.3005
R835 dvss.n512 dvss.n112 9.3005
R836 dvss.n514 dvss.n513 9.3005
R837 dvss.n515 dvss.n111 9.3005
R838 dvss.n517 dvss.n516 9.3005
R839 dvss.n519 dvss.n518 9.3005
R840 dvss.n250 dvss.n108 9.3005
R841 dvss.n252 dvss.n251 9.3005
R842 dvss.n254 dvss.n253 9.3005
R843 dvss.n255 dvss.n247 9.3005
R844 dvss.n258 dvss.n257 9.3005
R845 dvss.n259 dvss.n246 9.3005
R846 dvss.n261 dvss.n260 9.3005
R847 dvss.n262 dvss.n244 9.3005
R848 dvss.n265 dvss.n264 9.3005
R849 dvss.n266 dvss.n243 9.3005
R850 dvss.n268 dvss.n267 9.3005
R851 dvss.n269 dvss.n242 9.3005
R852 dvss.n273 dvss.n272 9.3005
R853 dvss.n274 dvss.n241 9.3005
R854 dvss.n276 dvss.n275 9.3005
R855 dvss.n277 dvss.n240 9.3005
R856 dvss.n279 dvss.n278 9.3005
R857 dvss.n280 dvss.n239 9.3005
R858 dvss.n282 dvss.n281 9.3005
R859 dvss.n283 dvss.n238 9.3005
R860 dvss.n285 dvss.n284 9.3005
R861 dvss.n286 dvss.n237 9.3005
R862 dvss.n288 dvss.n287 9.3005
R863 dvss.n290 dvss.n289 9.3005
R864 dvss.n291 dvss.n226 9.3005
R865 dvss.n293 dvss.n292 9.3005
R866 dvss.n297 dvss.n296 9.3005
R867 dvss.n298 dvss.n225 9.3005
R868 dvss.n300 dvss.n299 9.3005
R869 dvss.n301 dvss.n224 9.3005
R870 dvss.n662 dvss.n7 9.3005
R871 dvss.n667 dvss.n666 9.3005
R872 dvss.n673 dvss.n672 9.3005
R873 dvss.n671 dvss.n4 9.3005
R874 dvss.n670 dvss.n669 9.3005
R875 dvss.n668 dvss.n5 9.3005
R876 dvss.n665 dvss.n664 9.3005
R877 dvss.n674 dvss.n3 9.3005
R878 dvss.n676 dvss.n675 9.3005
R879 dvss.n640 dvss.n639 9.3005
R880 dvss.n24 dvss.n20 9.3005
R881 dvss.n26 dvss.n25 9.3005
R882 dvss.n644 dvss.n13 9.3005
R883 dvss.n77 dvss.n76 9.3005
R884 dvss.n73 dvss.n67 9.3005
R885 dvss.n635 dvss.n634 8.88939
R886 dvss.n68 dvss.n65 8.77764
R887 dvss.n528 dvss.n103 8.43597
R888 dvss.n271 dvss.n241 7.90638
R889 dvss.n500 dvss.n115 7.90638
R890 dvss.n460 dvss.n132 7.90638
R891 dvss.n412 dvss.n411 7.90638
R892 dvss.n373 dvss.n372 7.90638
R893 dvss.n334 dvss.n333 7.90638
R894 dvss.n620 dvss.n619 7.40556
R895 dvss.n621 dvss.n620 7.40556
R896 dvss.n603 dvss.n602 7.17831
R897 dvss.n75 dvss.n66 7.17078
R898 dvss.n26 dvss 7.15344
R899 dvss.n76 dvss 7.15344
R900 dvss.n569 dvss.n50 7.1196
R901 dvss.n257 dvss.n256 6.77697
R902 dvss.n486 dvss.n485 6.77697
R903 dvss.n446 dvss.n445 6.77697
R904 dvss.n427 dvss.n151 6.77697
R905 dvss.n387 dvss.n386 6.77697
R906 dvss.n348 dvss.n347 6.77697
R907 dvss.n538 dvss.n537 6.7205
R908 dvss.n216 dvss.n196 6.7005
R909 dvss.n679 dvss.n677 6.56103
R910 dvss.n525 dvss.n104 6.53261
R911 dvss.n230 dvss.n82 6.36591
R912 dvss.n602 dvss.n601 5.73579
R913 dvss.n621 dvss.n34 5.34031
R914 dvss.n598 dvss.n47 5.31835
R915 dvss.n565 dvss.n564 5.28896
R916 dvss.n572 dvss.n86 5.28896
R917 dvss.n609 dvss.n47 4.48642
R918 dvss.n555 dvss.t173 4.3505
R919 dvss.n555 dvss.t184 4.3505
R920 dvss.n556 dvss.t76 4.3505
R921 dvss.n556 dvss.t164 4.3505
R922 dvss.n548 dvss.t16 4.3505
R923 dvss.n548 dvss.t128 4.3505
R924 dvss.n547 dvss.t186 4.3505
R925 dvss.n547 dvss.t160 4.3505
R926 dvss.n529 dvss.n528 4.00961
R927 dvss.n577 dvss.n576 3.89404
R928 dvss.n583 dvss.n582 3.84425
R929 dvss.n602 dvss.n17 3.58941
R930 dvss.n579 dvss.n36 3.56414
R931 dvss.n584 dvss.n583 3.54405
R932 dvss.n251 dvss.n249 3.38874
R933 dvss.n480 dvss.n123 3.38874
R934 dvss.n440 dvss.n140 3.38874
R935 dvss.n150 dvss.n147 3.38874
R936 dvss.n393 dvss.n392 3.38874
R937 dvss.n354 dvss.n353 3.38874
R938 dvss.n666 dvss 3.29747
R939 dvss.n680 dvss.n1 3.21038
R940 dvss.n539 dvss.n96 3.01827
R941 dvss.n650 dvss.n649 2.88227
R942 dvss.n567 dvss.n566 2.75993
R943 dvss.n566 dvss.n565 2.75993
R944 dvss.n568 dvss.n87 2.75993
R945 dvss.n564 dvss.n87 2.75993
R946 dvss.n563 dvss.n91 2.64473
R947 dvss.n264 dvss.n263 2.63579
R948 dvss.n493 dvss.n492 2.63579
R949 dvss.n453 dvss.n452 2.63579
R950 dvss.n419 dvss.n154 2.63579
R951 dvss.n380 dvss.n172 2.63579
R952 dvss.n341 dvss.n189 2.63579
R953 dvss.n632 dvss.n22 2.47305
R954 dvss.n67 dvss.n65 2.41042
R955 dvss.n634 dvss.n22 2.33976
R956 dvss.n530 dvss.n96 2.3185
R957 dvss.n575 dvss.n82 1.98969
R958 dvss.n677 dvss.n1 1.93239
R959 dvss.n41 dvss.n36 1.92484
R960 dvss.n272 dvss.n271 1.88285
R961 dvss.n501 dvss.n500 1.88285
R962 dvss.n461 dvss.n460 1.88285
R963 dvss.n413 dvss.n412 1.88285
R964 dvss.n374 dvss.n373 1.88285
R965 dvss.n335 dvss.n334 1.88285
R966 dvss.n103 dvss.n102 1.85983
R967 dvss.n597 dvss.n46 1.80934
R968 dvss.n560 dvss.n559 1.57196
R969 dvss.n551 dvss.n550 1.57139
R970 dvss.n208 dvss.n194 1.5505
R971 dvss.n618 dvss.n18 1.48151
R972 dvss.n34 dvss.n18 1.48151
R973 dvss.n585 dvss.n584 1.46336
R974 dvss.n654 dvss.n14 1.32907
R975 dvss.n591 dvss.n590 1.32907
R976 dvss.n530 dvss.n529 1.21052
R977 dvss.n326 dvss.n196 1.11858
R978 dvss.n566 dvss.n87 1.10724
R979 dvss.n571 dvss.n88 1.10724
R980 dvss.n579 dvss.n37 1.01868
R981 dvss.n567 dvss.n89 0.899376
R982 dvss.n618 dvss.n19 0.804872
R983 dvss.n593 dvss.n38 0.778315
R984 dvss.n575 dvss.n574 0.774309
R985 dvss.n574 dvss.n573 0.774309
R986 dvss.n214 dvss.n208 0.649775
R987 dvss.n296 dvss.n295 0.630008
R988 dvss.n310 dvss.n205 0.630008
R989 dvss.n536 dvss.n89 0.629714
R990 dvss.n620 dvss.n18 0.538751
R991 dvss.n610 dvss.n46 0.533285
R992 dvss.n233 dvss.n232 0.519117
R993 dvss.n234 dvss.n233 0.519117
R994 dvss.n535 dvss.n533 0.482579
R995 dvss.t170 dvss.n657 0.474702
R996 dvss.n657 dvss.n656 0.447064
R997 dvss.n529 dvss.n100 0.443357
R998 dvss.n531 dvss.n530 0.443357
R999 dvss.n227 dvss.n104 0.428132
R1000 dvss.n227 dvss.n146 0.428132
R1001 dvss.n522 dvss.n104 0.411509
R1002 dvss.n616 dvss.n38 0.362946
R1003 dvss.n526 dvss.n90 0.355045
R1004 dvss.n211 dvss.n90 0.355045
R1005 dvss.n604 dvss.n601 0.336965
R1006 dvss.n600 dvss.n17 0.328522
R1007 dvss.n103 dvss 0.326572
R1008 dvss.n605 dvss.n600 0.326101
R1009 dvss.n592 dvss.n11 0.313726
R1010 dvss.n557 dvss.n82 0.277008
R1011 dvss.n662 dvss.n661 0.274194
R1012 dvss.n534 dvss.n51 0.271039
R1013 dvss.n583 dvss.n78 0.262597
R1014 dvss.n611 dvss.n610 0.2605
R1015 dvss.n612 dvss.n611 0.2605
R1016 dvss.n539 dvss.n538 0.248336
R1017 dvss.n81 dvss.n80 0.218682
R1018 dvss.n608 dvss.n48 0.210906
R1019 dvss.n642 dvss.n641 0.206439
R1020 dvss.n595 dvss.n48 0.202526
R1021 dvss.n187 dvss.t116 0.189075
R1022 dvss.n525 dvss.n524 0.181217
R1023 dvss.n633 dvss.n632 0.178278
R1024 dvss.n582 dvss.n581 0.170143
R1025 dvss.n607 dvss.n606 0.166164
R1026 dvss.n601 dvss.n600 0.155797
R1027 dvss dvss.n660 0.150986
R1028 dvss.n51 dvss.n50 0.145813
R1029 dvss.n325 dvss 0.142307
R1030 dvss.n222 dvss 0.140841
R1031 dvss.n660 dvss.n659 0.13579
R1032 dvss.n607 dvss.n599 0.130165
R1033 dvss.n223 dvss 0.127978
R1034 dvss.n223 dvss.n222 0.123227
R1035 dvss.n532 dvss.n531 0.122311
R1036 dvss.n523 dvss.n106 0.121873
R1037 dvss.n324 dvss.n323 0.120292
R1038 dvss.n323 dvss.n197 0.120292
R1039 dvss.n319 dvss.n197 0.120292
R1040 dvss.n319 dvss.n318 0.120292
R1041 dvss.n318 dvss.n317 0.120292
R1042 dvss.n313 dvss.n312 0.120292
R1043 dvss.n311 dvss.n203 0.120292
R1044 dvss.n307 dvss.n203 0.120292
R1045 dvss.n668 dvss.n667 0.120292
R1046 dvss.n669 dvss.n668 0.120292
R1047 dvss.n669 dvss.n4 0.120292
R1048 dvss.n673 dvss.n4 0.120292
R1049 dvss.n674 dvss.n673 0.120292
R1050 dvss.n675 dvss.n674 0.120292
R1051 dvss.n144 dvss.n143 0.104964
R1052 dvss.n312 dvss 0.104667
R1053 dvss.n594 dvss.n51 0.103194
R1054 dvss.n326 dvss 0.0999624
R1055 dvss.n667 dvss 0.0968542
R1056 dvss.n643 dvss 0.0941255
R1057 dvss.n606 dvss.n605 0.0879466
R1058 dvss.n648 dvss.n647 0.0850455
R1059 dvss.n66 dvss 0.080434
R1060 dvss.n221 dvss 0.0781256
R1061 dvss.n77 dvss.n66 0.0777204
R1062 dvss.n645 dvss 0.0770968
R1063 dvss.n578 dvss.n577 0.0749
R1064 dvss.n524 dvss.n523 0.0737044
R1065 dvss.n568 dvss.n567 0.0724101
R1066 dvss.n570 dvss.n569 0.0724101
R1067 dvss.t115 dvss.t114 0.070611
R1068 dvss.n560 dvss.n554 0.0678684
R1069 dvss.n658 dvss.t170 0.0675999
R1070 dvss.n552 dvss.n551 0.0671667
R1071 dvss.n595 dvss.n594 0.06684
R1072 dvss.n222 dvss.n221 0.0638562
R1073 dvss.n557 dvss 0.0633141
R1074 dvss.n581 dvss.n580 0.0614929
R1075 dvss.n659 dvss.t116 0.060491
R1076 dvss.n201 dvss 0.0603958
R1077 dvss.n313 dvss 0.0603958
R1078 dvss dvss.n306 0.0603958
R1079 dvss.n664 dvss 0.0603958
R1080 dvss.n657 dvss.n11 0.0595861
R1081 dvss.n221 dvss.n8 0.0586797
R1082 dvss.n98 dvss.n9 0.0559625
R1083 dvss.n143 dvss.n49 0.0535781
R1084 dvss.n608 dvss.n607 0.0533794
R1085 dvss.n1 dvss 0.0525833
R1086 dvss.n14 dvss 0.0515042
R1087 dvss.n25 dvss.n20 0.0480207
R1088 dvss.n643 dvss.n642 0.0476863
R1089 dvss.n524 dvss.n105 0.0461989
R1090 dvss.n550 dvss.n549 0.0457733
R1091 dvss.n325 dvss.n324 0.0447708
R1092 dvss.n658 dvss.n10 0.0405094
R1093 dvss.n642 dvss.n21 0.0402727
R1094 dvss.n593 dvss.n592 0.0393298
R1095 dvss.n531 dvss.n100 0.0374705
R1096 dvss.n619 dvss.n618 0.0354727
R1097 dvss dvss.n591 0.0347199
R1098 dvss.n559 dvss 0.0346686
R1099 dvss.n580 dvss.n579 0.0341957
R1100 dvss dvss.n201 0.0330521
R1101 dvss.n306 dvss 0.0330521
R1102 dvss.n19 dvss.n11 0.0323493
R1103 dvss.n656 dvss 0.0323446
R1104 dvss.n534 dvss.n89 0.0321327
R1105 dvss.n48 dvss.n46 0.0315
R1106 dvss.n581 dvss.n578 0.0306418
R1107 dvss.n532 dvss.n99 0.0284126
R1108 dvss dvss.n662 0.0271393
R1109 dvss.n592 dvss 0.0255
R1110 dvss.n641 dvss.n22 0.0247851
R1111 dvss.n641 dvss.n640 0.0242603
R1112 dvss.n25 dvss 0.0242603
R1113 dvss.n21 dvss 0.0242603
R1114 dvss.n536 dvss.n535 0.0239848
R1115 dvss.n664 dvss 0.0239375
R1116 dvss.n647 dvss.n645 0.0230951
R1117 dvss.n549 dvss.n10 0.0228519
R1118 dvss.n317 dvss 0.0226354
R1119 dvss.n307 dvss 0.0226354
R1120 dvss.n78 dvss 0.0215598
R1121 dvss.n8 dvss 0.0206613
R1122 dvss.n231 dvss.n9 0.0206307
R1123 dvss.n663 dvss 0.0199672
R1124 dvss.n523 dvss.n522 0.0192879
R1125 dvss.n521 dvss.n520 0.0189524
R1126 dvss.n596 dvss.n595 0.0189524
R1127 dvss.n558 dvss.n557 0.0184385
R1128 dvss.n67 dvss 0.0174837
R1129 dvss.n578 dvss.n79 0.0174213
R1130 dvss.n609 dvss.n608 0.0166458
R1131 dvss dvss.n311 0.016125
R1132 dvss.n432 dvss.n431 0.015957
R1133 dvss.n431 dvss.n430 0.015957
R1134 dvss.n430 dvss.n148 0.015957
R1135 dvss.n426 dvss.n148 0.015957
R1136 dvss.n426 dvss.n425 0.015957
R1137 dvss.n425 dvss.n152 0.015957
R1138 dvss.n421 dvss.n152 0.015957
R1139 dvss.n421 dvss.n420 0.015957
R1140 dvss.n420 dvss.n155 0.015957
R1141 dvss.n416 dvss.n155 0.015957
R1142 dvss.n416 dvss.n415 0.015957
R1143 dvss.n415 dvss.n414 0.015957
R1144 dvss.n414 dvss.n157 0.015957
R1145 dvss.n409 dvss.n157 0.015957
R1146 dvss.n409 dvss.n408 0.015957
R1147 dvss.n408 dvss.n407 0.015957
R1148 dvss.n407 dvss.n160 0.015957
R1149 dvss.n403 dvss.n160 0.015957
R1150 dvss.n403 dvss.n402 0.015957
R1151 dvss.n402 dvss.n401 0.015957
R1152 dvss.n401 dvss.n162 0.015957
R1153 dvss.n397 dvss.n162 0.015957
R1154 dvss.n395 dvss.n165 0.015957
R1155 dvss.n390 dvss.n165 0.015957
R1156 dvss.n390 dvss.n389 0.015957
R1157 dvss.n389 dvss.n388 0.015957
R1158 dvss.n388 dvss.n168 0.015957
R1159 dvss.n383 dvss.n168 0.015957
R1160 dvss.n383 dvss.n382 0.015957
R1161 dvss.n382 dvss.n381 0.015957
R1162 dvss.n381 dvss.n170 0.015957
R1163 dvss.n377 dvss.n170 0.015957
R1164 dvss.n377 dvss.n376 0.015957
R1165 dvss.n376 dvss.n375 0.015957
R1166 dvss.n375 dvss.n174 0.015957
R1167 dvss.n370 dvss.n174 0.015957
R1168 dvss.n370 dvss.n369 0.015957
R1169 dvss.n369 dvss.n368 0.015957
R1170 dvss.n368 dvss.n177 0.015957
R1171 dvss.n364 dvss.n177 0.015957
R1172 dvss.n364 dvss.n363 0.015957
R1173 dvss.n363 dvss.n362 0.015957
R1174 dvss.n362 dvss.n179 0.015957
R1175 dvss.n358 dvss.n179 0.015957
R1176 dvss.n356 dvss.n182 0.015957
R1177 dvss.n351 dvss.n182 0.015957
R1178 dvss.n351 dvss.n350 0.015957
R1179 dvss.n350 dvss.n349 0.015957
R1180 dvss.n349 dvss.n185 0.015957
R1181 dvss.n344 dvss.n185 0.015957
R1182 dvss.n344 dvss.n343 0.015957
R1183 dvss.n343 dvss.n342 0.015957
R1184 dvss.n339 dvss.n338 0.015957
R1185 dvss.n338 dvss.n337 0.015957
R1186 dvss.n337 dvss.n191 0.015957
R1187 dvss.n332 dvss.n191 0.015957
R1188 dvss.n332 dvss.n331 0.015957
R1189 dvss.n331 dvss.n330 0.015957
R1190 dvss.n326 dvss.n325 0.0141555
R1191 dvss.n644 dvss.n643 0.0140978
R1192 dvss.n640 dvss 0.0139298
R1193 dvss.n441 dvss.n141 0.0125293
R1194 dvss.n442 dvss.n441 0.0125293
R1195 dvss.n442 dvss.n138 0.0125293
R1196 dvss.n447 dvss.n138 0.0125293
R1197 dvss.n448 dvss.n447 0.0125293
R1198 dvss.n449 dvss.n448 0.0125293
R1199 dvss.n449 dvss.n135 0.0125293
R1200 dvss.n454 dvss.n135 0.0125293
R1201 dvss.n455 dvss.n454 0.0125293
R1202 dvss.n456 dvss.n455 0.0125293
R1203 dvss.n456 dvss.n133 0.0125293
R1204 dvss.n462 dvss.n133 0.0125293
R1205 dvss.n463 dvss.n462 0.0125293
R1206 dvss.n464 dvss.n463 0.0125293
R1207 dvss.n464 dvss.n131 0.0125293
R1208 dvss.n468 dvss.n131 0.0125293
R1209 dvss.n469 dvss.n468 0.0125293
R1210 dvss.n470 dvss.n469 0.0125293
R1211 dvss.n470 dvss.n129 0.0125293
R1212 dvss.n474 dvss.n129 0.0125293
R1213 dvss.n475 dvss.n474 0.0125293
R1214 dvss.n476 dvss.n475 0.0125293
R1215 dvss.n481 dvss.n124 0.0125293
R1216 dvss.n482 dvss.n481 0.0125293
R1217 dvss.n482 dvss.n121 0.0125293
R1218 dvss.n487 dvss.n121 0.0125293
R1219 dvss.n488 dvss.n487 0.0125293
R1220 dvss.n489 dvss.n488 0.0125293
R1221 dvss.n489 dvss.n118 0.0125293
R1222 dvss.n494 dvss.n118 0.0125293
R1223 dvss.n495 dvss.n494 0.0125293
R1224 dvss.n496 dvss.n495 0.0125293
R1225 dvss.n496 dvss.n116 0.0125293
R1226 dvss.n502 dvss.n116 0.0125293
R1227 dvss.n503 dvss.n502 0.0125293
R1228 dvss.n504 dvss.n503 0.0125293
R1229 dvss.n504 dvss.n114 0.0125293
R1230 dvss.n508 dvss.n114 0.0125293
R1231 dvss.n509 dvss.n508 0.0125293
R1232 dvss.n510 dvss.n509 0.0125293
R1233 dvss.n510 dvss.n112 0.0125293
R1234 dvss.n514 dvss.n112 0.0125293
R1235 dvss.n515 dvss.n514 0.0125293
R1236 dvss.n516 dvss.n515 0.0125293
R1237 dvss.n252 dvss.n250 0.0125293
R1238 dvss.n253 dvss.n252 0.0125293
R1239 dvss.n253 dvss.n247 0.0125293
R1240 dvss.n258 dvss.n247 0.0125293
R1241 dvss.n259 dvss.n258 0.0125293
R1242 dvss.n260 dvss.n259 0.0125293
R1243 dvss.n260 dvss.n244 0.0125293
R1244 dvss.n265 dvss.n244 0.0125293
R1245 dvss.n266 dvss.n265 0.0125293
R1246 dvss.n267 dvss.n266 0.0125293
R1247 dvss.n267 dvss.n242 0.0125293
R1248 dvss.n273 dvss.n242 0.0125293
R1249 dvss.n274 dvss.n273 0.0125293
R1250 dvss.n275 dvss.n274 0.0125293
R1251 dvss.n275 dvss.n240 0.0125293
R1252 dvss.n279 dvss.n240 0.0125293
R1253 dvss.n280 dvss.n279 0.0125293
R1254 dvss.n281 dvss.n280 0.0125293
R1255 dvss.n281 dvss.n238 0.0125293
R1256 dvss.n285 dvss.n238 0.0125293
R1257 dvss.n286 dvss.n285 0.0125293
R1258 dvss.n287 dvss.n286 0.0125293
R1259 dvss.n292 dvss.n291 0.0125293
R1260 dvss.n298 dvss.n297 0.0125293
R1261 dvss.n299 dvss.n298 0.0125293
R1262 dvss.n339 dvss.n187 0.0122608
R1263 dvss dvss.n558 0.0110353
R1264 dvss.n292 dvss 0.0109603
R1265 dvss.n78 dvss.n77 0.0106902
R1266 dvss.n659 dvss.t115 0.0106199
R1267 dvss.n580 dvss.n53 0.0101631
R1268 dvss.n327 dvss.n194 0.0099086
R1269 dvss.n661 dvss.n8 0.00990439
R1270 dvss.n660 dvss.n9 0.00933152
R1271 dvss.n675 dvss.n1 0.0083125
R1272 dvss.n642 dvss.n20 0.00824793
R1273 dvss.n535 dvss.n534 0.00822968
R1274 dvss.n432 dvss 0.00822849
R1275 dvss dvss.n396 0.00822849
R1276 dvss dvss.n395 0.00822849
R1277 dvss dvss.n357 0.00822849
R1278 dvss dvss.n356 0.00822849
R1279 dvss.n647 dvss.n646 0.00789958
R1280 dvss.n330 dvss.n194 0.00654839
R1281 dvss.n141 dvss 0.00651464
R1282 dvss dvss.n125 0.00651464
R1283 dvss dvss.n124 0.00651464
R1284 dvss.n250 dvss 0.00651464
R1285 dvss.n290 dvss 0.00651464
R1286 dvss.n291 dvss 0.00651464
R1287 dvss dvss.n224 0.00651464
R1288 dvss.n520 dvss.n519 0.00573013
R1289 dvss dvss.n1 0.00570833
R1290 dvss.n557 dvss.n10 0.00519818
R1291 dvss.n661 dvss 0.00481034
R1292 dvss dvss.n105 0.00470027
R1293 dvss.n396 dvss 0.00470027
R1294 dvss.n357 dvss 0.00470027
R1295 dvss.n342 dvss.n187 0.00419624
R1296 dvss.n645 dvss.n644 0.00411776
R1297 dvss dvss.n106 0.00376883
R1298 dvss.n125 dvss 0.00376883
R1299 dvss.n519 dvss 0.00376883
R1300 dvss dvss.n290 0.00376883
R1301 dvss.n224 dvss 0.00376883
R1302 dvss.t114 dvss.n658 0.00351108
R1303 dvss.n397 dvss 0.00335618
R1304 dvss.n358 dvss 0.00335618
R1305 dvss.n476 dvss 0.0027228
R1306 dvss.n516 dvss 0.0027228
R1307 dvss.n287 dvss 0.0027228
R1308 dvss.n299 dvss 0.0027228
R1309 dvss.n297 dvss 0.00206904
R1310 dvss dvss.n663 0.00180208
R1311 dvss.n533 dvss.n532 0.00156293
R1312 dvss.n663 dvss 0.00152459
R1313 dvss.n327 dvss.n326 0.00150806
R1314 dvss.n520 dvss 0.00128452
R1315 dvss dvss.n223 0.00077533
R1316 dvss.n646 dvss.n14 0.000632135
R1317 dvss.n591 dvss.n53 0.000588652
R1318 x7.stby_done_b.n8 x7.stby_done_b.t0 373.866
R1319 x7.stby_done_b.n6 x7.stby_done_b.t6 333.651
R1320 x7.stby_done_b.n6 x7.stby_done_b.t2 297.233
R1321 x7.stby_done_b.n1 x7.stby_done_b.t5 241.536
R1322 x7.stby_done_b x7.stby_done_b.t1 237.101
R1323 x7.stby_done_b.n4 x7.stby_done_b.t3 207.423
R1324 x7.stby_done_b.n3 x7.stby_done_b.t4 202.133
R1325 x7.stby_done_b x7.stby_done_b.n6 195.701
R1326 x7.stby_done_b.n1 x7.stby_done_b.t7 169.237
R1327 x7.stby_done_b.n5 x7.stby_done_b.n4 159.758
R1328 x7.stby_done_b.n3 x7.stby_done_b 154.91
R1329 x7.stby_done_b.n2 x7.stby_done_b.n1 152
R1330 x7.stby_done_b.n4 x7.stby_done_b.n3 36.8275
R1331 x7.stby_done_b x7.stby_done_b.n8 26.7478
R1332 x7.stby_done_b.n7 x7.stby_done_b 15.8995
R1333 x7.stby_done_b.n7 x7.stby_done_b.n0 15.8481
R1334 x7.stby_done_b.n0 x7.stby_done_b.n5 13.8109
R1335 x7.stby_done_b x7.stby_done_b.n2 13.3943
R1336 x7.stby_done_b.n8 x7.stby_done_b.n7 3.1005
R1337 x7.stby_done_b.n5 x7.stby_done_b 2.52171
R1338 x7.stby_done_b.n2 x7.stby_done_b 1.9205
R1339 x7.stby_done_b.n0 x7.stby_done_b 1.418
R1340 dvdd.n295 dvdd.n286 5128.23
R1341 dvdd.n295 dvdd.n287 5128.23
R1342 dvdd.n293 dvdd.n287 5128.23
R1343 dvdd.n293 dvdd.n286 5128.23
R1344 dvdd.n42 dvdd.n5 1736.47
R1345 dvdd.n45 dvdd.n4 1736.47
R1346 dvdd.n30 dvdd.n27 1736.47
R1347 dvdd.n33 dvdd.n29 1736.47
R1348 dvdd.n255 dvdd.t25 838.817
R1349 dvdd.n69 dvdd.t162 806.511
R1350 dvdd.n69 dvdd.t89 806.511
R1351 dvdd.n90 dvdd.t125 806.511
R1352 dvdd.n90 dvdd.t77 806.511
R1353 dvdd.n111 dvdd.t96 806.511
R1354 dvdd.n111 dvdd.t7 806.511
R1355 dvdd.n292 dvdd.n284 787.447
R1356 dvdd.n292 dvdd.n285 786.827
R1357 dvdd.n56 dvdd.t114 668.683
R1358 dvdd.n56 dvdd.t133 668.683
R1359 dvdd.n227 dvdd.t42 667.778
R1360 dvdd.n227 dvdd.t140 667.778
R1361 dvdd.n189 dvdd.t154 667.778
R1362 dvdd.n189 dvdd.t23 667.778
R1363 dvdd.n151 dvdd.t61 667.778
R1364 dvdd.n151 dvdd.t18 667.778
R1365 dvdd.n296 dvdd.n284 604.574
R1366 dvdd.n73 dvdd.n71 604.457
R1367 dvdd.n73 dvdd.n72 604.457
R1368 dvdd.n94 dvdd.n92 604.457
R1369 dvdd.n94 dvdd.n93 604.457
R1370 dvdd.n115 dvdd.n113 604.457
R1371 dvdd.n115 dvdd.n114 604.457
R1372 dvdd.n232 dvdd.n61 604.394
R1373 dvdd.n232 dvdd.n62 604.394
R1374 dvdd.n194 dvdd.n82 604.394
R1375 dvdd.n194 dvdd.n83 604.394
R1376 dvdd.n156 dvdd.n103 604.394
R1377 dvdd.n156 dvdd.n104 604.394
R1378 dvdd.n220 dvdd.n67 601.679
R1379 dvdd.n220 dvdd.n68 601.679
R1380 dvdd.n182 dvdd.n88 601.679
R1381 dvdd.n182 dvdd.n89 601.679
R1382 dvdd.n144 dvdd.n109 601.679
R1383 dvdd.n144 dvdd.n110 601.679
R1384 dvdd.n260 dvdd.n259 585
R1385 dvdd.t155 dvdd.t24 556.386
R1386 dvdd.n246 dvdd 538.664
R1387 dvdd.n18 dvdd 535.705
R1388 dvdd.n11 dvdd 535.705
R1389 dvdd.t86 dvdd 473.521
R1390 dvdd.t17 dvdd.t20 448.146
R1391 dvdd.t22 dvdd.t164 448.146
R1392 dvdd.t41 dvdd.t55 448.146
R1393 dvdd.n296 dvdd.n285 423.062
R1394 dvdd.t31 dvdd.t102 367.579
R1395 dvdd.t120 dvdd.t44 367.579
R1396 dvdd.t65 dvdd.t98 367.579
R1397 dvdd.n274 dvdd.t58 360.005
R1398 dvdd.t6 dvdd.t47 330.654
R1399 dvdd.t76 dvdd.t26 330.654
R1400 dvdd.t88 dvdd.t72 330.654
R1401 dvdd.n43 dvdd.n4 314.781
R1402 dvdd.n44 dvdd.n5 314.781
R1403 dvdd.n31 dvdd.n29 314.781
R1404 dvdd.n32 dvdd.n27 314.781
R1405 dvdd.n23 dvdd.n17 312.053
R1406 dvdd.n9 dvdd.n8 312.051
R1407 dvdd.n266 dvdd.n256 312.051
R1408 dvdd.t53 dvdd.t51 304.829
R1409 dvdd.t24 dvdd.t13 284.113
R1410 dvdd.t102 dvdd.t8 275.265
R1411 dvdd.t44 dvdd.t39 275.265
R1412 dvdd.t98 dvdd.t11 275.265
R1413 dvdd.t13 dvdd.t86 275.235
R1414 dvdd.n271 dvdd.t33 261.837
R1415 dvdd.t37 dvdd.t152 260.437
R1416 dvdd.t156 dvdd.t82 260.437
R1417 dvdd.n207 dvdd.n76 259.707
R1418 dvdd.n207 dvdd.n75 259.707
R1419 dvdd.n169 dvdd.n97 259.707
R1420 dvdd.n169 dvdd.n96 259.707
R1421 dvdd.n131 dvdd.n118 259.707
R1422 dvdd.n131 dvdd.n117 259.707
R1423 dvdd.t33 dvdd.t15 258.481
R1424 dvdd.n273 dvdd.t146 253.446
R1425 dvdd.n272 dvdd.t0 253.446
R1426 dvdd.t43 dvdd.t160 248.599
R1427 dvdd.t160 dvdd.t155 248.599
R1428 dvdd.n201 dvdd.n80 242.607
R1429 dvdd.n163 dvdd.n101 242.607
R1430 dvdd.n125 dvdd.n123 242.607
R1431 dvdd.n201 dvdd.n79 242.607
R1432 dvdd.n163 dvdd.n100 242.607
R1433 dvdd.n125 dvdd.n122 242.607
R1434 dvdd.t2 dvdd.t174 234.982
R1435 dvdd.t63 dvdd.t19 234.982
R1436 dvdd.t84 dvdd.t132 234.982
R1437 dvdd dvdd.n270 232.445
R1438 dvdd.n0 dvdd.t79 228.215
R1439 dvdd.n0 dvdd.t5 228.215
R1440 dvdd.n239 dvdd.n59 215.123
R1441 dvdd.n239 dvdd.n238 215.123
R1442 dvdd.t51 dvdd.t134 213.084
R1443 dvdd.n41 dvdd.n3 185.225
R1444 dvdd.n46 dvdd.n3 185.225
R1445 dvdd.n34 dvdd.n28 185.225
R1446 dvdd.n28 dvdd.n26 185.225
R1447 dvdd.t105 dvdd.t137 181.273
R1448 dvdd.t74 dvdd.t68 181.273
R1449 dvdd.t126 dvdd.t28 181.273
R1450 dvdd.t70 dvdd.t6 166.167
R1451 dvdd.t174 dvdd.t141 166.167
R1452 dvdd.t119 dvdd.t76 166.167
R1453 dvdd.t19 dvdd.t30 166.167
R1454 dvdd.t131 dvdd.t88 166.167
R1455 dvdd.t132 dvdd.t150 166.167
R1456 dvdd.t58 dvdd.t31 162.81
R1457 dvdd.t47 dvdd.t2 162.81
R1458 dvdd.t146 dvdd.t120 162.81
R1459 dvdd.t26 dvdd.t63 162.81
R1460 dvdd.t0 dvdd.t65 162.81
R1461 dvdd.t72 dvdd.t84 162.81
R1462 dvdd.t94 dvdd.n293 161.316
R1463 dvdd.n295 dvdd.t115 161.316
R1464 dvdd.t141 dvdd.t17 154.417
R1465 dvdd.t30 dvdd.t22 154.417
R1466 dvdd.t150 dvdd.t41 154.417
R1467 dvdd.t15 dvdd.t113 147.703
R1468 dvdd.n75 dvdd.t12 147.111
R1469 dvdd.n76 dvdd.t101 147.111
R1470 dvdd.n96 dvdd.t40 147.111
R1471 dvdd.n97 dvdd.t97 147.111
R1472 dvdd.n117 dvdd.t46 147.111
R1473 dvdd.n118 dvdd.t9 147.111
R1474 dvdd.t10 dvdd.t70 144.346
R1475 dvdd.t104 dvdd.t119 144.346
R1476 dvdd.t57 dvdd.t131 144.346
R1477 dvdd.t8 dvdd.t105 140.989
R1478 dvdd.t137 dvdd.t10 140.989
R1479 dvdd.t20 dvdd.t111 140.989
R1480 dvdd.t39 dvdd.t74 140.989
R1481 dvdd.t68 dvdd.t104 140.989
R1482 dvdd.t164 dvdd.t122 140.989
R1483 dvdd.t11 dvdd.t126 140.989
R1484 dvdd.t28 dvdd.t57 140.989
R1485 dvdd.t55 dvdd.t109 140.989
R1486 dvdd.t113 dvdd 132.597
R1487 dvdd dvdd.n273 125.883
R1488 dvdd dvdd.n272 125.883
R1489 dvdd dvdd.n271 125.883
R1490 dvdd.t144 dvdd.t94 121.245
R1491 dvdd.t142 dvdd.t144 121.245
R1492 dvdd.t49 dvdd.t142 121.245
R1493 dvdd.t169 dvdd.t49 121.245
R1494 dvdd.t92 dvdd.t117 121.245
R1495 dvdd.t80 dvdd.t92 121.245
R1496 dvdd.t35 dvdd.t80 121.245
R1497 dvdd.t115 dvdd.t35 121.245
R1498 dvdd.n71 dvdd.t60 119.608
R1499 dvdd.n72 dvdd.t29 119.608
R1500 dvdd.n92 dvdd.t69 119.608
R1501 dvdd.n93 dvdd.t136 119.608
R1502 dvdd.n113 dvdd.t138 119.608
R1503 dvdd.n114 dvdd.t171 119.608
R1504 dvdd.t111 dvdd 109.1
R1505 dvdd.t122 dvdd 109.1
R1506 dvdd.t109 dvdd 109.1
R1507 dvdd.n75 dvdd.t151 108.413
R1508 dvdd.n76 dvdd.t99 108.413
R1509 dvdd.n96 dvdd.t45 108.413
R1510 dvdd.n97 dvdd.t108 108.413
R1511 dvdd.n117 dvdd.t103 108.413
R1512 dvdd.n118 dvdd.t148 108.413
R1513 dvdd.n271 dvdd.n55 106.559
R1514 dvdd.n272 dvdd.n54 106.559
R1515 dvdd.n273 dvdd.n53 106.559
R1516 dvdd.n47 dvdd.n2 105.412
R1517 dvdd.n40 dvdd.n2 105.412
R1518 dvdd.n37 dvdd.n36 105.412
R1519 dvdd.n36 dvdd.n35 105.412
R1520 dvdd dvdd.t53 100.624
R1521 dvdd.n67 dvdd.t85 93.81
R1522 dvdd.n68 dvdd.t100 93.81
R1523 dvdd.n88 dvdd.t163 93.81
R1524 dvdd.n89 dvdd.t64 93.81
R1525 dvdd.n109 dvdd.t67 93.81
R1526 dvdd.n110 dvdd.t3 93.81
R1527 dvdd dvdd.t37 91.745
R1528 dvdd dvdd.t156 91.745
R1529 dvdd dvdd.t43 88.7855
R1530 dvdd.n259 dvdd.t54 86.7743
R1531 dvdd.n47 dvdd.n46 79.8123
R1532 dvdd.n41 dvdd.n40 79.8123
R1533 dvdd.n35 dvdd.n34 79.8123
R1534 dvdd.n37 dvdd.n26 79.8123
R1535 dvdd.n59 dvdd.t62 74.7554
R1536 dvdd.n238 dvdd.t16 74.7554
R1537 dvdd.n67 dvdd.t128 63.3219
R1538 dvdd.n68 dvdd.t73 63.3219
R1539 dvdd.n71 dvdd.t127 63.3219
R1540 dvdd.n72 dvdd.t129 63.3219
R1541 dvdd.n88 dvdd.t149 63.3219
R1542 dvdd.n89 dvdd.t27 63.3219
R1543 dvdd.n92 dvdd.t130 63.3219
R1544 dvdd.n93 dvdd.t75 63.3219
R1545 dvdd.n109 dvdd.t167 63.3219
R1546 dvdd.n110 dvdd.t48 63.3219
R1547 dvdd.n113 dvdd.t159 63.3219
R1548 dvdd.n114 dvdd.t106 63.3219
R1549 dvdd.n79 dvdd.t66 61.9829
R1550 dvdd.n100 dvdd.t121 61.9829
R1551 dvdd.n122 dvdd.t124 61.9829
R1552 dvdd.n80 dvdd.t90 61.9826
R1553 dvdd.n101 dvdd.t139 61.9826
R1554 dvdd.n123 dvdd.t32 61.9826
R1555 dvdd.n259 dvdd.t52 61.05
R1556 dvdd.n294 dvdd.t169 60.6225
R1557 dvdd.t117 dvdd.n294 60.6225
R1558 dvdd.n292 dvdd.t95 60.3236
R1559 dvdd.n296 dvdd.t116 60.3236
R1560 dvdd.n297 dvdd.n283 54.7085
R1561 dvdd.n298 dvdd.n282 54.7085
R1562 dvdd.n290 dvdd.n289 54.7085
R1563 dvdd.n291 dvdd.n288 54.7085
R1564 dvdd.n61 dvdd.t161 41.5552
R1565 dvdd.n61 dvdd.t173 41.5552
R1566 dvdd.n62 dvdd.t56 41.5552
R1567 dvdd.n62 dvdd.t110 41.5552
R1568 dvdd.n82 dvdd.t165 41.5552
R1569 dvdd.n82 dvdd.t172 41.5552
R1570 dvdd.n83 dvdd.t168 41.5552
R1571 dvdd.n83 dvdd.t123 41.5552
R1572 dvdd.n103 dvdd.t71 41.5552
R1573 dvdd.n103 dvdd.t112 41.5552
R1574 dvdd.n104 dvdd.t21 41.5552
R1575 dvdd.n104 dvdd.t135 41.5552
R1576 dvdd.n46 dvdd.n45 37.0005
R1577 dvdd.n42 dvdd.n41 37.0005
R1578 dvdd.n34 dvdd.n33 37.0005
R1579 dvdd.n30 dvdd.n26 37.0005
R1580 dvdd.n17 dvdd.t38 36.1587
R1581 dvdd.n17 dvdd.t153 36.1587
R1582 dvdd.n8 dvdd.t157 36.1587
R1583 dvdd.n8 dvdd.t83 36.1587
R1584 dvdd.n256 dvdd.t14 35.4605
R1585 dvdd.n250 dvdd.n249 34.6358
R1586 dvdd.n254 dvdd.n245 34.6358
R1587 dvdd.n265 dvdd.n257 34.6358
R1588 dvdd.n231 dvdd.n63 34.6358
R1589 dvdd.n221 dvdd.n65 34.6358
R1590 dvdd.n225 dvdd.n65 34.6358
R1591 dvdd.n226 dvdd.n225 34.6358
R1592 dvdd.n219 dvdd.n218 34.6358
R1593 dvdd.n213 dvdd.n212 34.6358
R1594 dvdd.n214 dvdd.n213 34.6358
R1595 dvdd.n200 dvdd.n199 34.6358
R1596 dvdd.n202 dvdd.n77 34.6358
R1597 dvdd.n206 dvdd.n77 34.6358
R1598 dvdd.n193 dvdd.n84 34.6358
R1599 dvdd.n183 dvdd.n86 34.6358
R1600 dvdd.n187 dvdd.n86 34.6358
R1601 dvdd.n188 dvdd.n187 34.6358
R1602 dvdd.n181 dvdd.n180 34.6358
R1603 dvdd.n175 dvdd.n174 34.6358
R1604 dvdd.n176 dvdd.n175 34.6358
R1605 dvdd.n162 dvdd.n161 34.6358
R1606 dvdd.n164 dvdd.n98 34.6358
R1607 dvdd.n168 dvdd.n98 34.6358
R1608 dvdd.n155 dvdd.n105 34.6358
R1609 dvdd.n145 dvdd.n107 34.6358
R1610 dvdd.n149 dvdd.n107 34.6358
R1611 dvdd.n150 dvdd.n149 34.6358
R1612 dvdd.n143 dvdd.n142 34.6358
R1613 dvdd.n137 dvdd.n136 34.6358
R1614 dvdd.n138 dvdd.n137 34.6358
R1615 dvdd.n124 dvdd.n52 34.6358
R1616 dvdd.n126 dvdd.n119 34.6358
R1617 dvdd.n130 dvdd.n119 34.6358
R1618 dvdd.n239 dvdd.n58 33.8829
R1619 dvdd.n227 dvdd.n226 32.377
R1620 dvdd.n189 dvdd.n188 32.377
R1621 dvdd.n151 dvdd.n150 32.377
R1622 dvdd.n214 dvdd.n69 32.0005
R1623 dvdd.n176 dvdd.n90 32.0005
R1624 dvdd.n138 dvdd.n111 32.0005
R1625 dvdd.n240 dvdd.n239 31.624
R1626 dvdd.n202 dvdd.n201 31.2476
R1627 dvdd.n164 dvdd.n163 31.2476
R1628 dvdd.n126 dvdd.n125 31.2476
R1629 dvdd.n5 dvdd.n3 30.8338
R1630 dvdd.n4 dvdd.n2 30.8338
R1631 dvdd.n36 dvdd.n27 30.8338
R1632 dvdd.n29 dvdd.n28 30.8338
R1633 dvdd.n79 dvdd.t1 30.1745
R1634 dvdd.n100 dvdd.t158 30.1745
R1635 dvdd.n122 dvdd.t166 30.1745
R1636 dvdd.n80 dvdd.t91 30.1738
R1637 dvdd.n101 dvdd.t147 30.1738
R1638 dvdd.n123 dvdd.t59 30.1738
R1639 dvdd.n208 dvdd.n73 30.1181
R1640 dvdd.n170 dvdd.n94 30.1181
R1641 dvdd.n132 dvdd.n115 30.1181
R1642 dvdd.n43 dvdd.n42 29.6618
R1643 dvdd.n45 dvdd.n44 29.6618
R1644 dvdd.n31 dvdd.n30 29.6618
R1645 dvdd.n33 dvdd.n32 29.6618
R1646 dvdd.n59 dvdd.t34 28.5349
R1647 dvdd.n238 dvdd.t107 28.5349
R1648 dvdd.n261 dvdd.n257 28.2952
R1649 dvdd dvdd.n245 27.8593
R1650 dvdd.n256 dvdd.t87 26.5955
R1651 dvdd.n260 dvdd.n258 25.2079
R1652 dvdd.n22 dvdd.n18 23.7181
R1653 dvdd.n11 dvdd.n10 23.7181
R1654 dvdd.n249 dvdd.n246 23.7181
R1655 dvdd.n233 dvdd.n55 23.7181
R1656 dvdd.n199 dvdd.n54 23.7181
R1657 dvdd.n195 dvdd.n54 23.7181
R1658 dvdd.n161 dvdd.n53 23.7181
R1659 dvdd.n157 dvdd.n53 23.7181
R1660 dvdd.n274 dvdd.n52 23.7181
R1661 dvdd.n58 dvdd.n55 23.7181
R1662 dvdd.n232 dvdd.n231 22.9652
R1663 dvdd.n194 dvdd.n193 22.9652
R1664 dvdd.n156 dvdd.n155 22.9652
R1665 dvdd.n267 dvdd.n255 22.5887
R1666 dvdd.n266 dvdd.n265 22.5887
R1667 dvdd.n267 dvdd.n266 21.8358
R1668 dvdd.n233 dvdd.n232 21.4593
R1669 dvdd.n195 dvdd.n194 21.4593
R1670 dvdd.n157 dvdd.n156 21.4593
R1671 dvdd.n212 dvdd.n73 20.3299
R1672 dvdd.n174 dvdd.n94 20.3299
R1673 dvdd.n136 dvdd.n115 20.3299
R1674 dvdd.n255 dvdd.n254 19.9534
R1675 dvdd.n240 dvdd.n56 19.577
R1676 dvdd.n270 dvdd.n56 18.4476
R1677 dvdd.n227 dvdd.n63 18.0711
R1678 dvdd.n189 dvdd.n84 18.0711
R1679 dvdd.n151 dvdd.n105 18.0711
R1680 dvdd.n23 dvdd 15.8123
R1681 dvdd dvdd.n9 15.8123
R1682 dvdd.n296 dvdd.n295 13.2148
R1683 dvdd.n293 dvdd.n292 13.2148
R1684 dvdd.n38 dvdd.n37 10.0436
R1685 dvdd.n35 dvdd.n1 9.59217
R1686 dvdd.n218 dvdd.n69 9.41227
R1687 dvdd.n180 dvdd.n90 9.41227
R1688 dvdd.n142 dvdd.n111 9.41227
R1689 dvdd.n19 dvdd.n18 9.3005
R1690 dvdd.n22 dvdd.n21 9.3005
R1691 dvdd.n10 dvdd.n6 9.3005
R1692 dvdd.n12 dvdd.n11 9.3005
R1693 dvdd.n40 dvdd.n39 9.3005
R1694 dvdd.n48 dvdd.n47 9.3005
R1695 dvdd.n262 dvdd.n261 9.3005
R1696 dvdd.n263 dvdd.n257 9.3005
R1697 dvdd.n265 dvdd.n264 9.3005
R1698 dvdd.n266 dvdd.n243 9.3005
R1699 dvdd.n255 dvdd.n244 9.3005
R1700 dvdd.n254 dvdd.n253 9.3005
R1701 dvdd.n252 dvdd.n245 9.3005
R1702 dvdd.n251 dvdd.n250 9.3005
R1703 dvdd.n249 dvdd.n248 9.3005
R1704 dvdd.n247 dvdd.n246 9.3005
R1705 dvdd.n270 dvdd.n269 9.3005
R1706 dvdd.n275 dvdd.n274 9.3005
R1707 dvdd.n120 dvdd.n52 9.3005
R1708 dvdd.n124 dvdd.n121 9.3005
R1709 dvdd.n127 dvdd.n126 9.3005
R1710 dvdd.n128 dvdd.n119 9.3005
R1711 dvdd.n130 dvdd.n129 9.3005
R1712 dvdd.n131 dvdd.n116 9.3005
R1713 dvdd.n133 dvdd.n132 9.3005
R1714 dvdd.n134 dvdd.n115 9.3005
R1715 dvdd.n136 dvdd.n135 9.3005
R1716 dvdd.n137 dvdd.n112 9.3005
R1717 dvdd.n139 dvdd.n138 9.3005
R1718 dvdd.n140 dvdd.n111 9.3005
R1719 dvdd.n142 dvdd.n141 9.3005
R1720 dvdd.n143 dvdd.n108 9.3005
R1721 dvdd.n146 dvdd.n145 9.3005
R1722 dvdd.n147 dvdd.n107 9.3005
R1723 dvdd.n149 dvdd.n148 9.3005
R1724 dvdd.n150 dvdd.n106 9.3005
R1725 dvdd.n152 dvdd.n151 9.3005
R1726 dvdd.n153 dvdd.n105 9.3005
R1727 dvdd.n155 dvdd.n154 9.3005
R1728 dvdd.n156 dvdd.n102 9.3005
R1729 dvdd.n158 dvdd.n157 9.3005
R1730 dvdd.n159 dvdd.n53 9.3005
R1731 dvdd.n161 dvdd.n160 9.3005
R1732 dvdd.n162 dvdd.n99 9.3005
R1733 dvdd.n165 dvdd.n164 9.3005
R1734 dvdd.n166 dvdd.n98 9.3005
R1735 dvdd.n168 dvdd.n167 9.3005
R1736 dvdd.n169 dvdd.n95 9.3005
R1737 dvdd.n171 dvdd.n170 9.3005
R1738 dvdd.n172 dvdd.n94 9.3005
R1739 dvdd.n174 dvdd.n173 9.3005
R1740 dvdd.n175 dvdd.n91 9.3005
R1741 dvdd.n177 dvdd.n176 9.3005
R1742 dvdd.n178 dvdd.n90 9.3005
R1743 dvdd.n180 dvdd.n179 9.3005
R1744 dvdd.n181 dvdd.n87 9.3005
R1745 dvdd.n184 dvdd.n183 9.3005
R1746 dvdd.n185 dvdd.n86 9.3005
R1747 dvdd.n187 dvdd.n186 9.3005
R1748 dvdd.n188 dvdd.n85 9.3005
R1749 dvdd.n190 dvdd.n189 9.3005
R1750 dvdd.n191 dvdd.n84 9.3005
R1751 dvdd.n193 dvdd.n192 9.3005
R1752 dvdd.n194 dvdd.n81 9.3005
R1753 dvdd.n196 dvdd.n195 9.3005
R1754 dvdd.n197 dvdd.n54 9.3005
R1755 dvdd.n199 dvdd.n198 9.3005
R1756 dvdd.n200 dvdd.n78 9.3005
R1757 dvdd.n203 dvdd.n202 9.3005
R1758 dvdd.n204 dvdd.n77 9.3005
R1759 dvdd.n206 dvdd.n205 9.3005
R1760 dvdd.n207 dvdd.n74 9.3005
R1761 dvdd.n209 dvdd.n208 9.3005
R1762 dvdd.n210 dvdd.n73 9.3005
R1763 dvdd.n212 dvdd.n211 9.3005
R1764 dvdd.n213 dvdd.n70 9.3005
R1765 dvdd.n215 dvdd.n214 9.3005
R1766 dvdd.n216 dvdd.n69 9.3005
R1767 dvdd.n218 dvdd.n217 9.3005
R1768 dvdd.n219 dvdd.n66 9.3005
R1769 dvdd.n222 dvdd.n221 9.3005
R1770 dvdd.n223 dvdd.n65 9.3005
R1771 dvdd.n225 dvdd.n224 9.3005
R1772 dvdd.n226 dvdd.n64 9.3005
R1773 dvdd.n228 dvdd.n227 9.3005
R1774 dvdd.n229 dvdd.n63 9.3005
R1775 dvdd.n231 dvdd.n230 9.3005
R1776 dvdd.n232 dvdd.n60 9.3005
R1777 dvdd.n234 dvdd.n233 9.3005
R1778 dvdd.n235 dvdd.n55 9.3005
R1779 dvdd.n236 dvdd.n58 9.3005
R1780 dvdd.n239 dvdd.n237 9.3005
R1781 dvdd.n239 dvdd.n57 9.3005
R1782 dvdd.n241 dvdd.n240 9.3005
R1783 dvdd.n242 dvdd.n56 9.3005
R1784 dvdd.n268 dvdd.n267 9.3005
R1785 dvdd.n208 dvdd.n207 9.03579
R1786 dvdd.n170 dvdd.n169 9.03579
R1787 dvdd.n132 dvdd.n131 9.03579
R1788 dvdd.n286 dvdd.n284 7.70883
R1789 dvdd.n294 dvdd.n286 7.70883
R1790 dvdd.n287 dvdd.n285 7.70883
R1791 dvdd.n294 dvdd.n287 7.70883
R1792 dvdd.n24 dvdd.n23 7.17001
R1793 dvdd.n9 dvdd.n7 7.15376
R1794 dvdd.n283 dvdd.t81 7.14175
R1795 dvdd.n283 dvdd.t36 7.14175
R1796 dvdd.n282 dvdd.t118 7.14175
R1797 dvdd.n282 dvdd.t93 7.14175
R1798 dvdd.n289 dvdd.t50 7.14175
R1799 dvdd.n289 dvdd.t170 7.14175
R1800 dvdd.n288 dvdd.t145 7.14175
R1801 dvdd.n288 dvdd.t143 7.14175
R1802 dvdd.n250 dvdd 6.77697
R1803 dvdd.n44 dvdd.t4 6.70818
R1804 dvdd.t4 dvdd.n43 6.70818
R1805 dvdd.n32 dvdd.t78 6.70818
R1806 dvdd.t78 dvdd.n31 6.70818
R1807 dvdd dvdd.n22 6.4005
R1808 dvdd.n10 dvdd 6.4005
R1809 dvdd.n221 dvdd.n220 6.02403
R1810 dvdd.n207 dvdd.n206 6.02403
R1811 dvdd.n183 dvdd.n182 6.02403
R1812 dvdd.n169 dvdd.n168 6.02403
R1813 dvdd.n145 dvdd.n144 6.02403
R1814 dvdd.n131 dvdd.n130 6.02403
R1815 dvdd.n220 dvdd.n219 3.76521
R1816 dvdd.n182 dvdd.n181 3.76521
R1817 dvdd.n144 dvdd.n143 3.76521
R1818 dvdd.n201 dvdd.n200 3.38874
R1819 dvdd.n163 dvdd.n162 3.38874
R1820 dvdd.n125 dvdd.n124 3.38874
R1821 dvdd.n297 dvdd.n296 1.66909
R1822 dvdd.n292 dvdd.n291 1.57188
R1823 dvdd.n36 dvdd.n0 1.32907
R1824 dvdd.n2 dvdd.n0 1.32907
R1825 dvdd.n261 dvdd.n260 1.23559
R1826 dvdd.n276 dvdd.n275 0.637387
R1827 dvdd.n276 dvdd.n51 0.496845
R1828 dvdd dvdd.n268 0.438
R1829 dvdd.n50 dvdd.n49 0.432317
R1830 dvdd.n16 dvdd 0.42713
R1831 dvdd dvdd.n16 0.32387
R1832 dvdd.n268 dvdd 0.313
R1833 dvdd.n247 dvdd.n51 0.280448
R1834 dvdd.n51 dvdd 0.232271
R1835 dvdd.n7 dvdd 0.203706
R1836 dvdd.n13 dvdd 0.167167
R1837 dvdd.n19 dvdd 0.164848
R1838 dvdd.n258 dvdd 0.159538
R1839 dvdd.n38 dvdd.n15 0.141704
R1840 dvdd.n262 dvdd.n258 0.141672
R1841 dvdd.n38 dvdd.n25 0.139389
R1842 dvdd.n14 dvdd.n6 0.127236
R1843 dvdd.n264 dvdd.n243 0.120292
R1844 dvdd.n252 dvdd.n251 0.120292
R1845 dvdd.n253 dvdd.n252 0.120292
R1846 dvdd.n253 dvdd.n244 0.120292
R1847 dvdd.n121 dvdd.n120 0.120292
R1848 dvdd.n127 dvdd.n121 0.120292
R1849 dvdd.n128 dvdd.n127 0.120292
R1850 dvdd.n129 dvdd.n128 0.120292
R1851 dvdd.n129 dvdd.n116 0.120292
R1852 dvdd.n133 dvdd.n116 0.120292
R1853 dvdd.n134 dvdd.n133 0.120292
R1854 dvdd.n135 dvdd.n134 0.120292
R1855 dvdd.n135 dvdd.n112 0.120292
R1856 dvdd.n139 dvdd.n112 0.120292
R1857 dvdd.n140 dvdd.n139 0.120292
R1858 dvdd.n141 dvdd.n140 0.120292
R1859 dvdd.n141 dvdd.n108 0.120292
R1860 dvdd.n146 dvdd.n108 0.120292
R1861 dvdd.n147 dvdd.n146 0.120292
R1862 dvdd.n148 dvdd.n147 0.120292
R1863 dvdd.n148 dvdd.n106 0.120292
R1864 dvdd.n152 dvdd.n106 0.120292
R1865 dvdd.n153 dvdd.n152 0.120292
R1866 dvdd.n154 dvdd.n153 0.120292
R1867 dvdd.n154 dvdd.n102 0.120292
R1868 dvdd.n158 dvdd.n102 0.120292
R1869 dvdd.n160 dvdd.n99 0.120292
R1870 dvdd.n165 dvdd.n99 0.120292
R1871 dvdd.n166 dvdd.n165 0.120292
R1872 dvdd.n167 dvdd.n166 0.120292
R1873 dvdd.n167 dvdd.n95 0.120292
R1874 dvdd.n171 dvdd.n95 0.120292
R1875 dvdd.n172 dvdd.n171 0.120292
R1876 dvdd.n173 dvdd.n172 0.120292
R1877 dvdd.n173 dvdd.n91 0.120292
R1878 dvdd.n177 dvdd.n91 0.120292
R1879 dvdd.n178 dvdd.n177 0.120292
R1880 dvdd.n179 dvdd.n178 0.120292
R1881 dvdd.n179 dvdd.n87 0.120292
R1882 dvdd.n184 dvdd.n87 0.120292
R1883 dvdd.n185 dvdd.n184 0.120292
R1884 dvdd.n186 dvdd.n185 0.120292
R1885 dvdd.n186 dvdd.n85 0.120292
R1886 dvdd.n190 dvdd.n85 0.120292
R1887 dvdd.n191 dvdd.n190 0.120292
R1888 dvdd.n192 dvdd.n191 0.120292
R1889 dvdd.n192 dvdd.n81 0.120292
R1890 dvdd.n196 dvdd.n81 0.120292
R1891 dvdd.n198 dvdd.n78 0.120292
R1892 dvdd.n203 dvdd.n78 0.120292
R1893 dvdd.n204 dvdd.n203 0.120292
R1894 dvdd.n205 dvdd.n204 0.120292
R1895 dvdd.n205 dvdd.n74 0.120292
R1896 dvdd.n209 dvdd.n74 0.120292
R1897 dvdd.n210 dvdd.n209 0.120292
R1898 dvdd.n211 dvdd.n210 0.120292
R1899 dvdd.n211 dvdd.n70 0.120292
R1900 dvdd.n215 dvdd.n70 0.120292
R1901 dvdd.n216 dvdd.n215 0.120292
R1902 dvdd.n217 dvdd.n216 0.120292
R1903 dvdd.n217 dvdd.n66 0.120292
R1904 dvdd.n222 dvdd.n66 0.120292
R1905 dvdd.n223 dvdd.n222 0.120292
R1906 dvdd.n224 dvdd.n223 0.120292
R1907 dvdd.n224 dvdd.n64 0.120292
R1908 dvdd.n228 dvdd.n64 0.120292
R1909 dvdd.n229 dvdd.n228 0.120292
R1910 dvdd.n230 dvdd.n229 0.120292
R1911 dvdd.n230 dvdd.n60 0.120292
R1912 dvdd.n234 dvdd.n60 0.120292
R1913 dvdd.n237 dvdd.n236 0.120292
R1914 dvdd.n241 dvdd.n57 0.120292
R1915 dvdd.n242 dvdd.n241 0.120292
R1916 dvdd.n277 dvdd.n276 0.109494
R1917 dvdd.n15 dvdd.n14 0.109053
R1918 dvdd.n268 dvdd.n244 0.107271
R1919 dvdd.n14 dvdd 0.0983618
R1920 dvdd dvdd.n262 0.0981562
R1921 dvdd.n251 dvdd 0.0968542
R1922 dvdd.n281 dvdd.n280 0.0944312
R1923 dvdd.n278 dvdd.n277 0.0856755
R1924 dvdd.n279 dvdd.n278 0.0856755
R1925 dvdd.n237 dvdd 0.0812292
R1926 dvdd dvdd.n6 0.0803611
R1927 dvdd.n280 dvdd.n279 0.0777774
R1928 dvdd.n14 dvdd.n7 0.070241
R1929 dvdd.n25 dvdd.n24 0.0685285
R1930 dvdd.n268 dvdd 0.063
R1931 dvdd.n264 dvdd 0.0603958
R1932 dvdd dvdd.n263 0.0603958
R1933 dvdd.n248 dvdd 0.0603958
R1934 dvdd.n120 dvdd 0.0603958
R1935 dvdd.n159 dvdd 0.0603958
R1936 dvdd.n160 dvdd 0.0603958
R1937 dvdd.n197 dvdd 0.0603958
R1938 dvdd.n198 dvdd 0.0603958
R1939 dvdd.n235 dvdd 0.0603958
R1940 dvdd.n236 dvdd 0.0603958
R1941 dvdd.n269 dvdd 0.0603958
R1942 dvdd dvdd.n13 0.0595278
R1943 dvdd.n21 dvdd.n16 0.0535523
R1944 dvdd.n12 dvdd 0.0508472
R1945 dvdd.n291 dvdd.n290 0.0456945
R1946 dvdd.n39 dvdd.n38 0.0456858
R1947 dvdd.n20 dvdd 0.0405
R1948 dvdd dvdd.n57 0.0395625
R1949 dvdd dvdd.n297 0.0385435
R1950 dvdd dvdd.n247 0.0382604
R1951 dvdd.n39 dvdd.n0 0.0379437
R1952 dvdd.n21 dvdd 0.0339302
R1953 dvdd.n13 dvdd.n12 0.0334861
R1954 dvdd.n275 dvdd 0.03175
R1955 dvdd dvdd.n159 0.03175
R1956 dvdd dvdd.n197 0.03175
R1957 dvdd dvdd.n235 0.03175
R1958 dvdd.n269 dvdd 0.03175
R1959 dvdd.n24 dvdd.n16 0.0300191
R1960 dvdd.n248 dvdd 0.0239375
R1961 dvdd.n49 dvdd.n0 0.0233041
R1962 dvdd.n263 dvdd 0.0226354
R1963 dvdd dvdd.n158 0.0226354
R1964 dvdd dvdd.n196 0.0226354
R1965 dvdd dvdd.n234 0.0226354
R1966 dvdd dvdd.n242 0.0226354
R1967 dvdd.n299 dvdd.n298 0.0219531
R1968 dvdd.n15 dvdd 0.0210592
R1969 dvdd.n20 dvdd.n19 0.0205
R1970 dvdd.n48 dvdd.n1 0.0182365
R1971 dvdd.n25 dvdd 0.0179419
R1972 dvdd.n49 dvdd.n48 0.0151396
R1973 dvdd.n290 dvdd.n281 0.0150881
R1974 dvdd dvdd.n20 0.0121279
R1975 dvdd.n299 dvdd.n281 0.00936728
R1976 dvdd.n268 dvdd.n243 0.0083125
R1977 dvdd.n277 dvdd.t178 0.0083125
R1978 dvdd.n278 dvdd.t177 0.0083125
R1979 dvdd.n279 dvdd.t176 0.0083125
R1980 dvdd.n50 dvdd.t175 0.0083125
R1981 dvdd.n298 dvdd 0.00765103
R1982 dvdd.n280 dvdd.n50 0.00754239
R1983 dvdd.n1 dvdd 0.00176689
R1984 dvdd.n299 dvdd 0.001125
R1985 a_20376_n2791.n1 a_20376_n2791.n0 926.024
R1986 a_20376_n2791.n1 a_20376_n2791.t2 82.0838
R1987 a_20376_n2791.n0 a_20376_n2791.t3 63.3338
R1988 a_20376_n2791.t0 a_20376_n2791.n1 63.3219
R1989 a_20376_n2791.n0 a_20376_n2791.t1 29.7268
R1990 a_19955_n2241.n1 a_19955_n2241.t7 530.01
R1991 a_19955_n2241.t0 a_19955_n2241.n5 421.021
R1992 a_19955_n2241.n0 a_19955_n2241.t2 337.142
R1993 a_19955_n2241.n3 a_19955_n2241.t1 280.223
R1994 a_19955_n2241.n4 a_19955_n2241.t3 263.173
R1995 a_19955_n2241.n4 a_19955_n2241.t5 227.826
R1996 a_19955_n2241.n0 a_19955_n2241.t4 199.762
R1997 a_19955_n2241.n2 a_19955_n2241.n1 170.81
R1998 a_19955_n2241.n2 a_19955_n2241.n0 167.321
R1999 a_19955_n2241.n5 a_19955_n2241.n4 152
R2000 a_19955_n2241.n1 a_19955_n2241.t6 141.923
R2001 a_19955_n2241.n3 a_19955_n2241.n2 10.8376
R2002 a_19955_n2241.n5 a_19955_n2241.n3 2.50485
R2003 a_20689_n2273.n3 a_20689_n2273.n2 647.119
R2004 a_20689_n2273.n1 a_20689_n2273.t4 350.253
R2005 a_20689_n2273.n2 a_20689_n2273.n0 260.339
R2006 a_20689_n2273.n2 a_20689_n2273.n1 246.119
R2007 a_20689_n2273.n1 a_20689_n2273.t5 189.588
R2008 a_20689_n2273.n3 a_20689_n2273.t2 89.1195
R2009 a_20689_n2273.n0 a_20689_n2273.t1 63.3338
R2010 a_20689_n2273.t3 a_20689_n2273.n3 41.0422
R2011 a_20689_n2273.n0 a_20689_n2273.t0 31.9797
R2012 a_21036_n1869.n3 a_21036_n1869.n2 636.953
R2013 a_21036_n1869.n1 a_21036_n1869.t5 366.856
R2014 a_21036_n1869.n2 a_21036_n1869.n0 300.2
R2015 a_21036_n1869.n2 a_21036_n1869.n1 225.036
R2016 a_21036_n1869.n1 a_21036_n1869.t4 174.056
R2017 a_21036_n1869.n0 a_21036_n1869.t0 70.0005
R2018 a_21036_n1869.n3 a_21036_n1869.t2 68.0124
R2019 a_21036_n1869.t1 a_21036_n1869.n3 63.3219
R2020 a_21036_n1869.n0 a_21036_n1869.t3 61.6672
R2021 a_10620_n8338.t0 a_10620_n8338.t1 83.9243
R2022 a_24220_n8172.t0 a_24220_n8172.t1 83.56
R2023 a_16620_n2791.n3 a_16620_n2791.n2 636.953
R2024 a_16620_n2791.n1 a_16620_n2791.t4 366.856
R2025 a_16620_n2791.n2 a_16620_n2791.n0 300.2
R2026 a_16620_n2791.n2 a_16620_n2791.n1 225.036
R2027 a_16620_n2791.n1 a_16620_n2791.t5 174.056
R2028 a_16620_n2791.n0 a_16620_n2791.t3 70.0005
R2029 a_16620_n2791.n3 a_16620_n2791.t2 68.0124
R2030 a_16620_n2791.t0 a_16620_n2791.n3 63.3219
R2031 a_16620_n2791.n0 a_16620_n2791.t1 61.6672
R2032 a_16974_n2791.t0 a_16974_n2791.t1 87.1434
R2033 a_16795_n2817.n4 a_16795_n2817.n0 746.659
R2034 a_16795_n2817.n5 a_16795_n2817.t3 389.183
R2035 a_16795_n2817.n1 a_16795_n2817.t7 256.988
R2036 a_16795_n2817.n6 a_16795_n2817.n5 251.167
R2037 a_16795_n2817.t0 a_16795_n2817.n6 223.571
R2038 a_16795_n2817.n3 a_16795_n2817.t5 212.081
R2039 a_16795_n2817.n4 a_16795_n2817.n3 181.942
R2040 a_16795_n2817.n5 a_16795_n2817.t8 174.891
R2041 a_16795_n2817.n1 a_16795_n2817.t4 163.803
R2042 a_16795_n2817.n2 a_16795_n2817.t6 139.78
R2043 a_16795_n2817.n2 a_16795_n2817.n1 129.264
R2044 a_16795_n2817.n0 a_16795_n2817.t1 63.3219
R2045 a_16795_n2817.n0 a_16795_n2817.t2 63.3219
R2046 a_16795_n2817.n6 a_16795_n2817.n4 24.6993
R2047 a_16795_n2817.n3 a_16795_n2817.n2 22.6399
R2048 ena_ip.t1 ena_ip.n0 744.115
R2049 ena_ip ena_ip.t1 732.75
R2050 ena_ip.n15 ena_ip.t7 408.63
R2051 ena_ip.n11 ena_ip.t13 408.63
R2052 ena_ip.n7 ena_ip.t4 408.63
R2053 ena_ip.n12 ena_ip.t6 347.577
R2054 ena_ip.n8 ena_ip.t8 347.577
R2055 ena_ip.n4 ena_ip.t16 347.577
R2056 ena_ip.n2 ena_ip.t14 332.752
R2057 ena_ip.t14 ena_ip.n1 332.752
R2058 ena_ip.n2 ena_ip.t17 332.411
R2059 ena_ip.t17 ena_ip.n1 332.411
R2060 ena_ip.n16 ena_ip.t19 239.505
R2061 ena_ip ena_ip.t0 216.155
R2062 ena_ip.n12 ena_ip.t9 193.337
R2063 ena_ip.n8 ena_ip.t10 193.337
R2064 ena_ip.n4 ena_ip.t18 193.337
R2065 ena_ip.n16 ena_ip.t11 167.204
R2066 ena_ip ena_ip.n15 165.089
R2067 ena_ip ena_ip.n11 165.089
R2068 ena_ip ena_ip.n7 165.089
R2069 ena_ip ena_ip.n16 157.12
R2070 ena_ip.n13 ena_ip.n12 152
R2071 ena_ip.n9 ena_ip.n8 152
R2072 ena_ip.n5 ena_ip.n4 152
R2073 ena_ip.n15 ena_ip.t3 132.282
R2074 ena_ip.n11 ena_ip.t5 132.282
R2075 ena_ip.n7 ena_ip.t15 132.282
R2076 ena_ip ena_ip.t2 59.9857
R2077 ena_ip ena_ip.t12 59.0936
R2078 ena_ip.n0 ena_ip 57.4755
R2079 ena_ip ena_ip.n17 13.8078
R2080 ena_ip.n17 ena_ip 9.82907
R2081 ena_ip ena_ip.n6 9.3005
R2082 ena_ip ena_ip.n10 9.3005
R2083 ena_ip ena_ip.n14 9.3005
R2084 ena_ip ena_ip.n18 8.84514
R2085 ena_ip.n17 ena_ip 5.71479
R2086 ena_ip.n3 ena_ip.n1 5.53161
R2087 ena_ip.n13 ena_ip 4.67077
R2088 ena_ip.n9 ena_ip 4.67077
R2089 ena_ip.n5 ena_ip 4.67077
R2090 ena_ip.n3 ena_ip.n2 4.67076
R2091 ena_ip.n18 ena_ip 4.17561
R2092 ena_ip.n0 ena_ip 3.62625
R2093 ena_ip ena_ip.n3 3.51723
R2094 ena_ip.n14 ena_ip 2.94104
R2095 ena_ip.n10 ena_ip 2.94104
R2096 ena_ip.n6 ena_ip 2.94104
R2097 ena_ip.n18 ena_ip 2.93705
R2098 ena_ip.n14 ena_ip.n13 2.76807
R2099 ena_ip.n10 ena_ip.n9 2.76807
R2100 ena_ip.n6 ena_ip.n5 2.76807
R2101 x3.in_b.n1 x3.in_b.n0 3.2348
R2102 x3.in_b.n1 x3.in_b.t3 166.376
R2103 x3.in_b.n1 x3.in_b.t2 166.207
R2104 x3.in_b.n0 x3.in_b.t0 228.429
R2105 x3.in_b.n0 x3.in_b.t1 83.9309
R2106 a_21211_n1943.n6 a_21211_n1943.n5 746.659
R2107 a_21211_n1943.n0 a_21211_n1943.t6 389.183
R2108 a_21211_n1943.n2 a_21211_n1943.t4 256.988
R2109 a_21211_n1943.n1 a_21211_n1943.n0 251.167
R2110 a_21211_n1943.n1 a_21211_n1943.t1 223.571
R2111 a_21211_n1943.n4 a_21211_n1943.t7 212.081
R2112 a_21211_n1943.n5 a_21211_n1943.n4 181.942
R2113 a_21211_n1943.n0 a_21211_n1943.t8 174.891
R2114 a_21211_n1943.n2 a_21211_n1943.t5 163.803
R2115 a_21211_n1943.n3 a_21211_n1943.t3 139.78
R2116 a_21211_n1943.n3 a_21211_n1943.n2 129.264
R2117 a_21211_n1943.t0 a_21211_n1943.n6 63.3219
R2118 a_21211_n1943.n6 a_21211_n1943.t2 63.3219
R2119 a_21211_n1943.n5 a_21211_n1943.n1 24.6993
R2120 a_21211_n1943.n4 a_21211_n1943.n3 22.6399
R2121 a_17913_n2791.t1 a_17913_n2791.n3 370.026
R2122 a_17913_n2791.n0 a_17913_n2791.t2 351.356
R2123 a_17913_n2791.n1 a_17913_n2791.t5 334.717
R2124 a_17913_n2791.n3 a_17913_n2791.t0 325.971
R2125 a_17913_n2791.n1 a_17913_n2791.t4 309.935
R2126 a_17913_n2791.n0 a_17913_n2791.t3 305.683
R2127 a_17913_n2791.n2 a_17913_n2791.n0 16.879
R2128 a_17913_n2791.n3 a_17913_n2791.n2 10.8867
R2129 a_17913_n2791.n2 a_17913_n2791.n1 9.3005
R2130 a_18481_n2549.n3 a_18481_n2549.n2 647.119
R2131 a_18481_n2549.n1 a_18481_n2549.t4 350.253
R2132 a_18481_n2549.n2 a_18481_n2549.n0 260.339
R2133 a_18481_n2549.n2 a_18481_n2549.n1 246.119
R2134 a_18481_n2549.n1 a_18481_n2549.t5 189.588
R2135 a_18481_n2549.n3 a_18481_n2549.t3 89.1195
R2136 a_18481_n2549.n0 a_18481_n2549.t1 63.3338
R2137 a_18481_n2549.t0 a_18481_n2549.n3 41.0422
R2138 a_18481_n2549.n0 a_18481_n2549.t2 31.9797
R2139 a_18828_n2791.n3 a_18828_n2791.n2 636.953
R2140 a_18828_n2791.n1 a_18828_n2791.t4 366.856
R2141 a_18828_n2791.n2 a_18828_n2791.n0 300.2
R2142 a_18828_n2791.n2 a_18828_n2791.n1 225.036
R2143 a_18828_n2791.n1 a_18828_n2791.t5 174.056
R2144 a_18828_n2791.n0 a_18828_n2791.t1 70.0005
R2145 a_18828_n2791.n3 a_18828_n2791.t3 68.0124
R2146 a_18828_n2791.t2 a_18828_n2791.n3 63.3219
R2147 a_18828_n2791.n0 a_18828_n2791.t0 61.6672
R2148 a_2130_n19848.t0 a_2130_n19848.t1 82.0028
R2149 a_24530_n20014.t0 a_24530_n20014.t1 81.9478
R2150 icnode.t0 icnode.t1 84.1171
R2151 a_11526_n12394.t0 a_11526_n12394.t1 78.7148
R2152 vbreg.n21 vbreg.t5 244.944
R2153 vbreg.n49 vbreg.n2 202.542
R2154 vbreg.n40 vbreg.n10 201.036
R2155 vbreg.n33 vbreg.n7 200.282
R2156 vbreg.n20 vbreg.n21 0.962138
R2157 vbreg.n35 vbreg.n10 179.201
R2158 vbreg.n2 vbreg.n24 178.447
R2159 vbreg.n35 vbreg.n7 176.941
R2160 vbreg.n42 vbreg.n24 160.376
R2161 vbreg.n35 vbreg.n19 116.609
R2162 vbreg.n35 vbreg.n15 116.609
R2163 vbreg.n30 vbreg.n10 116.609
R2164 vbreg.n17 vbreg.n10 116.609
R2165 vbreg.n44 vbreg.n24 116.609
R2166 vbreg.n56 vbreg.n24 116.609
R2167 vbreg.n53 vbreg.n2 116.609
R2168 vbreg.n2 vbreg.n25 116.609
R2169 vbreg.n18 vbreg.n7 116.609
R2170 vbreg.n16 vbreg.n7 116.609
R2171 vbreg.n42 vbreg.n26 115.005
R2172 vbreg.n42 vbreg.n40 110.683
R2173 vbreg.t13 vbreg.n31 86.3125
R2174 vbreg.n14 vbreg.t10 88.4838
R2175 vbreg.n18 vbreg.t14 86.3125
R2176 vbreg.t12 vbreg.n16 86.3125
R2177 vbreg.t23 vbreg.n12 88.4979
R2178 vbreg.n51 vbreg.t25 86.3125
R2179 vbreg.t17 vbreg.n38 86.3125
R2180 vbreg.n28 vbreg.t18 86.3125
R2181 vbreg.n15 vbreg.t9 86.3125
R2182 vbreg.n19 vbreg.t11 86.3125
R2183 vbreg.n37 vbreg.t15 86.3125
R2184 vbreg.n29 vbreg.t16 86.3125
R2185 vbreg.n57 vbreg.t6 86.3125
R2186 vbreg.n43 vbreg.t20 86.3125
R2187 vbreg.n55 vbreg.t19 86.3125
R2188 vbreg.n54 vbreg.t22 86.3125
R2189 vbreg.n47 vbreg.t21 86.3125
R2190 vbreg.n52 vbreg.t24 86.3125
R2191 vbreg.n16 vbreg.n14 2.64048
R2192 vbreg.n38 vbreg.n37 72.5338
R2193 vbreg.n12 vbreg.n47 2.18593
R2194 vbreg.n18 vbreg.n31 72.5338
R2195 vbreg.n29 vbreg.n28 72.5338
R2196 vbreg.n52 vbreg.n51 72.5338
R2197 vbreg.n15 vbreg.n17 71.7809
R2198 vbreg.n57 vbreg.n56 71.7809
R2199 vbreg.n19 vbreg.n30 71.7809
R2200 vbreg.n28 vbreg.n26 71.7809
R2201 vbreg.n44 vbreg.n43 71.7809
R2202 vbreg.n16 vbreg.n15 71.5299
R2203 vbreg.n13 vbreg.n18 2.62088
R2204 vbreg.n55 vbreg.n25 71.2789
R2205 vbreg.n54 vbreg.n53 71.2789
R2206 vbreg.n38 vbreg.n23 60.7378
R2207 vbreg.n11 vbreg.t7 60.1061
R2208 vbreg.n32 vbreg.t13 55.9125
R2209 vbreg.n32 vbreg.t10 55.9125
R2210 vbreg.t14 vbreg.n34 55.9125
R2211 vbreg.n34 vbreg.t12 55.9125
R2212 vbreg.n48 vbreg.t23 55.9125
R2213 vbreg.n48 vbreg.t25 55.9125
R2214 vbreg.n39 vbreg.t17 55.9125
R2215 vbreg.n39 vbreg.t18 55.9125
R2216 vbreg.t9 vbreg.n36 55.9125
R2217 vbreg.n36 vbreg.t11 55.9125
R2218 vbreg.n27 vbreg.t15 55.9125
R2219 vbreg.t16 vbreg.n27 55.9125
R2220 vbreg.n41 vbreg.t6 55.9125
R2221 vbreg.n41 vbreg.t20 55.9125
R2222 vbreg.n45 vbreg.t19 55.9125
R2223 vbreg.t22 vbreg.n45 55.9125
R2224 vbreg.t21 vbreg.n46 55.9125
R2225 vbreg.n46 vbreg.t24 55.9125
R2226 vbreg.n33 vbreg.n32 30.4005
R2227 vbreg.n49 vbreg.n48 30.4005
R2228 vbreg.n36 vbreg.n35 30.4005
R2229 vbreg.n27 vbreg.n10 30.4005
R2230 vbreg.n40 vbreg.n39 30.4005
R2231 vbreg.n42 vbreg.n41 30.4005
R2232 vbreg.n45 vbreg.n24 30.4005
R2233 vbreg.n46 vbreg.n2 30.4005
R2234 vbreg.n34 vbreg.n7 30.4005
R2235 vbreg.n21 vbreg.t2 22.4019
R2236 vbreg.n22 vbreg.t0 21.1527
R2237 vbreg.n21 vbreg.t1 21.0621
R2238 vbreg.n42 vbreg.n11 2.00645
R2239 vbreg.n11 vbreg.n23 15.0573
R2240 vbreg.n57 vbreg.n23 11.7966
R2241 vbreg.n21 vbreg.n22 0.632464
R2242 vbreg.n40 vbreg.n3 3.01598
R2243 vbreg.n51 vbreg.n50 2.92951
R2244 vbreg.n4 vbreg.n31 2.92951
R2245 vbreg.n50 vbreg.n49 2.3255
R2246 vbreg.n0 vbreg.n2 2.3255
R2247 vbreg.n38 vbreg.n3 2.3255
R2248 vbreg.n55 vbreg.n3 2.3255
R2249 vbreg.n0 vbreg.n54 2.3255
R2250 vbreg.n52 vbreg.n0 2.3255
R2251 vbreg.n4 vbreg.n33 2.3255
R2252 vbreg.n5 vbreg.n7 2.3255
R2253 vbreg.n37 vbreg.n9 2.3255
R2254 vbreg.n9 vbreg.n10 2.3255
R2255 vbreg.n29 vbreg.n9 2.3255
R2256 vbreg.n28 vbreg.n8 2.3255
R2257 vbreg.n43 vbreg.n8 2.3255
R2258 vbreg.n3 vbreg.n57 2.3255
R2259 vbreg.n8 vbreg.n11 1.77359
R2260 vbreg.n3 vbreg.n20 1.69825
R2261 vbreg.n47 vbreg.n25 1.2554
R2262 vbreg.n53 vbreg.n52 1.2554
R2263 vbreg.n20 vbreg.t8 21.8362
R2264 vbreg.n21 vbreg.t4 21.6418
R2265 vbreg.n22 vbreg.t3 21.6076
R2266 vbreg.n19 vbreg.n13 2.62088
R2267 vbreg.n9 vbreg.n15 2.82746
R2268 vbreg.n6 vbreg.n5 0.489702
R2269 vbreg.n9 vbreg.n6 0.553315
R2270 vbreg.n1 vbreg.n0 0.420519
R2271 vbreg.n9 vbreg.n8 1.22324
R2272 vbreg.n6 vbreg.n35 2.715
R2273 vbreg.n12 vbreg.n0 1.45199
R2274 vbreg.n50 vbreg.n0 1.13148
R2275 vbreg.n5 vbreg.n4 1.12454
R2276 vbreg.n1 vbreg.n3 0.237615
R2277 vbreg.n5 vbreg.n13 0.795018
R2278 vbreg.n14 vbreg.n5 0.776083
R2279 vbreg.n3 vbreg.n11 0.753999
R2280 vbreg.n37 vbreg.n17 0.753441
R2281 vbreg.n56 vbreg.n55 0.753441
R2282 vbreg.n30 vbreg.n29 0.753441
R2283 vbreg.n43 vbreg.n26 0.753441
R2284 vbreg.n54 vbreg.n44 0.753441
R2285 vbreg.n1 vbreg.n24 2.61619
R2286 a_15000_n2791.n2 a_15000_n2791.n1 682.193
R2287 a_15000_n2791.n0 a_15000_n2791.t4 279.142
R2288 a_15000_n2791.n1 a_15000_n2791.t1 250.526
R2289 a_15000_n2791.n0 a_15000_n2791.t3 145.958
R2290 a_15000_n2791.n1 a_15000_n2791.n0 118.642
R2291 a_15000_n2791.n2 a_15000_n2791.t2 70.3576
R2292 a_15000_n2791.t0 a_15000_n2791.n2 65.6672
R2293 x7.x2.x2.CLK x7.x2.x2.CLK.t0 721.571
R2294 x7.x2.x2.CLK.n2 x7.x2.x2.CLK.t0 707.66
R2295 x7.x2.x2.CLK.n0 x7.x2.x2.CLK.t2 294.557
R2296 x7.x2.x2.CLK.n1 x7.x2.x2.CLK.t1 271.777
R2297 x7.x2.x2.CLK.n0 x7.x2.x2.CLK.t3 211.01
R2298 x7.x2.x2.CLK x7.x2.x2.CLK.n0 152
R2299 x7.x2.x2.CLK.n2 x7.x2.x2.CLK.n1 38.2982
R2300 x7.x2.x2.CLK.n1 x7.x2.x2.CLK 32.5125
R2301 x7.x2.x2.CLK x7.x2.x2.CLK.n2 3.76521
R2302 x7.x1.Qb2.n4 x7.x1.Qb2.t1 372.361
R2303 x7.x1.Qb2.n2 x7.x1.Qb2.t2 333.651
R2304 x7.x1.Qb2.n2 x7.x1.Qb2.t5 297.233
R2305 x7.x1.Qb2.n0 x7.x1.Qb2.t3 294.557
R2306 x7.x1.Qb2.n5 x7.x1.Qb2.t0 231.921
R2307 x7.x1.Qb2.n0 x7.x1.Qb2.t4 211.01
R2308 x7.x1.Qb2 x7.x1.Qb2.n2 195.701
R2309 x7.x1.Qb2.n1 x7.x1.Qb2.n0 152
R2310 x7.x1.Qb2.n5 x7.x1.Qb2.n1 41.5091
R2311 x7.x1.Qb2.n5 x7.x1.Qb2.n4 18.1966
R2312 x7.x1.Qb2.n4 x7.x1.Qb2.n3 9.36092
R2313 x7.x1.Qb2.n3 x7.x1.Qb2 6.49269
R2314 x7.x1.Qb2.n1 x7.x1.Qb2 4.20621
R2315 x7.x1.Qb2.n3 x7.x1.Qb2 3.52967
R2316 x7.x1.Qb2 x7.x1.Qb2.n5 2.5605
R2317 a_18168_n1881.n1 a_18168_n1881.n0 926.024
R2318 a_18168_n1881.n1 a_18168_n1881.t2 82.0838
R2319 a_18168_n1881.n0 a_18168_n1881.t3 63.3338
R2320 a_18168_n1881.t0 a_18168_n1881.n1 63.3219
R2321 a_18168_n1881.n0 a_18168_n1881.t1 29.7268
R2322 vbp vbp.t9 165.465
R2323 vbp.n8 vbp 165.078
R2324 vbp.n2 vbp.t13 164.613
R2325 vbp.n4 vbp 163.965
R2326 vbp.n1 vbp 109.079
R2327 vbp vbp.t11 64.4412
R2328 vbp vbp.n0 83.6272
R2329 vbp.n0 vbp 83.2005
R2330 vbp.t0 vbp 62.2125
R2331 vbp.t7 vbp 62.2125
R2332 vbp vbp.t5 62.2125
R2333 vbp vbp.t10 62.2125
R2334 vbp.t15 vbp 65.3588
R2335 vbp.t12 vbp 62.2125
R2336 vbp.n0 vbp.t2 62.2125
R2337 vbp.n2 vbp.t6 62.2125
R2338 vbp vbp.t14 62.2125
R2339 vbp vbp.t4 62.2125
R2340 vbp vbp.t1 62.2125
R2341 vbp.t8 vbp 62.2125
R2342 vbp.t3 vbp 65.3497
R2343 vbp.n0 vbp 37.5472
R2344 vbp.n10 vbp.t0 31.8125
R2345 vbp.n10 vbp.t7 31.8125
R2346 vbp.n7 vbp.t5 31.8125
R2347 vbp.t10 vbp.n7 31.8125
R2348 vbp.n8 vbp.t15 31.8125
R2349 vbp.t9 vbp.n8 31.8125
R2350 vbp.n9 vbp.t12 31.8125
R2351 vbp.t2 vbp.n9 31.8125
R2352 vbp.n3 vbp.t6 31.8125
R2353 vbp.t11 vbp.n3 31.8125
R2354 vbp.t14 vbp.n5 31.8125
R2355 vbp.n5 vbp.t4 31.8125
R2356 vbp.t1 vbp.n6 31.8125
R2357 vbp.n6 vbp.t8 31.8125
R2358 vbp.n4 vbp.t3 31.8125
R2359 vbp.t13 vbp.n4 31.8125
R2360 vbp.n9 vbp 30.4005
R2361 vbp.n7 vbp 30.4005
R2362 vbp.n5 vbp.n1 30.4005
R2363 vbp.n3 vbp 30.4005
R2364 vbp.n6 vbp 30.4005
R2365 vbp vbp.n10 30.4005
R2366 vbp.n2 vbp 18.4815
R2367 vbp vbp.n1 15.0659
R2368 vbp vbp.n0 10.3663
R2369 dvdd_ip.n75 dvdd_ip.n54 36575
R2370 dvdd_ip.n76 dvdd_ip.n75 36575
R2371 dvdd_ip.n77 dvdd_ip.n76 36575
R2372 dvdd_ip.n77 dvdd_ip.n54 36575
R2373 dvdd_ip.n74 dvdd_ip.n52 18251.4
R2374 dvdd_ip.n74 dvdd_ip.n53 18251.4
R2375 dvdd_ip.n78 dvdd_ip.n53 18251.4
R2376 dvdd_ip.n78 dvdd_ip.n52 18251.4
R2377 dvdd_ip.n109 dvdd_ip.n33 10440
R2378 dvdd_ip.n111 dvdd_ip.n33 10440
R2379 dvdd_ip.n111 dvdd_ip.n34 10440
R2380 dvdd_ip.n109 dvdd_ip.n34 10440
R2381 dvdd_ip.n59 dvdd_ip.n51 4516.33
R2382 dvdd_ip.n79 dvdd_ip.n51 4243.24
R2383 dvdd_ip.n62 dvdd_ip.n58 4030.59
R2384 dvdd_ip.n65 dvdd_ip.n57 4030.59
R2385 dvdd_ip.n107 dvdd_ip.n42 4030.59
R2386 dvdd_ip.n104 dvdd_ip.n43 4030.59
R2387 dvdd_ip.n55 dvdd_ip.n4 3741.35
R2388 dvdd_ip.n73 dvdd_ip.n55 3618.82
R2389 dvdd_ip.n100 dvdd_ip.n96 3190.03
R2390 dvdd_ip.n100 dvdd_ip.n97 3190.03
R2391 dvdd_ip.n98 dvdd_ip.n97 3190.03
R2392 dvdd_ip.n98 dvdd_ip.n96 3190.03
R2393 dvdd_ip.n84 dvdd_ip.n16 2795.29
R2394 dvdd_ip.n81 dvdd_ip.n50 2795.29
R2395 dvdd_ip.n87 dvdd_ip.n86 2417.65
R2396 dvdd_ip.n89 dvdd_ip.n86 2417.65
R2397 dvdd_ip.n89 dvdd_ip.n85 2417.65
R2398 dvdd_ip.n87 dvdd_ip.n85 2417.65
R2399 dvdd_ip.n105 dvdd_ip.n42 1199.77
R2400 dvdd_ip.n106 dvdd_ip.n43 1199.77
R2401 dvdd_ip.n82 dvdd_ip.n16 703.912
R2402 dvdd_ip.n83 dvdd_ip.n50 703.912
R2403 dvdd_ip.n60 dvdd_ip.n59 654.165
R2404 dvdd_ip.n46 dvdd_ip.t37 642.13
R2405 dvdd_ip.n67 dvdd_ip.t46 642.13
R2406 dvdd_ip.n103 dvdd_ip.t42 642.13
R2407 dvdd_ip.n10 dvdd_ip.n47 594.953
R2408 dvdd_ip.n10 dvdd_ip.n48 594.301
R2409 dvdd_ip.n61 dvdd_ip.n56 429.93
R2410 dvdd_ip.n61 dvdd_ip.n60 429.93
R2411 dvdd_ip.t19 dvdd_ip.t5 397.805
R2412 dvdd_ip.t13 dvdd_ip.t19 397.805
R2413 dvdd_ip.t15 dvdd_ip.t13 397.805
R2414 dvdd_ip.t8 dvdd_ip.t23 397.805
R2415 dvdd_ip.t17 dvdd_ip.t8 397.805
R2416 dvdd_ip.t10 dvdd_ip.t17 397.805
R2417 dvdd_ip.n66 dvdd_ip.n56 340.42
R2418 dvdd_ip.t0 dvdd_ip.n85 327.8
R2419 dvdd_ip.t35 dvdd_ip.n86 327.8
R2420 dvdd_ip.t54 dvdd_ip.t52 312.123
R2421 dvdd_ip.t38 dvdd_ip.t49 312.123
R2422 dvdd_ip.t52 dvdd_ip.n96 259.716
R2423 dvdd_ip.t49 dvdd_ip.n97 259.716
R2424 dvdd_ip.t5 dvdd_ip.n109 250.107
R2425 dvdd_ip.n111 dvdd_ip.t10 250.107
R2426 dvdd_ip.n101 dvdd_ip.n1 221.308
R2427 dvdd_ip.n110 dvdd_ip.t15 198.903
R2428 dvdd_ip.t23 dvdd_ip.n110 198.903
R2429 dvdd_ip.n88 dvdd_ip.t0 159.988
R2430 dvdd_ip.n88 dvdd_ip.t35 159.988
R2431 dvdd_ip.n99 dvdd_ip.t54 156.062
R2432 dvdd_ip.n99 dvdd_ip.t38 156.062
R2433 dvdd_ip.n21 dvdd_ip.n30 146.071
R2434 dvdd_ip.n108 dvdd_ip.n39 138.667
R2435 dvdd_ip.n27 dvdd_ip.t24 126.082
R2436 dvdd_ip.n31 dvdd_ip.t18 115.43
R2437 dvdd_ip.n28 dvdd_ip.t27 115.43
R2438 dvdd_ip.n35 dvdd_ip.t28 115.43
R2439 dvdd_ip.n37 dvdd_ip.t20 115.43
R2440 dvdd_ip.n0 dvdd_ip.t14 113.624
R2441 dvdd_ip.n3 dvdd_ip.t32 113.624
R2442 dvdd_ip.n18 dvdd_ip.t29 113.624
R2443 dvdd_ip.n0 dvdd_ip.t26 113.501
R2444 dvdd_ip.n3 dvdd_ip.t16 113.501
R2445 dvdd_ip.n32 dvdd_ip.t31 111.784
R2446 dvdd_ip.n31 dvdd_ip.t30 111.784
R2447 dvdd_ip.n29 dvdd_ip.t12 111.784
R2448 dvdd_ip.n28 dvdd_ip.t11 111.784
R2449 dvdd_ip.n35 dvdd_ip.t22 111.784
R2450 dvdd_ip.n36 dvdd_ip.t21 111.784
R2451 dvdd_ip.n37 dvdd_ip.t7 111.784
R2452 dvdd_ip.n38 dvdd_ip.t6 111.784
R2453 dvdd_ip.n19 dvdd_ip.t9 111.784
R2454 dvdd_ip.n19 dvdd_ip.t33 111.784
R2455 dvdd_ip.n27 dvdd_ip.t25 111.784
R2456 dvdd_ip.n64 dvdd_ip.n58 106.282
R2457 dvdd_ip.n63 dvdd_ip.n57 106.282
R2458 dvdd_ip.n24 dvdd_ip 1.37849
R2459 dvdd_ip.n94 dvdd_ip.n40 89.4643
R2460 dvdd_ip.n108 dvdd_ip.n26 64.1367
R2461 dvdd_ip.n25 dvdd_ip.t3 60.3236
R2462 dvdd_ip.n48 dvdd_ip.t1 57.1305
R2463 dvdd_ip.n48 dvdd_ip.t36 57.1305
R2464 dvdd_ip.n47 dvdd_ip.t4 57.1305
R2465 dvdd_ip.n47 dvdd_ip.t53 57.1305
R2466 dvdd_ip.n92 dvdd_ip.n44 55.1223
R2467 dvdd_ip.n20 dvdd_ip.n72 54.7105
R2468 dvdd_ip.n20 dvdd_ip.n69 54.7105
R2469 dvdd_ip.n20 dvdd_ip.n71 54.7085
R2470 dvdd_ip.n20 dvdd_ip.n70 54.7085
R2471 dvdd_ip.n20 dvdd_ip.n68 54.7085
R2472 dvdd_ip.n49 dvdd_ip.n46 53.6981
R2473 dvdd_ip.n66 dvdd_ip.n13 46.6446
R2474 dvdd_ip.n91 dvdd_ip.n43 46.2505
R2475 dvdd_ip.n102 dvdd_ip.n42 46.2505
R2476 dvdd_ip.n66 dvdd_ip.n65 46.2505
R2477 dvdd_ip.n62 dvdd_ip.n61 46.2505
R2478 dvdd_ip.n65 dvdd_ip.n64 44.5206
R2479 dvdd_ip.n63 dvdd_ip.n62 44.5206
R2480 dvdd_ip.n15 dvdd_ip.n23 0.871339
R2481 dvdd_ip.n102 dvdd_ip.n41 37.2058
R2482 dvdd_ip.n50 dvdd_ip.n14 37.0005
R2483 dvdd_ip.n4 dvdd_ip.n16 37.0005
R2484 dvdd_ip.n92 dvdd_ip.n45 33.5615
R2485 dvdd_ip.n7 dvdd_ip.n8 1.04644
R2486 dvdd_ip.n94 dvdd_ip.n41 31.3351
R2487 dvdd_ip.n85 dvdd_ip.n14 26.4291
R2488 dvdd_ip.n86 dvdd_ip.n45 26.4291
R2489 dvdd_ip.n104 dvdd_ip.n9 12.8793
R2490 dvdd_ip.n59 dvdd_ip.n13 23.3225
R2491 dvdd_ip.n5 dvdd_ip.n41 22.576
R2492 dvdd_ip.n87 dvdd_ip.n44 20.5561
R2493 dvdd_ip.n88 dvdd_ip.n87 20.5561
R2494 dvdd_ip.n90 dvdd_ip.n89 20.5561
R2495 dvdd_ip.n89 dvdd_ip.n88 20.5561
R2496 dvdd_ip.n90 dvdd_ip.n49 19.0763
R2497 dvdd_ip.n39 dvdd_ip.n1 18.9635
R2498 dvdd_ip.n46 dvdd_ip.n45 17.7956
R2499 dvdd_ip.n80 dvdd_ip.n4 17.833
R2500 dvdd_ip.n80 dvdd_ip.n17 17.8749
R2501 dvdd_ip.n36 dvdd_ip.n35 14.6565
R2502 dvdd_ip.n38 dvdd_ip.n37 14.6565
R2503 dvdd_ip.n29 dvdd_ip.n28 14.6565
R2504 dvdd_ip.n32 dvdd_ip.n31 14.6565
R2505 dvdd_ip.n23 dvdd_ip.n93 10.2385
R2506 dvdd_ip.n25 dvdd_ip.n11 0.591844
R2507 dvdd_ip.n17 dvdd_ip.n44 13.513
R2508 dvdd_ip.n81 dvdd_ip.n80 13.2148
R2509 dvdd_ip.n25 dvdd_ip.n84 13.2148
R2510 dvdd_ip.n96 dvdd_ip.n95 12.3338
R2511 dvdd_ip.n97 dvdd_ip.n39 12.3338
R2512 dvdd_ip.n21 dvdd_ip.n111 11.563
R2513 dvdd_ip.n102 dvdd_ip.n93 11.1792
R2514 dvdd_ip.n12 dvdd_ip.n6 1.8903
R2515 dvdd_ip.n15 dvdd_ip.n94 11.0012
R2516 dvdd_ip.n22 dvdd_ip.n30 139.684
R2517 dvdd_ip.n82 dvdd_ip.n81 9.84115
R2518 dvdd_ip.n84 dvdd_ip.n83 9.84115
R2519 dvdd_ip.n7 dvdd_ip.n46 9.4314
R2520 dvdd_ip dvdd_ip.n67 9.39134
R2521 dvdd_ip.n15 dvdd_ip.n103 9.30175
R2522 dvdd_ip.n22 dvdd_ip.n1 1.1019
R2523 dvdd_ip.n26 dvdd_ip.n40 8.03454
R2524 dvdd_ip.n33 dvdd_ip.n24 15.3109
R2525 dvdd_ip.n5 dvdd_ip.n107 7.4005
R2526 dvdd_ip.n57 dvdd_ip.n56 7.4005
R2527 dvdd_ip.n60 dvdd_ip.n58 7.4005
R2528 dvdd_ip.n9 dvdd_ip.n15 0.167749
R2529 dvdd_ip.n72 dvdd_ip.t50 7.14175
R2530 dvdd_ip.n72 dvdd_ip.t39 7.14175
R2531 dvdd_ip.n71 dvdd_ip.t43 7.14175
R2532 dvdd_ip.n71 dvdd_ip.t40 7.14175
R2533 dvdd_ip.n70 dvdd_ip.t34 7.14175
R2534 dvdd_ip.n70 dvdd_ip.t47 7.14175
R2535 dvdd_ip.n69 dvdd_ip.t55 7.14175
R2536 dvdd_ip.n69 dvdd_ip.t48 7.14175
R2537 dvdd_ip.n68 dvdd_ip.t44 7.14175
R2538 dvdd_ip.n68 dvdd_ip.t51 7.14175
R2539 dvdd_ip.n101 dvdd_ip.n100 6.37981
R2540 dvdd_ip.n100 dvdd_ip.n99 6.37981
R2541 dvdd_ip.n98 dvdd_ip.n40 6.37981
R2542 dvdd_ip.n99 dvdd_ip.n98 6.37981
R2543 dvdd_ip.n92 dvdd_ip.n91 5.51614
R2544 dvdd_ip.n105 dvdd_ip.n104 5.18874
R2545 dvdd_ip.n107 dvdd_ip.n106 5.18874
R2546 dvdd_ip.n12 dvdd_ip.n79 5.53168
R2547 dvdd_ip.n73 dvdd_ip.n13 4.95261
R2548 dvdd_ip.n108 dvdd_ip.n22 3.23758
R2549 dvdd_ip.n17 dvdd_ip.n6 0.738278
R2550 dvdd_ip.n6 dvdd_ip.n90 3.8204
R2551 dvdd_ip.n21 dvdd_ip 3.55088
R2552 dvdd_ip.t2 dvdd_ip.n82 3.32862
R2553 dvdd_ip.n83 dvdd_ip.t2 3.32862
R2554 dvdd_ip.n7 dvdd_ip.n92 3.14232
R2555 dvdd_ip.n1 dvdd_ip.n36 3.1045
R2556 dvdd_ip.n1 dvdd_ip.n38 3.1045
R2557 dvdd_ip.n21 dvdd_ip.n32 3.1045
R2558 dvdd_ip.n11 dvdd_ip.n6 0.0238734
R2559 dvdd_ip.n110 dvdd_ip.n33 2.76169
R2560 dvdd_ip.n34 dvdd_ip.n30 2.76169
R2561 dvdd_ip.n110 dvdd_ip.n34 2.76169
R2562 dvdd_ip.n91 dvdd_ip.n8 2.74244
R2563 dvdd_ip.n95 dvdd_ip.n15 2.32363
R2564 dvdd_ip.n106 dvdd_ip.t41 2.20373
R2565 dvdd_ip.t41 dvdd_ip.n105 2.20373
R2566 dvdd_ip.n74 dvdd_ip.n73 2.07915
R2567 dvdd_ip.n75 dvdd_ip.n74 2.07915
R2568 dvdd_ip.n79 dvdd_ip.n78 2.07915
R2569 dvdd_ip.n78 dvdd_ip.n77 2.07915
R2570 dvdd_ip.n8 dvdd_ip.n49 9.20625
R2571 dvdd_ip.n18 dvdd_ip.n27 1.71757
R2572 dvdd_ip.n1 dvdd_ip.n24 1.42317
R2573 dvdd_ip.n67 dvdd_ip.n66 1.51323
R2574 dvdd_ip.n23 dvdd_ip.n101 82.9703
R2575 dvdd_ip.n21 dvdd_ip.n29 3.23543
R2576 dvdd_ip.t45 dvdd_ip.n63 1.22055
R2577 dvdd_ip.n64 dvdd_ip.t45 1.22055
R2578 dvdd_ip.n7 dvdd_ip.n5 1.02666
R2579 dvdd_ip.n7 dvdd_ip.n6 0.868735
R2580 dvdd_ip.n103 dvdd_ip.n102 0.83013
R2581 dvdd_ip.n26 dvdd_ip.n15 0.810159
R2582 dvdd_ip.n55 dvdd_ip.n52 0.768135
R2583 dvdd_ip.n54 dvdd_ip.n52 0.768135
R2584 dvdd_ip.n53 dvdd_ip.n51 0.768135
R2585 dvdd_ip.n76 dvdd_ip.n53 0.768135
R2586 dvdd_ip dvdd_ip.n2 0.748986
R2587 dvdd_ip.n0 dvdd_ip.n3 0.726273
R2588 dvdd_ip.n95 dvdd_ip.n93 0.70655
R2589 dvdd_ip.n2 dvdd_ip.n18 0.67791
R2590 dvdd_ip.n6 dvdd_ip.n10 0.621489
R2591 dvdd_ip dvdd_ip.n20 0.569502
R2592 dvdd_ip.n109 dvdd_ip.n1 11.6172
R2593 dvdd_ip.n26 dvdd_ip.n1 1.64329
R2594 dvdd_ip.n13 dvdd_ip 0.563996
R2595 dvdd_ip.n9 dvdd_ip.n7 0.547509
R2596 dvdd_ip.n2 dvdd_ip.n19 0.721964
R2597 dvdd_ip.n6 dvdd_ip.t56 0.442304
R2598 dvdd_ip.n1 dvdd_ip.n0 0.719176
R2599 dvdd_ip.n11 dvdd_ip.n14 1.41519
R2600 dvdd_ip.n4 dvdd_ip.n12 1.39615
R2601 dvdd_ip.n0 dvdd_ip.n2 1.26452
R2602 tail.n2 tail.t3 113.688
R2603 tail tail.t4 113.688
R2604 tail tail.t6 113.624
R2605 tail.n0 tail.t2 113.562
R2606 tail.n0 tail.t7 113.562
R2607 tail.n1 tail.t5 113.562
R2608 tail.n1 tail.t0 113.562
R2609 tail tail.t1 113.501
R2610 tail.n2 tail.t8 113.438
R2611 tail tail.t9 113.438
R2612 tail tail.n3 53.5531
R2613 tail.n3 tail.t11 6.92425
R2614 tail.n3 tail.t10 6.92425
R2615 tail tail.n1 1.9055
R2616 tail.n1 tail.n0 1.13844
R2617 tail tail.n2 1.13636
R2618 a_16273_n2549.n3 a_16273_n2549.n2 647.119
R2619 a_16273_n2549.n1 a_16273_n2549.t4 350.253
R2620 a_16273_n2549.n2 a_16273_n2549.n0 260.339
R2621 a_16273_n2549.n2 a_16273_n2549.n1 246.119
R2622 a_16273_n2549.n1 a_16273_n2549.t5 189.588
R2623 a_16273_n2549.n3 a_16273_n2549.t1 89.1195
R2624 a_16273_n2549.n0 a_16273_n2549.t3 63.3338
R2625 a_16273_n2549.t0 a_16273_n2549.n3 41.0422
R2626 a_16273_n2549.n0 a_16273_n2549.t2 31.9797
R2627 a_16151_n2791.t0 a_16151_n2791.t1 198.571
R2628 a_16317_n2791.t0 a_16317_n2791.t1 60.0005
R2629 standby_b.n18 standby_b.t14 408.63
R2630 standby_b.n20 standby_b.t25 408.63
R2631 standby_b.n22 standby_b.t11 408.63
R2632 standby_b.n12 standby_b.t6 401.051
R2633 standby_b.t6 standby_b.n11 401.051
R2634 standby_b.t19 standby_b.n3 401.051
R2635 standby_b.n4 standby_b.t19 401.051
R2636 standby_b.n12 standby_b.t16 371.31
R2637 standby_b.t16 standby_b.n11 371.31
R2638 standby_b.t18 standby_b.n13 371.31
R2639 standby_b.n14 standby_b.t18 371.31
R2640 standby_b.t0 standby_b.n10 371.31
R2641 standby_b.n15 standby_b.t0 371.31
R2642 standby_b.n17 standby_b.t3 371.31
R2643 standby_b.t3 standby_b.n16 371.31
R2644 standby_b.n9 standby_b.t21 371.31
R2645 standby_b.t21 standby_b.n8 371.31
R2646 standby_b.t23 standby_b.n2 371.31
R2647 standby_b.n7 standby_b.t23 371.31
R2648 standby_b.t7 standby_b.n5 371.31
R2649 standby_b.n6 standby_b.t7 371.31
R2650 standby_b.n4 standby_b.t17 371.31
R2651 standby_b.t17 standby_b.n3 371.31
R2652 standby_b.n26 standby_b.t13 347.577
R2653 standby_b.n25 standby_b.t15 347.577
R2654 standby_b.n24 standby_b.t2 347.577
R2655 standby_b.n0 standby_b.t12 332.752
R2656 standby_b.t12 x4.in_b 332.752
R2657 standby_b.n0 standby_b.t4 332.411
R2658 standby_b.t4 x4.in_b 332.411
R2659 standby_b.n27 standby_b.t24 236.552
R2660 standby_b.n26 standby_b.t8 193.337
R2661 standby_b.n25 standby_b.t9 193.337
R2662 standby_b.n24 standby_b.t22 193.337
R2663 x7.x2.x4.RESET_B standby_b.n18 165.089
R2664 x7.x2.x4.RESET_B standby_b.n20 165.089
R2665 x7.x2.x4.RESET_B standby_b.n22 165.089
R2666 standby_b.n27 standby_b.t10 164.251
R2667 x7.x3.A1 standby_b.n27 154.47
R2668 x7.x2.x2.RESET_B standby_b.n26 152
R2669 x7.x2.x3.RESET_B standby_b.n25 152
R2670 x7.x2.x4.RESET_B standby_b.n24 152
R2671 standby_b.n18 standby_b.t1 132.282
R2672 standby_b.n20 standby_b.t5 132.282
R2673 standby_b.n22 standby_b.t20 132.282
R2674 standby_b.n6 standby_b.n3 29.7417
R2675 standby_b.n7 standby_b.n6 29.7417
R2676 standby_b.n8 standby_b.n7 29.7417
R2677 standby_b.n16 standby_b.n15 29.7417
R2678 standby_b.n15 standby_b.n14 29.7417
R2679 standby_b.n14 standby_b.n11 29.7417
R2680 standby_b.n5 standby_b.n4 29.7417
R2681 standby_b.n5 standby_b.n2 29.7417
R2682 standby_b.n9 standby_b.n2 29.7417
R2683 standby_b.n17 standby_b.n10 29.7417
R2684 standby_b.n13 standby_b.n10 29.7417
R2685 standby_b.n13 standby_b.n12 29.7417
R2686 standby_b.n8 standby_b.n1 17.6946
R2687 standby_b.n1 standby_b.n9 17.5064
R2688 standby_b.n19 x7.x2.x4.RESET_B 16.7098
R2689 standby_b.n1 x7.stby_b 15.0825
R2690 x7.x2.x2.RESET_B standby_b.n19 14.0185
R2691 x7.x2.x3.RESET_B standby_b.n21 14.0185
R2692 x7.x2.x4.RESET_B standby_b.n23 14.0185
R2693 x7.stby_b x7.x3.A1 13.8064
R2694 standby_b.n1 standby_b.n17 12.2358
R2695 standby_b.n16 standby_b.n1 12.0476
R2696 standby_b.n19 x7.x2.x2.RESET_B 11.4672
R2697 standby_b.n21 x7.x2.x3.RESET_B 11.4672
R2698 standby_b.n23 x7.x2.x4.RESET_B 11.4672
R2699 x4.in_b standby_b.n0 11.1417
R2700 x7.stby_b x7.x2.x4.RESET_B 10.5569
R2701 x4.in_b standby_b.n1 10.4718
R2702 standby_b.n23 x7.x2.x4.RESET_B 9.3005
R2703 x7.x2.x4.RESET_B x7.x2.x3.RESET_B 9.3005
R2704 standby_b.n21 x7.x2.x4.RESET_B 9.3005
R2705 x7.x2.x4.RESET_B x7.x2.x2.RESET_B 9.3005
R2706 a_9120_n9346.n1 a_9120_n9346.t3 649.659
R2707 a_9120_n9346.n0 a_9120_n9346.t1 227.685
R2708 a_9120_n9346.t4 a_9120_n9346.n2 44.6806
R2709 a_9120_n9346.n1 a_9120_n9346.t2 5.45407
R2710 a_9120_n9346.n0 a_9120_n9346.t0 5.07473
R2711 a_9120_n9346.n2 a_9120_n9346.n0 0.639781
R2712 a_9120_n9346.n2 a_9120_n9346.n1 0.0621233
R2713 a_24220_n9832.t0 a_24220_n9832.t1 83.56
R2714 a_16974_n1881.t0 a_16974_n1881.t1 87.1434
R2715 a_16795_n1943.n6 a_16795_n1943.n5 746.659
R2716 a_16795_n1943.n0 a_16795_n1943.t8 389.183
R2717 a_16795_n1943.n2 a_16795_n1943.t4 256.988
R2718 a_16795_n1943.n1 a_16795_n1943.n0 251.167
R2719 a_16795_n1943.n1 a_16795_n1943.t1 223.571
R2720 a_16795_n1943.n4 a_16795_n1943.t5 212.081
R2721 a_16795_n1943.n5 a_16795_n1943.n4 181.942
R2722 a_16795_n1943.n0 a_16795_n1943.t7 174.891
R2723 a_16795_n1943.n2 a_16795_n1943.t6 163.803
R2724 a_16795_n1943.n3 a_16795_n1943.t3 139.78
R2725 a_16795_n1943.n3 a_16795_n1943.n2 129.264
R2726 a_16795_n1943.t0 a_16795_n1943.n6 63.3219
R2727 a_16795_n1943.n6 a_16795_n1943.t2 63.3219
R2728 a_16795_n1943.n5 a_16795_n1943.n1 24.6993
R2729 a_16795_n1943.n4 a_16795_n1943.n3 22.6399
R2730 a_21775_n2247.t0 a_21775_n2247.n1 386.31
R2731 a_21775_n2247.n1 a_21775_n2247.t1 249.956
R2732 a_21775_n2247.n0 a_21775_n2247.t2 239.04
R2733 a_21775_n2247.n1 a_21775_n2247.n0 175.661
R2734 a_21775_n2247.n0 a_21775_n2247.t3 166.739
R2735 x7.ena_done_b.n8 x7.ena_done_b.t0 373.866
R2736 x7.ena_done_b.n6 x7.ena_done_b.t5 333.651
R2737 x7.ena_done_b.n6 x7.ena_done_b.t6 297.233
R2738 x7.ena_done_b x7.ena_done_b.t1 247.159
R2739 x7.ena_done_b.n0 x7.ena_done_b.t3 241.536
R2740 x7.ena_done_b.n2 x7.ena_done_b.t4 207.423
R2741 x7.ena_done_b.n3 x7.ena_done_b.t7 202.133
R2742 x7.ena_done_b x7.ena_done_b.n6 195.701
R2743 x7.ena_done_b.n0 x7.ena_done_b.t2 169.237
R2744 x7.ena_done_b.n5 x7.ena_done_b.n2 159.758
R2745 x7.ena_done_b.n1 x7.ena_done_b.n0 155.84
R2746 x7.ena_done_b.n4 x7.ena_done_b.n3 152
R2747 x7.ena_done_b.n3 x7.ena_done_b.n2 36.8275
R2748 x7.ena_done_b x7.ena_done_b.n8 16.6907
R2749 x7.ena_done_b.n7 x7.ena_done_b 15.8995
R2750 x7.ena_done_b.n7 x7.ena_done_b 15.6656
R2751 x7.ena_done_b x7.ena_done_b.n5 13.8109
R2752 x7.ena_done_b x7.ena_done_b.n1 11.2245
R2753 x7.ena_done_b.n5 x7.ena_done_b.n4 5.4308
R2754 x7.ena_done_b.n4 x7.ena_done_b 3.68535
R2755 x7.ena_done_b.n1 x7.ena_done_b 3.2005
R2756 x7.ena_done_b.n8 x7.ena_done_b.n7 3.1005
R2757 a_20121_n2241.t0 a_20121_n2241.n3 370.026
R2758 a_20121_n2241.n0 a_20121_n2241.t2 351.356
R2759 a_20121_n2241.n1 a_20121_n2241.t4 334.717
R2760 a_20121_n2241.n3 a_20121_n2241.t1 325.971
R2761 a_20121_n2241.n1 a_20121_n2241.t5 309.935
R2762 a_20121_n2241.n0 a_20121_n2241.t3 305.683
R2763 a_20121_n2241.n2 a_20121_n2241.n0 16.879
R2764 a_20121_n2241.n3 a_20121_n2241.n2 10.8867
R2765 a_20121_n2241.n2 a_20121_n2241.n1 9.3005
R2766 a_2130_n21176.t0 a_2130_n21176.t1 82.0028
R2767 a_24530_n21342.t0 a_24530_n21342.t1 81.9492
R2768 standby_33.n0 standby_33.t0 227.886
R2769 standby_33 standby_33.t3 216.05
R2770 standby_33.n0 standby_33.n1 25.0903
R2771 standby_33.n0 standby_33.t4 12.7763
R2772 standby_33.n1 standby_33.t2 5.5105
R2773 standby_33.n1 standby_33.t1 5.5105
R2774 standby_33.n0 standby_33 1.67737
R2775 ibias.n7 ibias.n1 1544.9
R2776 ibias.n4 ibias.n3 1544.9
R2777 ibias.n2 ibias.n0 300.425
R2778 ibias.n8 ibias.n2 300.425
R2779 ibias.n9 ibias.n0 177.746
R2780 ibias.n9 ibias.n8 177.746
R2781 ibias.n5 ibias.n1 139.143
R2782 ibias.n6 ibias.n3 139.143
R2783 ibias.n9 ibias.t1 60.1061
R2784 ibias.n4 ibias.n0 46.2505
R2785 ibias.n8 ibias.n7 46.2505
R2786 ibias.n5 ibias.n4 40.8622
R2787 ibias.n7 ibias.n6 40.8622
R2788 ibias.n3 ibias.n2 12.3338
R2789 ibias.n9 ibias.n1 12.3338
R2790 ibias.n6 ibias.t0 4.16651
R2791 ibias.t0 ibias.n5 4.16651
R2792 ibias ibias.n9 1.58676
R2793 ibias_ip ibias_ip.t13 31.8332
R2794 ibias_ip.t12 ibias_ip 31.4808
R2795 ibias_ip ibias_ip.t10 61.7027
R2796 ibias_ip.t0 ibias_ip 31.3394
R2797 ibias_ip ibias_ip.t1 39.498
R2798 ibias_ip.n0 ibias_ip.t11 31.8633
R2799 ibias_ip ibias_ip.t6 31.1832
R2800 ibias_ip.n1 ibias_ip.t2 31.1727
R2801 ibias_ip.n0 ibias_ip.t8 31.193
R2802 ibias_ip.n0 ibias_ip.t4 31.1967
R2803 ibias_ip.t3 ibias_ip.n1 39.8957
R2804 ibias_ip ibias_ip.t7 39.8329
R2805 ibias_ip.t5 ibias_ip.n0 39.8506
R2806 ibias_ip.n0 ibias_ip.t9 39.8715
R2807 ibias_ip ibias_ip.n1 1.87886
R2808 ibias_ip ibias_ip.n0 1.34188
R2809 avdd_ip.n81 avdd_ip.n73 58547.9
R2810 avdd_ip.n81 avdd_ip.n80 58547.9
R2811 avdd_ip.n79 avdd_ip.n73 58547.9
R2812 avdd_ip.n80 avdd_ip.n79 58547.9
R2813 avdd_ip.n43 avdd_ip.n42 54381
R2814 avdd_ip.n82 avdd_ip.n71 28978.4
R2815 avdd_ip.n82 avdd_ip.n72 28978.4
R2816 avdd_ip.n78 avdd_ip.n71 28978.4
R2817 avdd_ip.n78 avdd_ip.n72 28978.4
R2818 avdd_ip.n93 avdd_ip.n26 7296
R2819 avdd_ip.n91 avdd_ip.n26 7296
R2820 avdd_ip.n93 avdd_ip.n27 7296
R2821 avdd_ip.n91 avdd_ip.n27 7296
R2822 avdd_ip.n77 avdd_ip.n75 5062.04
R2823 avdd_ip.n75 avdd_ip.n74 3209.98
R2824 avdd_ip.n76 avdd_ip.n62 1005.14
R2825 avdd_ip.n44 avdd_ip.n36 857.648
R2826 avdd_ip.n40 avdd_ip.n37 857.648
R2827 avdd_ip.n44 avdd_ip.n37 857.648
R2828 avdd_ip.n55 avdd_ip.n54 857.648
R2829 avdd_ip.n57 avdd_ip.n50 857.648
R2830 avdd_ip.n43 avdd_ip.t3 337.433
R2831 avdd_ip.n77 avdd_ip.n76 269.44
R2832 avdd_ip.n57 avdd_ip.n56 267.182
R2833 avdd_ip.n54 avdd_ip.n51 267.182
R2834 avdd_ip.n41 avdd_ip.n40 267.182
R2835 avdd_ip.n84 avdd_ip.n63 212.139
R2836 avdd_ip.n90 avdd_ip.n89 202.696
R2837 avdd_ip.n88 avdd_ip.n29 134.065
R2838 avdd_ip.n74 avdd_ip.n29 110.358
R2839 avdd_ip.t7 avdd_ip.n26 105.665
R2840 avdd_ip.t11 avdd_ip.n27 105.665
R2841 avdd_ip.n85 avdd_ip.n84 96.3051
R2842 avdd_ip.n58 avdd_ip.n57 92.5005
R2843 avdd_ip.n55 avdd_ip.n49 92.5005
R2844 avdd_ip.n54 avdd_ip.n53 92.5005
R2845 avdd_ip.n52 avdd_ip.n50 92.5005
R2846 avdd_ip.n45 avdd_ip.n44 92.5005
R2847 avdd_ip.n44 avdd_ip.n43 92.5005
R2848 avdd_ip.n38 avdd_ip.n37 92.5005
R2849 avdd_ip.t3 avdd_ip.n37 92.5005
R2850 avdd_ip.n40 avdd_ip.n39 92.5005
R2851 avdd_ip.n36 avdd_ip.n35 92.5005
R2852 avdd_ip.n39 avdd_ip.n35 91.4862
R2853 avdd_ip.n53 avdd_ip.n49 91.4829
R2854 avdd_ip.n92 avdd_ip.t7 79.5673
R2855 avdd_ip.n92 avdd_ip.t11 79.5673
R2856 avdd_ip.n85 avdd_ip.n62 73.3959
R2857 avdd_ip.n39 avdd_ip.n38 66.8321
R2858 avdd_ip.n53 avdd_ip.n52 66.3131
R2859 avdd_ip.n59 avdd_ip.n49 63.936
R2860 avdd_ip.n46 avdd_ip.n35 63.936
R2861 avdd_ip.n2 avdd_ip.t6 62.0945
R2862 avdd_ip.n17 avdd_ip.t23 61.1041
R2863 avdd_ip.n15 avdd_ip.t24 60.1061
R2864 avdd_ip.n14 avdd_ip.t21 60.1061
R2865 avdd_ip.n21 avdd_ip.t26 60.1061
R2866 avdd_ip.n24 avdd_ip.t20 60.1061
R2867 avdd_ip.n89 avdd_ip.t15 60.1061
R2868 avdd_ip.n89 avdd_ip.t12 60.1061
R2869 avdd_ip.n89 avdd_ip.t13 60.1061
R2870 avdd_ip.n63 avdd_ip.t10 60.1061
R2871 avdd_ip.n63 avdd_ip.t8 60.1061
R2872 avdd_ip.n63 avdd_ip.t9 60.1061
R2873 avdd_ip.n31 avdd_ip.t16 60.1061
R2874 avdd_ip.n31 avdd_ip.t14 60.1061
R2875 avdd_ip.n30 avdd_ip.t18 60.1061
R2876 avdd_ip.n30 avdd_ip.t17 60.1061
R2877 avdd_ip.n65 avdd_ip.t27 60.1061
R2878 avdd_ip.n65 avdd_ip.t19 60.1061
R2879 avdd_ip.n64 avdd_ip.t28 60.1061
R2880 avdd_ip.n64 avdd_ip.t22 60.1061
R2881 avdd_ip.n16 avdd_ip.t25 60.1061
R2882 avdd_ip.n41 avdd_ip.n36 57.4849
R2883 avdd_ip.n56 avdd_ip.n55 57.4849
R2884 avdd_ip.n51 avdd_ip.n50 57.4849
R2885 avdd_ip.n2 avdd_ip.n1 55.1707
R2886 avdd_ip.n2 avdd_ip.n0 54.9038
R2887 avdd_ip.n69 avdd_ip.n13 44.6614
R2888 avdd_ip.n58 avdd_ip.n48 43.3376
R2889 avdd_ip.n45 avdd_ip.n34 43.3376
R2890 avdd_ip.n83 avdd_ip.n70 30.1747
R2891 avdd_ip.n51 avdd_ip.t5 28.8172
R2892 avdd_ip.n56 avdd_ip.t5 28.8172
R2893 avdd_ip.t3 avdd_ip.n41 28.8172
R2894 avdd_ip.n90 avdd_ip.n28 10.6324
R2895 avdd_ip.n74 avdd_ip.n25 8.37369
R2896 avdd_ip.n16 avdd_ip.n15 7.25561
R2897 avdd_ip.n0 avdd_ip.t1 6.92425
R2898 avdd_ip.n0 avdd_ip.t4 6.92425
R2899 avdd_ip.n1 avdd_ip.t0 6.92425
R2900 avdd_ip.n1 avdd_ip.t2 6.92425
R2901 avdd_ip.n91 avdd_ip.n90 6.37981
R2902 avdd_ip.n92 avdd_ip.n91 6.37981
R2903 avdd_ip.n94 avdd_ip.n93 6.37981
R2904 avdd_ip.n93 avdd_ip.n92 6.37981
R2905 avdd_ip.n24 avdd_ip.n23 6.17839
R2906 avdd_ip.n78 avdd_ip.n77 6.15262
R2907 avdd_ip.n94 avdd_ip.n25 5.31953
R2908 avdd_ip.n52 avdd_ip.n48 4.38907
R2909 avdd_ip.n38 avdd_ip.n34 4.38907
R2910 avdd_ip.n95 avdd_ip.n94 3.87825
R2911 avdd_ip.n84 avdd_ip.n83 3.6009
R2912 avdd_ip.n60 avdd_ip.n48 2.4925
R2913 avdd_ip.n47 avdd_ip.n34 2.44611
R2914 avdd_ip.n29 avdd_ip.n27 2.43471
R2915 avdd_ip.n70 avdd_ip.n26 2.43471
R2916 avdd_ip.n59 avdd_ip.n58 2.37764
R2917 avdd_ip.n46 avdd_ip.n45 2.37764
R2918 avdd_ip.n60 avdd_ip.n59 2.3255
R2919 avdd_ip.n47 avdd_ip.n46 2.3255
R2920 avdd_ip.n22 avdd_ip.n21 1.87566
R2921 avdd_ip.n95 avdd_ip.n13 1.41891
R2922 avdd_ip.n4 avdd_ip.n3 1.18871
R2923 avdd_ip.n23 avdd_ip.n14 1.07773
R2924 avdd_ip.n79 avdd_ip.n78 1.05764
R2925 avdd_ip.n83 avdd_ip.n82 1.05764
R2926 avdd_ip.n82 avdd_ip.n81 1.05764
R2927 avdd_ip.n86 avdd_ip.n85 1.02375
R2928 avdd_ip.n21 avdd_ip.n20 0.982678
R2929 avdd_ip.n20 avdd_ip.n14 0.919312
R2930 avdd_ip.n17 avdd_ip.n16 0.90347
R2931 avdd_ip.n23 avdd_ip.n22 0.845955
R2932 avdd_ip.n11 avdd_ip.n4 0.827286
R2933 avdd_ip avdd_ip.n11 0.808179
R2934 avdd_ip.n66 avdd_ip.n64 0.65712
R2935 avdd_ip.n32 avdd_ip.n30 0.652725
R2936 avdd_ip.n88 avdd_ip.n87 0.613954
R2937 avdd_ip.n76 avdd_ip.n72 0.530586
R2938 avdd_ip.n80 avdd_ip.n72 0.530586
R2939 avdd_ip.n75 avdd_ip.n71 0.530586
R2940 avdd_ip.n73 avdd_ip.n71 0.530586
R2941 avdd_ip.n3 avdd_ip.n2 0.507794
R2942 avdd_ip.n70 avdd_ip.n69 0.448948
R2943 avdd_ip.n19 avdd_ip.n18 0.402976
R2944 avdd_ip.n33 avdd_ip.n32 0.319749
R2945 avdd_ip.n87 avdd_ip.n86 0.319015
R2946 avdd_ip.n67 avdd_ip.n66 0.319015
R2947 avdd_ip.n18 avdd_ip.n12 0.319015
R2948 avdd_ip.n20 avdd_ip.n19 0.282318
R2949 avdd_ip.n11 avdd_ip.n10 0.255087
R2950 avdd_ip.n32 avdd_ip.n31 0.25137
R2951 avdd_ip.n66 avdd_ip.n65 0.25137
R2952 avdd_ip.n96 avdd_ip.n12 0.243945
R2953 avdd_ip avdd_ip.n97 0.213307
R2954 avdd_ip.n87 avdd_ip.n28 0.211864
R2955 avdd_ip.n18 avdd_ip.n17 0.211864
R2956 avdd_ip.n97 avdd_ip 0.18211
R2957 avdd_ip.n25 avdd_ip.n24 0.174542
R2958 avdd_ip.n15 avdd_ip.n13 0.174542
R2959 avdd_ip.n62 avdd_ip.n61 0.166571
R2960 avdd_ip.n67 avdd_ip.n12 0.150396
R2961 avdd_ip.n86 avdd_ip.n33 0.150396
R2962 avdd_ip.n3 avdd_ip.t33 0.125045
R2963 avdd_ip.n7 avdd_ip.n4 0.123905
R2964 avdd_ip.n68 avdd_ip.n33 0.117461
R2965 avdd_ip.n10 avdd_ip.n9 0.111971
R2966 avdd_ip.n8 avdd_ip.n7 0.110265
R2967 avdd_ip.n68 avdd_ip.n67 0.108384
R2968 avdd_ip.n6 avdd_ip.n5 0.106696
R2969 avdd_ip.n9 avdd_ip.n8 0.106696
R2970 avdd_ip.n61 avdd_ip.n47 0.0839309
R2971 avdd_ip.n61 avdd_ip.n60 0.0812962
R2972 avdd_ip.n5 avdd_ip.t30 0.0180781
R2973 avdd_ip.n9 avdd_ip.t32 0.0180781
R2974 avdd_ip.n8 avdd_ip.t29 0.0180781
R2975 avdd_ip.n6 avdd_ip.t31 0.0180781
R2976 avdd_ip.n10 avdd_ip.n5 0.0174228
R2977 avdd_ip.n96 avdd_ip.n95 0.0173478
R2978 avdd_ip.n63 avdd_ip.n28 0.0154184
R2979 avdd_ip.n89 avdd_ip.n88 0.0154184
R2980 avdd_ip.n7 avdd_ip.n6 0.0150053
R2981 avdd_ip.n69 avdd_ip.n68 0.0108333
R2982 avdd_ip.n97 avdd_ip.n96 0.00292843
R2983 avdd_ip.n22 avdd_ip.n19 0.000885802
R2984 xout.n29 xout.t26 594.784
R2985 xout.n29 xout.t24 194.649
R2986 xout.n25 xout.t23 124.457
R2987 xout.n25 xout.t25 106.793
R2988 xout.t23 xout.n24 86.3125
R2989 xout.t25 xout.n23 86.3125
R2990 xout.n3 xout.t18 62.0071
R2991 xout.n4 xout.t16 62.0071
R2992 xout.n3 xout.t11 60.1061
R2993 xout.n4 xout.t12 60.1061
R2994 xout.n8 xout.t14 60.1061
R2995 xout.n8 xout.t13 60.1061
R2996 xout.n10 xout.t17 60.1061
R2997 xout.n10 xout.t15 60.1061
R2998 xout.n0 xout.t20 60.1061
R2999 xout.n0 xout.t22 60.1061
R3000 xout.n1 xout.t19 60.1061
R3001 xout.n1 xout.t21 60.1061
R3002 xout.n24 xout.n23 58.6245
R3003 xout.n22 xout.t3 43.5339
R3004 xout.n28 xout.n27 21.3269
R3005 xout.n16 xout.n15 18.5533
R3006 xout.n20 xout.n13 18.553
R3007 xout.n19 xout.n18 18.4723
R3008 xout.n19 xout.n17 18.4564
R3009 xout.n16 xout.n14 18.4564
R3010 xout.n27 xout.n23 12.2455
R3011 xout.n18 xout.t9 4.133
R3012 xout.n18 xout.t5 4.133
R3013 xout.n17 xout.t6 4.133
R3014 xout.n17 xout.t10 4.133
R3015 xout.n15 xout.t8 4.133
R3016 xout.n15 xout.t2 4.133
R3017 xout.n14 xout.t0 4.133
R3018 xout.n14 xout.t4 4.133
R3019 xout.n13 xout.t1 4.133
R3020 xout.n13 xout.t7 4.133
R3021 xout.n5 xout.n4 3.64406
R3022 xout.n5 xout.n3 3.61238
R3023 xout.n26 xout.n24 3.56553
R3024 xout.n22 xout.n21 2.24362
R3025 xout.n29 xout.n28 2.18092
R3026 xout.n28 xout.n22 1.03102
R3027 xout.n27 xout.n26 0.742745
R3028 xout.n26 xout.n25 0.715885
R3029 xout.n21 xout.n12 0.464586
R3030 xout.n2 xout.n0 0.424187
R3031 xout.n11 xout.n9 0.402558
R3032 xout xout.n29 0.377063
R3033 xout.n6 xout.n2 0.316998
R3034 xout.n2 xout.n1 0.310571
R3035 xout.n12 xout.n7 0.273717
R3036 xout.n7 xout.n6 0.261913
R3037 xout.n9 xout.n8 0.254998
R3038 xout.n11 xout.n10 0.25137
R3039 xout.n6 xout.n5 0.143668
R3040 xout.n9 xout.n7 0.126918
R3041 xout.n12 xout.n11 0.125886
R3042 xout.n21 xout.n20 0.0947164
R3043 xout.n20 xout.n16 0.0657574
R3044 xout.n20 xout.n19 0.0480746
R3045 inv_in.n19 inv_in.t0 47.4896
R3046 inv_in.n18 inv_in.t3 6.48745
R3047 inv_in.n19 inv_in.t1 6.24255
R3048 inv_in inv_in.n17 2.2182
R3049 inv_in.n18 inv_in 0.342687
R3050 inv_in inv_in.n18 0.217687
R3051 inv_in.n5 inv_in.n4 0.110198
R3052 inv_in.n7 inv_in.n6 0.110101
R3053 inv_in.n10 inv_in.n9 0.110101
R3054 inv_in.n8 inv_in.n2 0.110101
R3055 inv_in.n16 inv_in.n15 0.109734
R3056 inv_in.n14 inv_in.n0 0.109734
R3057 inv_in.n13 inv_in.n12 0.109709
R3058 inv_in.n11 inv_in.n1 0.109709
R3059 inv_in.n9 inv_in.n7 0.109325
R3060 inv_in.n9 inv_in.n8 0.109325
R3061 inv_in.n12 inv_in.n11 0.109325
R3062 inv_in.n11 inv_in.n3 0.109325
R3063 inv_in.n15 inv_in.n14 0.1086
R3064 inv_in.n16 inv_in.n0 0.1086
R3065 inv_in.n4 inv_in.n3 0.10222
R3066 inv_in.n7 inv_in.n5 0.101755
R3067 inv_in inv_in.n19 0.09425
R3068 inv_in.n18 inv_in 0.063
R3069 inv_in.n0 inv_in.t11 0.00880157
R3070 inv_in.n7 inv_in.t9 0.00848368
R3071 inv_in.n9 inv_in.t10 0.00848368
R3072 inv_in.n8 inv_in.t2 0.00848368
R3073 inv_in.n5 inv_in.t12 0.00838586
R3074 inv_in.n4 inv_in.t14 0.0083125
R3075 inv_in.n6 inv_in.t13 0.0083125
R3076 inv_in.n2 inv_in.t6 0.0083125
R3077 inv_in.n10 inv_in.t4 0.0083125
R3078 inv_in.n1 inv_in.t5 0.0083125
R3079 inv_in.n13 inv_in.t8 0.0083125
R3080 inv_in.n17 inv_in.t7 0.0083125
R3081 inv_in.n6 inv_in.n3 0.00106244
R3082 inv_in.n12 inv_in.n2 0.00106244
R3083 inv_in.n11 inv_in.n10 0.00106244
R3084 inv_in.n17 inv_in.n16 0.000989074
R3085 inv_in.n15 inv_in.n1 0.000548907
R3086 inv_in.n14 inv_in.n13 0.000548907
R3087 inv_m1.t0 inv_m1.n0 229.685
R3088 inv_m1.n0 inv_m1.t1 652.083
R3089 inv_m1 inv_m1.n0 4.5555
R3090 inv_m1 inv_m1.n3 1.058
R3091 inv_m1.n3 inv_m1.n2 24.8426
R3092 inv_m1.n2 inv_m1.t4 20.438
R3093 inv_m1.n2 inv_m1.t3 20.4375
R3094 inv_m1.n3 inv_m1.n1 24.7082
R3095 inv_m1.n1 inv_m1.t5 21.9207
R3096 inv_m1.n1 inv_m1.t2 21.9202
R3097 a_2132_n15590.t0 a_2132_n15590.t1 82.3309
R3098 a_18932_n15756.t0 a_18932_n15756.t1 83.5579
R3099 inv_m2 inv_m2.t1 651.861
R3100 inv_m2 inv_m2.t0 229.522
R3101 inv_m2 inv_m2.t2 108.124
R3102 inv_m2.t5 inv_m2 108.124
R3103 inv_m2.n0 inv_m2 80.6505
R3104 inv_m2.t2 inv_m2.n0 27.4745
R3105 inv_m2.n0 inv_m2.t5 27.4745
R3106 inv_m2 inv_m2.n1 24.0208
R3107 inv_m2.n1 inv_m2.t3 20.4885
R3108 inv_m2.n1 inv_m2.t4 20.387
R3109 dout_ip.n0 dout_ip.t2 651.692
R3110 dout_ip.n0 dout_ip.t3 651.431
R3111 dout_ip.n1 dout_ip.t9 288.204
R3112 dout_ip.n5 dout_ip.t5 264.103
R3113 dout_ip.n2 dout_ip.t6 264.103
R3114 dout_ip.n0 dout_ip.t1 229.352
R3115 dout_ip.n0 dout_ip.t0 229.101
R3116 dout_ip.n1 dout_ip.t7 195.017
R3117 x7.x2.clkin dout_ip.n5 159.236
R3118 x7.x1.clkin dout_ip.n2 159.236
R3119 x7.x5.A dout_ip.n1 153.153
R3120 dout_ip.n4 x7.x2.x1.A 152
R3121 x7.x1.x1.A dout_ip.n3 152
R3122 dout_ip.n4 dout_ip.t8 145.209
R3123 dout_ip.n3 dout_ip.t4 145.209
R3124 dout_ip.n7 dout_ip.n6 117.519
R3125 dout_ip.n6 x7.x1.clkin 68.1959
R3126 dout_ip.n5 dout_ip.n4 37.6741
R3127 dout_ip.n3 dout_ip.n2 37.6741
R3128 x7.clkin dout_ip.n7 31.6505
R3129 dout_ip.n7 x7.x5.A 24.4485
R3130 x7.clkin dout_ip.n0 11.4719
R3131 x7.x2.clkin x7.x2.x1.A 10.3444
R3132 x7.x1.clkin x7.x1.x1.A 10.3444
R3133 dout_ip.n6 x7.x2.clkin 9.3005
R3134 a_20689_n2549.n3 a_20689_n2549.n2 647.119
R3135 a_20689_n2549.n1 a_20689_n2549.t4 350.253
R3136 a_20689_n2549.n2 a_20689_n2549.n0 260.339
R3137 a_20689_n2549.n2 a_20689_n2549.n1 246.119
R3138 a_20689_n2549.n1 a_20689_n2549.t5 189.588
R3139 a_20689_n2549.n3 a_20689_n2549.t3 89.1195
R3140 a_20689_n2549.n0 a_20689_n2549.t2 63.3338
R3141 a_20689_n2549.t0 a_20689_n2549.n3 41.0422
R3142 a_20689_n2549.n0 a_20689_n2549.t1 31.9797
R3143 a_20567_n2791.t0 a_20567_n2791.t1 198.571
R3144 a_20733_n2791.t0 a_20733_n2791.t1 60.0005
R3145 xin_buf.n0 xin_buf.t1 9.98044
R3146 xin_buf.n1 xin_buf.t4 6.0819
R3147 xin_buf.n0 xin_buf.t0 3.49292
R3148 xin_buf.n1 xin_buf.t2 2.23853
R3149 xin_buf.n1 xin_buf.t3 10.3359
R3150 xin_buf.n0 xin_buf.t3 28.8094
R3151 a_15000_n1881.n2 a_15000_n1881.n1 682.193
R3152 a_15000_n1881.n0 a_15000_n1881.t4 279.142
R3153 a_15000_n1881.n1 a_15000_n1881.t2 250.737
R3154 a_15000_n1881.n0 a_15000_n1881.t3 145.958
R3155 a_15000_n1881.n1 a_15000_n1881.n0 118.45
R3156 a_15000_n1881.n2 a_15000_n1881.t1 70.3576
R3157 a_15000_n1881.t0 a_15000_n1881.n2 65.6672
R3158 x7.x1.x2.CLK x7.x1.x2.CLK.t0 716.451
R3159 x7.x1.x2.CLK.t0 x7.x1.x2.CLK.n3 707.66
R3160 x7.x1.x2.CLK.n0 x7.x1.x2.CLK.t2 294.557
R3161 x7.x1.x2.CLK.n2 x7.x1.x2.CLK.t1 271.777
R3162 x7.x1.x2.CLK.n0 x7.x1.x2.CLK.t3 211.01
R3163 x7.x1.x2.CLK.n1 x7.x1.x2.CLK.n0 152
R3164 x7.x1.x2.CLK.n3 x7.x1.x2.CLK.n2 38.2982
R3165 x7.x1.x2.CLK.n2 x7.x1.x2.CLK.n1 33.0611
R3166 x7.x1.x2.CLK x7.x1.x2.CLK.n3 8.88521
R3167 x7.x1.x2.CLK.n1 x7.x1.x2.CLK 4.20621
R3168 a_16151_n1869.t0 a_16151_n1869.t1 198.571
R3169 a_16317_n1881.t0 a_16317_n1881.t1 60.0005
R3170 a_21775_n2791.t0 a_21775_n2791.n1 386.31
R3171 a_21775_n2791.n1 a_21775_n2791.t1 249.956
R3172 a_21775_n2791.n0 a_21775_n2791.t3 239.04
R3173 a_21775_n2791.n1 a_21775_n2791.n0 175.661
R3174 a_21775_n2791.n0 a_21775_n2791.t2 166.739
R3175 x7.clk_disable.n3 x7.clk_disable.t0 319.219
R3176 x7.clk_disable.n1 x7.clk_disable.t4 268.313
R3177 x7.clk_disable x7.clk_disable.t1 249.867
R3178 x7.clk_disable.n2 x7.clk_disable.t2 206.19
R3179 x7.clk_disable.n1 x7.clk_disable.t5 186.374
R3180 x7.clk_disable x7.clk_disable.n2 152
R3181 x7.clk_disable.n2 x7.clk_disable.n1 148.35
R3182 x7.clk_disable x7.clk_disable.n0 32.2121
R3183 x7.clk_disable x7.clk_disable.t3 21.881
R3184 x7.clk_disable.n3 x7.clk_disable 21.8175
R3185 x7.clk_disable.n0 x7.clk_disable 11.0708
R3186 x7.clk_disable.n0 x7.clk_disable 8.03187
R3187 x7.clk_disable x7.clk_disable.n3 4.14393
R3188 a_14009_n2701.t0 a_14009_n2701.n0 753.673
R3189 a_14009_n2701.n0 a_14009_n2701.t2 354.81
R3190 a_14009_n2701.n0 a_14009_n2701.t1 303.562
R3191 standby_ip.t1 standby_ip.n3 368.26
R3192 standby_ip.n2 standby_ip.n3 1.85916
R3193 standby_ip.n17 standby_ip.t4 405.389
R3194 standby_ip.t4 standby_ip.n16 405.389
R3195 standby_ip.t15 standby_ip.n8 405.389
R3196 standby_ip.n9 standby_ip.t15 405.389
R3197 standby_ip.n17 standby_ip.t6 375.649
R3198 standby_ip.t6 standby_ip.n16 375.649
R3199 standby_ip.t17 standby_ip.n18 375.649
R3200 standby_ip.n19 standby_ip.t17 375.649
R3201 standby_ip.t18 standby_ip.n15 375.649
R3202 standby_ip.n20 standby_ip.t18 375.649
R3203 standby_ip.n22 standby_ip.t5 375.649
R3204 standby_ip.t5 standby_ip.n21 375.649
R3205 standby_ip.n14 standby_ip.t11 375.649
R3206 standby_ip.t11 standby_ip.n13 375.649
R3207 standby_ip.t12 standby_ip.n7 375.649
R3208 standby_ip.n12 standby_ip.t12 375.649
R3209 standby_ip.t8 standby_ip.n10 375.649
R3210 standby_ip.n11 standby_ip.t8 375.649
R3211 standby_ip.n9 standby_ip.t9 375.649
R3212 standby_ip.t9 standby_ip.n8 375.649
R3213 standby_ip.t13 standby_ip.n23 332.752
R3214 standby_ip.n24 standby_ip.t13 332.75
R3215 standby_ip.t7 standby_ip.n23 332.411
R3216 standby_ip.n24 standby_ip.t7 332.411
R3217 standby_ip.n4 standby_ip.t3 231.718
R3218 standby_ip standby_ip.t0 216.155
R3219 standby_ip standby_ip.n5 161.314
R3220 standby_ip.n4 standby_ip.t14 159.417
R3221 standby_ip.n5 standby_ip.n4 152
R3222 standby_ip standby_ip.t16 59.9857
R3223 standby_ip standby_ip.t2 59.3654
R3224 standby_ip standby_ip.n2 46.2227
R3225 standby_ip.n11 standby_ip.n8 29.7417
R3226 standby_ip.n12 standby_ip.n11 29.7417
R3227 standby_ip.n13 standby_ip.n12 29.7417
R3228 standby_ip.n21 standby_ip.n20 29.7417
R3229 standby_ip.n20 standby_ip.n19 29.7417
R3230 standby_ip.n19 standby_ip.n16 29.7417
R3231 standby_ip.n10 standby_ip.n9 29.7417
R3232 standby_ip.n10 standby_ip.n7 29.7417
R3233 standby_ip.n14 standby_ip.n7 29.7417
R3234 standby_ip.n22 standby_ip.n15 29.7417
R3235 standby_ip.n18 standby_ip.n15 29.7417
R3236 standby_ip.n18 standby_ip.n17 29.7417
R3237 standby_ip.n13 standby_ip.n6 16.7534
R3238 standby_ip.n0 standby_ip.n14 16.7534
R3239 standby_ip.n1 standby_ip 13.0593
R3240 standby_ip.n21 standby_ip.n6 12.9887
R3241 standby_ip.n0 standby_ip.n22 12.9887
R3242 standby_ip standby_ip.t10 12.6603
R3243 standby_ip standby_ip.n26 9.27339
R3244 standby_ip.n25 standby_ip.n23 5.53161
R3245 standby_ip.n26 standby_ip.n2 5.46183
R3246 standby_ip standby_ip.n1 5.4255
R3247 standby_ip.n25 standby_ip.n24 4.67076
R3248 standby_ip.n3 standby_ip 1.88798
R3249 standby_ip standby_ip.n25 3.51723
R3250 standby_ip.n2 standby_ip 2.98717
R3251 standby_ip.n1 standby_ip.n6 2.80971
R3252 standby_ip.n26 standby_ip 2.78266
R3253 standby_ip.n5 standby_ip 2.74336
R3254 standby_ip.n1 standby_ip.n0 2.49791
R3255 a_2971_n1521.t0 a_2971_n1521.n1 405.735
R3256 a_2971_n1521.n1 a_2971_n1521.t1 294.611
R3257 a_2971_n1521.n0 a_2971_n1521.t3 254.389
R3258 a_2971_n1521.n0 a_2971_n1521.t2 211.01
R3259 a_2971_n1521.n1 a_2971_n1521.n0 152
R3260 a_14035_n1997.t0 a_14035_n1997.t1 38.7697
R3261 a_2132_n17582.t0 a_2132_n17582.t1 83.9053
R3262 a_18932_n17416.t0 a_18932_n17416.t1 83.5579
R3263 avss.n20 avss.n19 18580.7
R3264 avss.n38 avss.n37 15308.7
R3265 avss.n76 avss.n20 12246.6
R3266 avss.n40 avss.n35 3599.36
R3267 avss.n41 avss.n35 3599.36
R3268 avss.n41 avss.n34 3599.36
R3269 avss.n40 avss.n34 3599.36
R3270 avss.n67 avss.n25 2489.59
R3271 avss.n67 avss.n26 2489.59
R3272 avss.n69 avss.n26 2489.59
R3273 avss.n69 avss.n25 2489.59
R3274 avss.n28 avss.n21 2489.59
R3275 avss.n28 avss.n22 2489.59
R3276 avss.n74 avss.n22 2489.59
R3277 avss.n74 avss.n21 2489.59
R3278 avss.n78 avss.n13 2489.59
R3279 avss.n78 avss.n14 2489.59
R3280 avss.n16 avss.n14 2489.59
R3281 avss.n16 avss.n13 2489.59
R3282 avss.n88 avss.n6 2489.59
R3283 avss.n90 avss.n6 2489.59
R3284 avss.n90 avss.n5 2489.59
R3285 avss.n88 avss.n5 2489.59
R3286 avss.n36 avss.n20 2342.14
R3287 avss.n77 avss.n76 930.542
R3288 avss.n76 avss.n75 930.542
R3289 avss.n43 avss.n42 881.42
R3290 avss.n19 avss.t6 633.244
R3291 avss.n15 avss.t4 633.244
R3292 avss.t20 avss.n17 633.244
R3293 avss.n77 avss.t22 633.244
R3294 avss.n75 avss.t10 633.244
R3295 avss.n29 avss.t12 633.244
R3296 avss.t0 avss.n30 633.244
R3297 avss.n37 avss.t2 633.244
R3298 avss.t24 avss.n36 412.863
R3299 avss.t14 avss.n38 397.358
R3300 avss.n17 avss.n15 362.704
R3301 avss.n30 avss.n29 362.704
R3302 avss.t18 avss.t24 306.255
R3303 avss.t8 avss.t18 306.255
R3304 avss.t8 avss.t16 306.255
R3305 avss.t16 avss.t14 306.255
R3306 avss.n39 avss.n32 295.807
R3307 avss.n66 avss.n65 289.13
R3308 avss.n87 avss.n3 289.13
R3309 avss.n92 avss.n91 288.753
R3310 avss.n70 avss.n24 288.753
R3311 avss.n89 avss.t6 234.865
R3312 avss.n89 avss.t4 234.865
R3313 avss.n18 avss.t20 234.865
R3314 avss.t22 avss.n18 234.865
R3315 avss.n27 avss.t10 234.865
R3316 avss.t12 avss.n27 234.865
R3317 avss.n68 avss.t0 234.865
R3318 avss.n68 avss.t2 234.865
R3319 avss.n31 avss.n10 152.73
R3320 avss.n73 avss.n72 152.73
R3321 avss.n80 avss.n7 152.73
R3322 avss.n79 avss.n12 152.73
R3323 avss.n39 avss.n33 118.081
R3324 avss.n91 avss.n4 103.529
R3325 avss.n64 avss.n31 103.529
R3326 avss.n72 avss.n71 103.529
R3327 avss.n66 avss.n64 103.529
R3328 avss.n71 avss.n70 103.529
R3329 avss.n86 avss.n7 103.529
R3330 avss.n12 avss.n4 103.529
R3331 avss.n87 avss.n86 103.529
R3332 avss.n88 avss.n87 97.5005
R3333 avss.n89 avss.n88 97.5005
R3334 avss.n91 avss.n90 97.5005
R3335 avss.n90 avss.n89 97.5005
R3336 avss.n13 avss.n7 97.5005
R3337 avss.n18 avss.n13 97.5005
R3338 avss.n14 avss.n12 97.5005
R3339 avss.n18 avss.n14 97.5005
R3340 avss.n31 avss.n21 97.5005
R3341 avss.n27 avss.n21 97.5005
R3342 avss.n72 avss.n22 97.5005
R3343 avss.n27 avss.n22 97.5005
R3344 avss.n70 avss.n69 97.5005
R3345 avss.n69 avss.n68 97.5005
R3346 avss.n67 avss.n66 97.5005
R3347 avss.n68 avss.n67 97.5005
R3348 avss.n42 avss.n33 69.8003
R3349 avss.n38 avss.n35 54.5071
R3350 avss.n5 avss.n3 48.7505
R3351 avss.n19 avss.n5 48.7505
R3352 avss.n8 avss.n6 48.7505
R3353 avss.n15 avss.n6 48.7505
R3354 avss.n16 avss.n8 48.7505
R3355 avss.n17 avss.n16 48.7505
R3356 avss.n79 avss.n78 48.7505
R3357 avss.n78 avss.n77 48.7505
R3358 avss.n74 avss.n73 48.7505
R3359 avss.n75 avss.n74 48.7505
R3360 avss.n28 avss.n23 48.7505
R3361 avss.n29 avss.n28 48.7505
R3362 avss.n25 avss.n23 48.7505
R3363 avss.n30 avss.n25 48.7505
R3364 avss.n65 avss.n26 48.7505
R3365 avss.n37 avss.n26 48.7505
R3366 avss.n40 avss.n39 45.0005
R3367 avss.t8 avss.n40 45.0005
R3368 avss.n42 avss.n41 45.0005
R3369 avss.n41 avss.t8 45.0005
R3370 avss.n64 avss.n63 40.3697
R3371 avss.n71 avss.n23 40.3697
R3372 avss.n86 avss.n85 40.3697
R3373 avss.n8 avss.n4 40.3697
R3374 avss.n94 avss.n1 39.7977
R3375 avss.n34 avss.n33 39.0005
R3376 avss.n36 avss.n34 39.0005
R3377 avss.n35 avss.n32 39.0005
R3378 avss.n94 avss 33.7505
R3379 avss.n84 avss.t21 29.9199
R3380 avss.n62 avss.t1 29.9199
R3381 avss.n62 avss.t13 29.9199
R3382 avss.n84 avss.t5 29.9199
R3383 avss.n2 avss.t7 29.798
R3384 avss.n57 avss.t3 29.798
R3385 avss.n11 avss.t23 29.798
R3386 avss.n11 avss.t11 29.798
R3387 avss.n32 avss.t15 20.9512
R3388 avss.n46 avss.n45 18.8362
R3389 avss.n46 avss.n44 18.6458
R3390 avss.n44 avss.t9 4.133
R3391 avss.n44 avss.t17 4.133
R3392 avss.n45 avss.t25 4.133
R3393 avss.n45 avss.t19 4.133
R3394 avss.n47 avss.n43 1.61679
R3395 avss.n55 avss 1.33946
R3396 avss.n58 avss.n24 1.21803
R3397 avss.n93 avss.n92 1.21803
R3398 avss.n54 avss.n47 0.8655
R3399 avss.n63 avss.n62 0.664786
R3400 avss.n81 avss.n10 0.664786
R3401 avss.n81 avss.n80 0.664786
R3402 avss.n85 avss.n84 0.664786
R3403 avss.n55 avss.n54 0.53175
R3404 avss.n56 avss.n9 0.434977
R3405 avss.n95 avss.n0 0.433066
R3406 avss.n61 avss.n59 0.433066
R3407 avss.n61 avss.n60 0.433066
R3408 avss.n60 avss.n0 0.433066
R3409 avss.n65 avss.n24 0.376971
R3410 avss.n92 avss.n3 0.376971
R3411 avss.n84 avss.n0 0.299413
R3412 avss.n62 avss.n61 0.299413
R3413 avss.n62 avss.n9 0.247783
R3414 avss.n84 avss.n83 0.247783
R3415 avss.n83 avss 0.245943
R3416 avss.n59 avss.n58 0.231236
R3417 avss.n82 avss.n9 0.201672
R3418 avss.n83 avss.n82 0.201672
R3419 avss.n2 avss.n1 0.2005
R3420 avss.n95 avss.n94 0.2005
R3421 avss.n47 avss.n46 0.1855
R3422 avss.n49 avss.n48 0.122162
R3423 avss.n82 avss.n81 0.120904
R3424 avss.n50 avss.n49 0.105544
R3425 avss.n51 avss.n50 0.101695
R3426 avss.n73 avss.n10 0.1005
R3427 avss.n80 avss.n79 0.1005
R3428 avss.n60 avss.n11 0.0997647
R3429 avss.n53 avss.n48 0.0989292
R3430 avss.n56 avss.n55 0.096886
R3431 avss.n54 avss.n53 0.0847138
R3432 avss.n63 avss.n23 0.0825513
R3433 avss.n85 avss.n8 0.0825513
R3434 avss.n51 avss.n48 0.0586846
R3435 avss.n57 avss.n56 0.0480171
R3436 avss avss.n95 0.0332586
R3437 avss.n59 avss 0.0330342
R3438 avss.n94 avss.n93 0.0328276
R3439 avss.n43 avss.n32 0.0328232
R3440 avss.n53 avss.n52 0.0277801
R3441 avss.n50 avss.t28 0.0083125
R3442 avss.n49 avss.t29 0.0083125
R3443 avss.n48 avss.t26 0.0083125
R3444 avss.n52 avss.t27 0.0083125
R3445 avss avss.n1 0.00342969
R3446 avss.n93 avss.n2 0.000931034
R3447 avss.n58 avss.n57 0.000928082
R3448 avss.n81 avss.n11 0.000683824
R3449 avss.n52 avss.n51 0.000622332
R3450 avdd.n92 avdd.n91 15807.9
R3451 avdd.n93 avdd.n92 15807.9
R3452 avdd.n93 avdd.n28 15807.9
R3453 avdd.n91 avdd.n28 15807.9
R3454 avdd.n90 avdd.n27 8112.97
R3455 avdd.n94 avdd.n27 8112.97
R3456 avdd.n94 avdd.n26 8112.97
R3457 avdd.n90 avdd.n26 8112.97
R3458 avdd.n98 avdd.n6 2166
R3459 avdd.n97 avdd.n6 2166
R3460 avdd.n98 avdd.n7 2166
R3461 avdd.n97 avdd.n7 2166
R3462 avdd.n78 avdd.n77 1643.17
R3463 avdd.n77 avdd.n76 1643.17
R3464 avdd.n74 avdd.n69 1643.17
R3465 avdd.n80 avdd.n69 1643.17
R3466 avdd.n52 avdd.n37 1643.17
R3467 avdd.n60 avdd.n37 1643.17
R3468 avdd.n55 avdd.n54 1643.17
R3469 avdd.n58 avdd.n55 1643.17
R3470 avdd.n89 avdd.n88 1439.4
R3471 avdd.n89 avdd.n29 1352.37
R3472 avdd.n66 avdd.n25 1313.54
R3473 avdd.n71 avdd.n70 1106.59
R3474 avdd.n70 avdd.n68 1106.59
R3475 avdd.n40 avdd.n39 1106.59
R3476 avdd.n39 avdd.n36 1106.59
R3477 avdd.n78 avdd.n68 536.587
R3478 avdd.n76 avdd.n71 536.587
R3479 avdd.n74 avdd.n71 536.587
R3480 avdd.n80 avdd.n68 536.587
R3481 avdd.n52 avdd.n40 536.587
R3482 avdd.n54 avdd.n40 536.587
R3483 avdd.n58 avdd.n36 536.587
R3484 avdd.n60 avdd.n36 536.587
R3485 avdd.n75 avdd.t2 382.582
R3486 avdd.n79 avdd.t2 382.582
R3487 avdd.n53 avdd.t0 382.582
R3488 avdd.n59 avdd.t0 382.582
R3489 avdd.n73 avdd.n30 319.248
R3490 avdd.n57 avdd.n56 319.248
R3491 avdd.n88 avdd.n31 287.265
R3492 avdd.n38 avdd.n29 287.265
R3493 avdd.n88 avdd.n30 276.295
R3494 avdd.n56 avdd.n29 276.295
R3495 avdd.n86 avdd.t3 227.377
R3496 avdd.n1 avdd.t6 227.377
R3497 avdd.n34 avdd.t1 227.377
R3498 avdd.n43 avdd.t17 227.377
R3499 avdd.n66 avdd.n3 205.554
R3500 avdd.n72 avdd.n31 189.742
R3501 avdd.n38 avdd.n35 189.742
R3502 avdd.n101 avdd.n3 186.73
R3503 avdd.t4 avdd.n6 157.492
R3504 avdd.t18 avdd.n7 157.492
R3505 avdd.n25 avdd.n4 118.862
R3506 avdd.n100 avdd.n4 115.031
R3507 avdd.n73 avdd.n72 108.569
R3508 avdd.n57 avdd.n35 108.569
R3509 avdd.t9 avdd.t4 107.677
R3510 avdd.t7 avdd.t9 107.677
R3511 avdd.t7 avdd.t15 107.677
R3512 avdd.t15 avdd.t18 107.677
R3513 avdd.n62 avdd.n5 63.4672
R3514 avdd.n23 avdd.t5 60.1061
R3515 avdd.n21 avdd.n20 54.9038
R3516 avdd.n21 avdd.n19 54.9038
R3517 avdd.n72 avdd.n2 32.2138
R3518 avdd.n61 avdd.n35 32.2138
R3519 avdd.n101 avdd.n100 31.7005
R3520 avdd.n102 avdd.n101 30.3938
R3521 avdd.n76 avdd.n73 26.4291
R3522 avdd.n76 avdd.n75 26.4291
R3523 avdd.n74 avdd.n2 26.4291
R3524 avdd.n75 avdd.n74 26.4291
R3525 avdd.n78 avdd.n32 26.4291
R3526 avdd.n79 avdd.n78 26.4291
R3527 avdd.n81 avdd.n80 26.4291
R3528 avdd.n80 avdd.n79 26.4291
R3529 avdd.n58 avdd.n57 26.4291
R3530 avdd.n59 avdd.n58 26.4291
R3531 avdd.n61 avdd.n60 26.4291
R3532 avdd.n60 avdd.n59 26.4291
R3533 avdd.n54 avdd.n41 26.4291
R3534 avdd.n54 avdd.n53 26.4291
R3535 avdd.n52 avdd.n51 26.4291
R3536 avdd.n53 avdd.n52 26.4291
R3537 avdd.n96 avdd.n24 15.6997
R3538 avdd.n97 avdd.n96 14.2313
R3539 avdd.t7 avdd.n97 14.2313
R3540 avdd.n99 avdd.n98 14.2313
R3541 avdd.n98 avdd.t7 14.2313
R3542 avdd.n77 avdd.n30 13.2148
R3543 avdd.n77 avdd.t2 13.2148
R3544 avdd.n70 avdd.n31 13.2148
R3545 avdd.n70 avdd.t2 13.2148
R3546 avdd.n69 avdd.n3 13.2148
R3547 avdd.t2 avdd.n69 13.2148
R3548 avdd.n39 avdd.n38 13.2148
R3549 avdd.n39 avdd.t0 13.2148
R3550 avdd.n56 avdd.n55 13.2148
R3551 avdd.n55 avdd.t0 13.2148
R3552 avdd.n49 avdd.n37 13.2148
R3553 avdd.t0 avdd.n37 13.2148
R3554 avdd.n7 avdd.n4 12.3338
R3555 avdd.n47 avdd.n6 12.3338
R3556 avdd.n100 avdd.n99 8.13132
R3557 avdd.n95 avdd.n25 7.54184
R3558 avdd.n82 avdd.n32 7.30037
R3559 avdd.n46 avdd.n41 7.22016
R3560 avdd.n20 avdd.t10 6.92425
R3561 avdd.n20 avdd.t8 6.92425
R3562 avdd.n19 avdd.t16 6.92425
R3563 avdd.n19 avdd.t19 6.92425
R3564 avdd.n48 avdd.n47 6.88003
R3565 avdd.n99 avdd.n5 6.16704
R3566 avdd.n67 avdd.n66 3.51587
R3567 avdd.n50 avdd.n49 3.30818
R3568 avdd.n82 avdd.n81 2.8599
R3569 avdd.n90 avdd.n89 2.84665
R3570 avdd.n91 avdd.n90 2.84665
R3571 avdd.n95 avdd.n94 2.84665
R3572 avdd.n94 avdd.n93 2.84665
R3573 avdd.n51 avdd.n46 2.78239
R3574 avdd.n48 avdd.n5 2.51338
R3575 avdd.n49 avdd.n48 2.33395
R3576 avdd.n67 avdd.n27 2.28445
R3577 avdd.n92 avdd.n27 2.28445
R3578 avdd.n50 avdd.n26 2.28445
R3579 avdd.n28 avdd.n26 2.28445
R3580 avdd.n84 avdd 1.89829
R3581 avdd.n23 avdd.n22 1.87575
R3582 avdd.n102 avdd.n2 1.70717
R3583 avdd.n62 avdd.n61 1.70717
R3584 avdd.n81 avdd.n67 1.56476
R3585 avdd.n51 avdd.n50 1.54047
R3586 avdd.n85 avdd.n1 1.11161
R3587 avdd.n96 avdd.n95 1.03878
R3588 avdd.n65 avdd.n33 0.909856
R3589 avdd.n87 avdd.n65 0.871595
R3590 avdd.n42 avdd.n29 0.517167
R3591 avdd.n63 avdd.n62 0.517167
R3592 avdd.n103 avdd.n102 0.517167
R3593 avdd.n88 avdd.n87 0.517167
R3594 avdd.n83 avdd.n1 0.457832
R3595 avdd.n88 avdd.n32 0.30326
R3596 avdd.n41 avdd.n29 0.29856
R3597 avdd.n44 avdd.n34 0.277965
R3598 avdd.n44 avdd.n43 0.242141
R3599 avdd.n13 avdd.n12 0.221624
R3600 avdd.n45 avdd.n44 0.191202
R3601 avdd.n15 avdd.n8 0.171
R3602 avdd.n64 avdd 0.165618
R3603 avdd.n18 avdd.n8 0.158572
R3604 avdd.n45 avdd.n33 0.155105
R3605 avdd.n22 avdd.n18 0.129984
R3606 avdd.n65 avdd.n64 0.124867
R3607 avdd.n24 avdd.n23 0.0960224
R3608 avdd.n18 avdd.n17 0.0860931
R3609 avdd.n16 avdd.n15 0.0718577
R3610 avdd.n15 avdd.n14 0.0677409
R3611 avdd.n46 avdd.n45 0.058264
R3612 avdd.n83 avdd.n82 0.058264
R3613 avdd.n86 avdd.n85 0.0482015
R3614 avdd avdd.n63 0.0421667
R3615 avdd avdd.n0 0.035342
R3616 avdd.n12 avdd.n0 0.0293462
R3617 avdd.n22 avdd.n21 0.0285269
R3618 avdd.n17 avdd.n16 0.0255438
R3619 avdd.n14 avdd.n13 0.0253723
R3620 avdd.n12 avdd.n8 0.0246031
R3621 avdd.n85 avdd.n84 0.0240664
R3622 avdd.n11 avdd.t13 0.0122401
R3623 avdd avdd.n103 0.0122337
R3624 avdd.n17 avdd.t11 0.0122173
R3625 avdd.n10 avdd.t14 0.0113908
R3626 avdd.n9 avdd.t12 0.011362
R3627 avdd.n63 avdd.n34 0.0105575
R3628 avdd.n103 avdd.n1 0.0105575
R3629 avdd.n17 avdd.n9 0.00991802
R3630 avdd.n11 avdd.n10 0.00930403
R3631 avdd.n47 avdd.n24 0.00805162
R3632 avdd.n64 avdd 0.00600766
R3633 avdd.n43 avdd.n42 0.00573256
R3634 avdd.n42 avdd.n33 0.00515116
R3635 avdd.n87 avdd.n86 0.00333375
R3636 avdd.n14 avdd.n9 0.00220261
R3637 avdd.n16 avdd.n10 0.00176706
R3638 avdd.n84 avdd.n83 0.00111075
R3639 avdd.n64 avdd.n0 0.00109866
R3640 avdd.n13 avdd.n11 0.000671533
R3641 a_10620_n9666.t0 a_10620_n9666.t1 83.9243
R3642 a_20567_n1869.t0 a_20567_n1869.t1 198.571
R3643 a_20733_n1881.t0 a_20733_n1881.t1 60.0005
R3644 a_15539_n2791.n1 a_15539_n2791.t6 530.01
R3645 a_15539_n2791.t0 a_15539_n2791.n5 421.021
R3646 a_15539_n2791.n0 a_15539_n2791.t5 337.142
R3647 a_15539_n2791.n3 a_15539_n2791.t1 280.223
R3648 a_15539_n2791.n4 a_15539_n2791.t2 263.173
R3649 a_15539_n2791.n4 a_15539_n2791.t4 227.826
R3650 a_15539_n2791.n0 a_15539_n2791.t7 199.762
R3651 a_15539_n2791.n2 a_15539_n2791.n1 170.81
R3652 a_15539_n2791.n2 a_15539_n2791.n0 167.321
R3653 a_15539_n2791.n5 a_15539_n2791.n4 152
R3654 a_15539_n2791.n1 a_15539_n2791.t3 141.923
R3655 a_15539_n2791.n3 a_15539_n2791.n2 10.8376
R3656 a_15539_n2791.n5 a_15539_n2791.n3 2.50485
R3657 a_15705_n2791.t0 a_15705_n2791.n3 370.026
R3658 a_15705_n2791.n0 a_15705_n2791.t5 351.356
R3659 a_15705_n2791.n1 a_15705_n2791.t3 334.717
R3660 a_15705_n2791.n3 a_15705_n2791.t1 325.971
R3661 a_15705_n2791.n1 a_15705_n2791.t4 309.935
R3662 a_15705_n2791.n0 a_15705_n2791.t2 305.683
R3663 a_15705_n2791.n2 a_15705_n2791.n0 16.879
R3664 a_15705_n2791.n3 a_15705_n2791.n2 10.8867
R3665 a_15705_n2791.n2 a_15705_n2791.n1 9.3005
R3666 a_16782_n2425.t0 a_16782_n2425.t1 126.644
R3667 standby.n1 standby.t0 260.322
R3668 standby.n0 standby.t1 194.635
R3669 standby.n1 standby.t2 175.169
R3670 standby.n2 standby.n1 152
R3671 standby.n2 standby.n0 69.674
R3672 standby standby.n2 1.55726
R3673 standby.n0 standby 0.748625
R3674 a_4857_n1521.t0 a_4857_n1521.n1 405.735
R3675 a_4857_n1521.n1 a_4857_n1521.t1 294.611
R3676 a_4857_n1521.n0 a_4857_n1521.t2 254.389
R3677 a_4857_n1521.n0 a_4857_n1521.t3 211.01
R3678 a_4857_n1521.n1 a_4857_n1521.n0 152
R3679 x3.out_b.n5 x3.out_b.t8 397.163
R3680 x3.out_b.n3 x3.out_b.t4 397.163
R3681 x3.out_b.n6 x3.out_b.t8 396.286
R3682 x3.out_b.n4 x3.out_b.t4 396.286
R3683 x3.out_b.t3 x3.out_b.n5 375.649
R3684 x3.out_b.n6 x3.out_b.t3 375.649
R3685 x3.out_b.n0 x3.out_b.t6 375.649
R3686 x3.out_b.n7 x3.out_b.t6 375.649
R3687 x3.out_b.t7 x3.out_b.n3 375.649
R3688 x3.out_b.n4 x3.out_b.t7 375.649
R3689 x3.out_b.n2 x3.out_b.t0 227.887
R3690 x3.out_b.n2 x3.out_b.n8 25.0905
R3691 x3.out_b.n5 x3.out_b.n0 21.5154
R3692 x3.out_b.n3 x3.out_b.n0 21.1069
R3693 x3.out_b.n7 x3.out_b.n4 20.6372
R3694 x3.out_b.n7 x3.out_b.n6 20.6372
R3695 x3.out_b.n2 x3.out_b.t5 12.777
R3696 x3.out_b.n8 x3.out_b.t1 5.5105
R3697 x3.out_b.n8 x3.out_b.t2 5.5105
R3698 x3.out_b.n1 x3.out_b.n0 5.32901
R3699 x3.out_b.n1 x3.out_b.n7 2.74252
R3700 x3.out_b.n2 x3.out_b.n1 1.06508
R3701 a_19955_n2791.n1 a_19955_n2791.t4 530.01
R3702 a_19955_n2791.t1 a_19955_n2791.n5 421.021
R3703 a_19955_n2791.n0 a_19955_n2791.t3 337.142
R3704 a_19955_n2791.n3 a_19955_n2791.t0 280.223
R3705 a_19955_n2791.n4 a_19955_n2791.t6 263.173
R3706 a_19955_n2791.n4 a_19955_n2791.t2 227.826
R3707 a_19955_n2791.n0 a_19955_n2791.t5 199.762
R3708 a_19955_n2791.n2 a_19955_n2791.n1 170.81
R3709 a_19955_n2791.n2 a_19955_n2791.n0 167.321
R3710 a_19955_n2791.n5 a_19955_n2791.n4 152
R3711 a_19955_n2791.n1 a_19955_n2791.t7 141.923
R3712 a_19955_n2791.n3 a_19955_n2791.n2 10.8376
R3713 a_19955_n2791.n5 a_19955_n2791.n3 2.50485
R3714 a_20121_n2791.t0 a_20121_n2791.n3 370.026
R3715 a_20121_n2791.n0 a_20121_n2791.t4 351.356
R3716 a_20121_n2791.n1 a_20121_n2791.t3 334.717
R3717 a_20121_n2791.n3 a_20121_n2791.t1 325.971
R3718 a_20121_n2791.n1 a_20121_n2791.t2 309.935
R3719 a_20121_n2791.n0 a_20121_n2791.t5 305.683
R3720 a_20121_n2791.n2 a_20121_n2791.n0 16.879
R3721 a_20121_n2791.n3 a_20121_n2791.n2 10.8867
R3722 a_20121_n2791.n2 a_20121_n2791.n1 9.3005
R3723 a_19567_n2247.t1 a_19567_n2247.n1 386.31
R3724 a_19567_n2247.n1 a_19567_n2247.t0 249.956
R3725 a_19567_n2247.n0 a_19567_n2247.t3 239.04
R3726 a_19567_n2247.n1 a_19567_n2247.n0 175.661
R3727 a_19567_n2247.n0 a_19567_n2247.t2 166.739
R3728 ena.n0 ena.t2 260.322
R3729 ena.n2 ena.t0 194.63
R3730 ena.n0 ena.t1 175.169
R3731 ena.n1 ena.n0 152
R3732 ena.n3 ena.n2 51.6747
R3733 ena ena.n3 4.94983
R3734 ena.n3 ena.n1 3.45996
R3735 ena.n1 ena 1.55726
R3736 ena.n2 ena 0.746125
R3737 a_19003_n2817.n6 a_19003_n2817.n5 746.659
R3738 a_19003_n2817.n0 a_19003_n2817.t5 389.183
R3739 a_19003_n2817.n2 a_19003_n2817.t3 256.988
R3740 a_19003_n2817.n1 a_19003_n2817.n0 251.167
R3741 a_19003_n2817.n1 a_19003_n2817.t2 223.571
R3742 a_19003_n2817.n4 a_19003_n2817.t8 212.081
R3743 a_19003_n2817.n5 a_19003_n2817.n4 181.942
R3744 a_19003_n2817.n0 a_19003_n2817.t4 174.891
R3745 a_19003_n2817.n2 a_19003_n2817.t6 163.803
R3746 a_19003_n2817.n3 a_19003_n2817.t7 139.78
R3747 a_19003_n2817.n3 a_19003_n2817.n2 129.264
R3748 a_19003_n2817.n6 a_19003_n2817.t1 63.3219
R3749 a_19003_n2817.t0 a_19003_n2817.n6 63.3219
R3750 a_19003_n2817.n5 a_19003_n2817.n1 24.6993
R3751 a_19003_n2817.n4 a_19003_n2817.n3 22.6399
R3752 a_19567_n2791.t0 a_19567_n2791.n1 386.31
R3753 a_19567_n2791.n1 a_19567_n2791.t1 249.956
R3754 a_19567_n2791.n0 a_19567_n2791.t3 239.04
R3755 a_19567_n2791.n1 a_19567_n2791.n0 175.661
R3756 a_19567_n2791.n0 a_19567_n2791.t2 166.739
R3757 vg1.n10 vg1.t1 85.228
R3758 vg1.n0 vg1.t3 61.1305
R3759 vg1.n7 vg1.t5 54.828
R3760 vg1.n7 vg1.t1 54.828
R3761 vg1.n5 vg1.t0 42.6599
R3762 vg1.n8 vg1.n7 32.9015
R3763 vg1.n10 vg1.n9 30.9745
R3764 vg1.n9 vg1.t2 20.9512
R3765 vg1.n6 vg1.n5 3.63479
R3766 vg1.n11 vg1.n10 2.3255
R3767 vg1.n12 vg1.n0 0.471594
R3768 vg1.n5 vg1.n4 0.390524
R3769 vg1.n9 vg1.n8 0.238607
R3770 vg1.n11 vg1.n6 0.176742
R3771 vg1 vg1.n12 0.133236
R3772 vg1.n1 vg1.t9 0.0767969
R3773 vg1.n2 vg1.n1 0.0752537
R3774 vg1.n3 vg1.n2 0.0752537
R3775 vg1.n4 vg1.t8 0.0717511
R3776 vg1.n0 vg1 0.0387813
R3777 vg1.n12 vg1.n11 0.0257152
R3778 vg1.n8 vg1.n6 0.0123355
R3779 vg1.n4 vg1.n3 0.00554581
R3780 vg1.n1 vg1.t4 0.00204321
R3781 vg1.n2 vg1.t7 0.00204321
R3782 vg1.n3 vg1.t6 0.00204321
R3783 a_21145_n1869.n0 a_21145_n1869.t0 68.3338
R3784 a_21145_n1869.n0 a_21145_n1869.t1 26.3935
R3785 a_21145_n1869.n1 a_21145_n1869.n0 14.4005
R3786 a_21211_n2817.n4 a_21211_n2817.n0 746.659
R3787 a_21211_n2817.n5 a_21211_n2817.t8 389.183
R3788 a_21211_n2817.n1 a_21211_n2817.t6 256.988
R3789 a_21211_n2817.n6 a_21211_n2817.n5 251.167
R3790 a_21211_n2817.t0 a_21211_n2817.n6 223.571
R3791 a_21211_n2817.n3 a_21211_n2817.t5 212.081
R3792 a_21211_n2817.n4 a_21211_n2817.n3 181.942
R3793 a_21211_n2817.n5 a_21211_n2817.t7 174.891
R3794 a_21211_n2817.n1 a_21211_n2817.t3 163.803
R3795 a_21211_n2817.n2 a_21211_n2817.t4 139.78
R3796 a_21211_n2817.n2 a_21211_n2817.n1 129.264
R3797 a_21211_n2817.n0 a_21211_n2817.t1 63.3219
R3798 a_21211_n2817.n0 a_21211_n2817.t2 63.3219
R3799 a_21211_n2817.n6 a_21211_n2817.n4 24.6993
R3800 a_21211_n2817.n3 a_21211_n2817.n2 22.6399
R3801 xin.n36 xin.t8 594.832
R3802 xin.t18 xin.n5 380.808
R3803 xin.n6 xin.t18 380.808
R3804 xin.n6 xin.t15 380.611
R3805 xin.t15 xin.n5 380.611
R3806 xin.t13 xin.n7 380.611
R3807 xin.n8 xin.t13 380.611
R3808 xin.t19 xin.n4 380.611
R3809 xin.n9 xin.t19 380.611
R3810 xin.n11 xin.t16 380.611
R3811 xin.t16 xin.n10 380.611
R3812 xin.n12 xin.t11 380.611
R3813 xin.t11 xin.n3 380.611
R3814 xin.t10 xin.n13 380.611
R3815 xin.n14 xin.t10 380.611
R3816 xin.t17 xin.n2 380.611
R3817 xin.n15 xin.t17 380.611
R3818 xin.n17 xin.t14 380.611
R3819 xin.t14 xin.n16 380.611
R3820 xin.n18 xin.t12 380.611
R3821 xin.t12 xin.n1 380.611
R3822 xin.t9 xin.n19 380.611
R3823 xin.n20 xin.t9 380.611
R3824 xin.n21 xin.t6 380.611
R3825 xin.t6 xin.n0 380.611
R3826 xin.n36 xin.t21 194.639
R3827 xin.n25 xin.t20 124.457
R3828 xin.n25 xin.t7 106.793
R3829 xin.t7 xin.n23 86.3125
R3830 xin.t20 xin.n24 86.3125
R3831 xin.n24 xin.n23 58.6245
R3832 xin.n30 xin.t0 45.927
R3833 xin.n28 xin.n27 20.1298
R3834 xin.n27 xin.n23 12.2455
R3835 xin.n35 xin.n34 4.04311
R3836 xin.n26 xin.n24 3.56553
R3837 xin.n34 xin.n29 3.51336
R3838 xin.n30 xin.n29 3.51061
R3839 xin.n28 xin.n22 1.95915
R3840 xin.n35 xin.n28 1.1106
R3841 xin.n22 xin.n21 0.8105
R3842 xin.n22 xin.n0 0.7905
R3843 xin.n27 xin.n26 0.741791
R3844 xin.n26 xin.n25 0.715885
R3845 xin.n36 xin.n35 0.4755
R3846 xin xin.n36 0.377063
R3847 xin.n8 xin.n5 0.198
R3848 xin.n9 xin.n8 0.198
R3849 xin.n10 xin.n9 0.198
R3850 xin.n10 xin.n3 0.198
R3851 xin.n14 xin.n3 0.198
R3852 xin.n15 xin.n14 0.198
R3853 xin.n16 xin.n15 0.198
R3854 xin.n16 xin.n1 0.198
R3855 xin.n20 xin.n1 0.198
R3856 xin.n21 xin.n20 0.198
R3857 xin.n7 xin.n6 0.198
R3858 xin.n7 xin.n4 0.198
R3859 xin.n11 xin.n4 0.198
R3860 xin.n12 xin.n11 0.198
R3861 xin.n13 xin.n12 0.198
R3862 xin.n13 xin.n2 0.198
R3863 xin.n17 xin.n2 0.198
R3864 xin.n18 xin.n17 0.198
R3865 xin.n19 xin.n18 0.198
R3866 xin.n19 xin.n0 0.198
R3867 xin.t4 xin.t2 0.0760058
R3868 xin.n31 xin.n30 0.0410952
R3869 xin.n32 xin.n29 0.0410952
R3870 xin.n34 xin.n33 0.0410952
R3871 xin.n32 xin.t5 0.0264927
R3872 xin.n31 xin.t1 0.0264885
R3873 xin.n33 xin.t4 0.0264703
R3874 xin.n33 xin.t3 0.0264296
R3875 xin.t3 xin.n32 0.0264114
R3876 xin.t5 xin.n31 0.0264072
R3877 a_19182_n2791.t0 a_19182_n2791.t1 87.1434
R3878 a_2132_n17250.t0 a_2132_n17250.t1 82.3314
R3879 a_24220_n9500.t0 a_24220_n9500.t1 83.56
R3880 a_17913_n2241.t1 a_17913_n2241.n3 370.026
R3881 a_17913_n2241.n0 a_17913_n2241.t3 351.356
R3882 a_17913_n2241.n1 a_17913_n2241.t2 334.717
R3883 a_17913_n2241.n3 a_17913_n2241.t0 325.971
R3884 a_17913_n2241.n1 a_17913_n2241.t4 309.935
R3885 a_17913_n2241.n0 a_17913_n2241.t5 305.683
R3886 a_17913_n2241.n2 a_17913_n2241.n0 16.879
R3887 a_17913_n2241.n3 a_17913_n2241.n2 10.8867
R3888 a_17913_n2241.n2 a_17913_n2241.n1 9.3005
R3889 a_18263_n1869.n3 a_18263_n1869.n2 674.338
R3890 a_18263_n1869.n1 a_18263_n1869.t4 332.58
R3891 a_18263_n1869.n2 a_18263_n1869.n0 284.012
R3892 a_18263_n1869.n2 a_18263_n1869.n1 253.648
R3893 a_18263_n1869.n1 a_18263_n1869.t5 168.701
R3894 a_18263_n1869.t0 a_18263_n1869.n3 96.1553
R3895 a_18263_n1869.n3 a_18263_n1869.t1 65.6672
R3896 a_18263_n1869.n0 a_18263_n1869.t3 65.0005
R3897 a_18263_n1869.n0 a_18263_n1869.t2 45.0005
R3898 a_18359_n1869.t1 a_18359_n1869.t0 198.571
R3899 vg2.n2 vg2.t9 87.8852
R3900 vg2.n9 vg2.t5 87.8852
R3901 vg2.n5 vg2.t6 85.228
R3902 vg2.n12 vg2.t7 85.228
R3903 vg2.n15 vg2.t8 67.0783
R3904 vg2.n4 vg2.t9 54.828
R3905 vg2.t6 vg2.n4 54.828
R3906 vg2.n11 vg2.t5 54.828
R3907 vg2.t7 vg2.n11 54.828
R3908 vg2.n16 vg2.t4 42.6015
R3909 vg2.n4 vg2.n3 30.4005
R3910 vg2.n11 vg2.n10 30.4005
R3911 vg2.n3 vg2.n1 29.1205
R3912 vg2.n5 vg2.n1 29.1205
R3913 vg2.n10 vg2.n8 29.1205
R3914 vg2.n12 vg2.n8 29.1205
R3915 vg2.n6 vg2.n5 2.3255
R3916 vg2.n13 vg2.n12 2.3255
R3917 vg2.n3 vg2.n2 2.13477
R3918 vg2.n10 vg2.n9 2.13477
R3919 vg2 vg2.n14 0.742464
R3920 vg2.n16 vg2.n15 0.714193
R3921 vg2.n14 vg2.n6 0.474719
R3922 vg2.n14 vg2.n13 0.474719
R3923 vg2.n1 vg2.n0 0.423227
R3924 vg2.n8 vg2.n7 0.423227
R3925 vg2.n2 vg2.n0 0.308459
R3926 vg2.n9 vg2.n7 0.308459
R3927 vg2.n6 vg2.n0 0.284875
R3928 vg2.n13 vg2.n7 0.284875
R3929 vg2.n15 vg2.t2 0.170134
R3930 vg2 vg2.n16 0.119455
R3931 vg2.t0 vg2.t1 0.0652716
R3932 vg2.t3 vg2.t0 0.0652716
R3933 vg2.t2 vg2.t3 0.0652716
R3934 vrb.n2 vrb.t0 43.1048
R3935 vrb.n0 vrb.t4 22.3777
R3936 vrb.n1 vrb.t1 22.1989
R3937 vrb.n1 vrb.t3 21.3671
R3938 vrb.n0 vrb.t2 21.3663
R3939 vrb.n3 vrb.n2 1.11856
R3940 vrb.n3 vrb.n0 0.759192
R3941 vrb.n2 vrb.n1 0.758408
R3942 vrb vrb.n3 0.0491111
R3943 a_18359_n2791.t0 a_18359_n2791.t1 198.571
R3944 a_18525_n2791.t0 a_18525_n2791.t1 60.0005
R3945 a_2130_n20844.t0 a_2130_n20844.t1 82.0028
R3946 a_24530_n21010.t0 a_24530_n21010.t1 81.9478
R3947 a_15083_n2791.t0 a_15083_n2791.t1 60.0005
R3948 a_18932_n15424.t0 a_18932_n15424.t1 83.5579
R3949 a_14285_n2281.n1 a_14285_n2281.n0 953.039
R3950 a_14285_n2281.t0 a_14285_n2281.n1 33.4905
R3951 a_14285_n2281.n1 a_14285_n2281.t1 31.5205
R3952 a_14285_n2281.n0 a_14285_n2281.t3 26.5955
R3953 a_14285_n2281.n0 a_14285_n2281.t2 26.5955
R3954 a_14285_n2079.t0 a_14285_n2079.n0 1201.3
R3955 a_14285_n2079.n0 a_14285_n2079.t2 26.5955
R3956 a_14285_n2079.n0 a_14285_n2079.t1 26.5955
R3957 a_18828_n1869.n3 a_18828_n1869.n2 636.953
R3958 a_18828_n1869.n1 a_18828_n1869.t4 366.856
R3959 a_18828_n1869.n2 a_18828_n1869.n0 300.2
R3960 a_18828_n1869.n2 a_18828_n1869.n1 225.036
R3961 a_18828_n1869.n1 a_18828_n1869.t5 174.056
R3962 a_18828_n1869.n0 a_18828_n1869.t1 70.0005
R3963 a_18828_n1869.n3 a_18828_n1869.t3 68.0124
R3964 a_18828_n1869.t0 a_18828_n1869.n3 63.3219
R3965 a_18828_n1869.n0 a_18828_n1869.t2 61.6672
R3966 a_19182_n1881.t0 a_19182_n1881.t1 87.1434
R3967 a_19003_n1943.n6 a_19003_n1943.n5 746.659
R3968 a_19003_n1943.n0 a_19003_n1943.t8 389.183
R3969 a_19003_n1943.n2 a_19003_n1943.t5 256.988
R3970 a_19003_n1943.n1 a_19003_n1943.n0 251.167
R3971 a_19003_n1943.n1 a_19003_n1943.t2 223.571
R3972 a_19003_n1943.n4 a_19003_n1943.t7 212.081
R3973 a_19003_n1943.n5 a_19003_n1943.n4 181.942
R3974 a_19003_n1943.n0 a_19003_n1943.t3 174.891
R3975 a_19003_n1943.n2 a_19003_n1943.t6 163.803
R3976 a_19003_n1943.n3 a_19003_n1943.t4 139.78
R3977 a_19003_n1943.n3 a_19003_n1943.n2 129.264
R3978 a_19003_n1943.n6 a_19003_n1943.t1 63.3219
R3979 a_19003_n1943.t0 a_19003_n1943.n6 63.3219
R3980 a_19003_n1943.n5 a_19003_n1943.n1 24.6993
R3981 a_19003_n1943.n4 a_19003_n1943.n3 22.6399
R3982 vn.t9 vn.n3 182.935
R3983 vn.t2 vn.n0 144.126
R3984 vn.n8 vn.n5 97.2442
R3985 vn.n9 vn.n3 97.2442
R3986 vn.n4 vn.t9 88.2031
R3987 vn.t8 vn.n3 85.228
R3988 vn.n5 vn.t8 85.228
R3989 vn.n9 vn.t0 85.228
R3990 vn.t0 vn.n8 85.228
R3991 vn.n1 vn.t2 85.228
R3992 vn vn.t6 64.2147
R3993 vn.n7 vn.n1 58.8987
R3994 vn vn.n2 56.3112
R3995 vn vn.t4 21.1687
R3996 vn.n8 vn.n7 17.975
R3997 vn.n9 vn.n0 17.975
R3998 vn vn.n6 16.8187
R3999 vn.n2 vn.t7 6.92425
R4000 vn.n2 vn.t5 6.92425
R4001 vn.n6 vn.t1 4.3505
R4002 vn.n6 vn.t3 4.3505
R4003 vn.n4 vn 3.29454
R4004 vn vn.n1 2.80102
R4005 vn.n8 vn 2.44682
R4006 vn.n3 vn 2.3255
R4007 vn vn.n9 2.3255
R4008 vn.n5 vn.n4 2.20282
R4009 vn.n7 vn 2.69718
R4010 vn vn.n0 2.67028
R4011 a_10620_n7674.t0 a_10620_n7674.t1 82.5973
R4012 a_24220_n7840.t0 a_24220_n7840.t1 83.56
R4013 x7.x2.Qb1.n4 x7.x2.Qb1.t0 372.361
R4014 x7.x2.Qb1.n2 x7.x2.Qb1.t5 333.651
R4015 x7.x2.Qb1.n2 x7.x2.Qb1.t2 297.233
R4016 x7.x2.Qb1.n1 x7.x2.Qb1.t3 294.557
R4017 x7.x2.Qb1.n5 x7.x2.Qb1.t1 231.921
R4018 x7.x2.Qb1.n1 x7.x2.Qb1.t4 211.01
R4019 x7.x2.Qb1 x7.x2.Qb1.n2 195.701
R4020 x7.x2.Qb1.n0 x7.x2.Qb1.n1 152
R4021 x7.x2.Qb1.n5 x7.x2.Qb1.n0 40.9605
R4022 x7.x2.Qb1.n5 x7.x2.Qb1.n4 18.1966
R4023 x7.x2.Qb1.n0 x7.x2.Qb1 10.4234
R4024 x7.x2.Qb1.n4 x7.x2.Qb1.n3 9.35675
R4025 x7.x2.Qb1.n3 x7.x2.Qb1 6.49269
R4026 x7.x2.Qb1.n3 x7.x2.Qb1 3.52967
R4027 x7.x2.Qb1 x7.x2.Qb1.n5 2.5605
R4028 x7.x2.Qb1.n0 x7.x2.Qb1 2.01193
R4029 a_15960_n2791.n1 a_15960_n2791.n0 926.024
R4030 a_15960_n2791.n1 a_15960_n2791.t3 82.0838
R4031 a_15960_n2791.n0 a_15960_n2791.t0 63.3338
R4032 a_15960_n2791.t1 a_15960_n2791.n1 63.3219
R4033 a_15960_n2791.n0 a_15960_n2791.t2 29.7268
R4034 a_2130_n19516.t0 a_2130_n19516.t1 82.0028
R4035 a_24530_n19682.t0 a_24530_n19682.t1 81.9478
R4036 a_20579_n2247.n0 a_20579_n2247.t1 1327.82
R4037 a_20579_n2247.n0 a_20579_n2247.t2 194.655
R4038 a_20579_n2247.t0 a_20579_n2247.n0 63.3219
R4039 a_15083_n1881.t0 a_15083_n1881.t1 60.0005
R4040 a_18481_n2273.n3 a_18481_n2273.n2 647.119
R4041 a_18481_n2273.n1 a_18481_n2273.t4 350.253
R4042 a_18481_n2273.n2 a_18481_n2273.n0 260.339
R4043 a_18481_n2273.n2 a_18481_n2273.n1 246.119
R4044 a_18481_n2273.n1 a_18481_n2273.t5 189.588
R4045 a_18481_n2273.n3 a_18481_n2273.t3 89.1195
R4046 a_18481_n2273.n0 a_18481_n2273.t0 63.3338
R4047 a_18481_n2273.t1 a_18481_n2273.n3 41.0422
R4048 a_18481_n2273.n0 a_18481_n2273.t2 31.9797
R4049 a_18525_n1881.t0 a_18525_n1881.t1 60.0005
R4050 x7.x2.Qb2.n4 x7.x2.Qb2.t0 372.361
R4051 x7.x2.Qb2.n2 x7.x2.Qb2.t5 333.651
R4052 x7.x2.Qb2.n2 x7.x2.Qb2.t2 297.233
R4053 x7.x2.Qb2.n1 x7.x2.Qb2.t3 294.557
R4054 x7.x2.Qb2.n5 x7.x2.Qb2.t1 231.921
R4055 x7.x2.Qb2.n1 x7.x2.Qb2.t4 211.01
R4056 x7.x2.Qb2 x7.x2.Qb2.n2 195.701
R4057 x7.x2.Qb2.n0 x7.x2.Qb2.n1 152
R4058 x7.x2.Qb2.n5 x7.x2.Qb2.n0 40.9605
R4059 x7.x2.Qb2.n5 x7.x2.Qb2.n4 18.1966
R4060 x7.x2.Qb2.n0 x7.x2.Qb2 10.4234
R4061 x7.x2.Qb2.n4 x7.x2.Qb2.n3 9.36092
R4062 x7.x2.Qb2.n3 x7.x2.Qb2 6.49269
R4063 x7.x2.Qb2.n3 x7.x2.Qb2 3.52967
R4064 x7.x2.Qb2 x7.x2.Qb2.n5 2.5605
R4065 x7.x2.Qb2.n0 x7.x2.Qb2 2.01193
R4066 a_18168_n2791.n1 a_18168_n2791.n0 926.024
R4067 a_18168_n2791.n1 a_18168_n2791.t3 82.0838
R4068 a_18168_n2791.n0 a_18168_n2791.t0 63.3338
R4069 a_18168_n2791.t1 a_18168_n2791.n1 63.3219
R4070 a_18168_n2791.n0 a_18168_n2791.t2 29.7268
R4071 a_16055_n2791.n3 a_16055_n2791.n2 674.338
R4072 a_16055_n2791.n1 a_16055_n2791.t4 332.58
R4073 a_16055_n2791.n2 a_16055_n2791.n0 284.012
R4074 a_16055_n2791.n2 a_16055_n2791.n1 253.648
R4075 a_16055_n2791.n1 a_16055_n2791.t5 168.701
R4076 a_16055_n2791.t0 a_16055_n2791.n3 96.1553
R4077 a_16055_n2791.n3 a_16055_n2791.t2 65.6672
R4078 a_16055_n2791.n0 a_16055_n2791.t1 65.0005
R4079 a_16055_n2791.n0 a_16055_n2791.t3 45.0005
R4080 x7.x1.x4.Q x7.x1.x4.Q.t0 240.05
R4081 x7.x1.x4.Q x7.x1.x4.Q.t1 155.386
R4082 a_14009_n2404.t2 a_14009_n2404.n3 669.389
R4083 a_14009_n2404.n0 a_14009_n2404.t3 326.493
R4084 a_14009_n2404.n0 a_14009_n2404.t1 249.615
R4085 a_14009_n2404.n1 a_14009_n2404.t0 249.615
R4086 a_14009_n2404.n2 a_14009_n2404.t4 241.536
R4087 a_14009_n2404.n2 a_14009_n2404.t5 169.237
R4088 a_14009_n2404.n3 a_14009_n2404.n2 152
R4089 a_14009_n2404.n3 a_14009_n2404.n1 108.529
R4090 a_14009_n2404.n1 a_14009_n2404.n0 26.6245
R4091 a_24530_n20678.t0 a_24530_n20678.t1 81.9478
R4092 a_15539_n2241.n1 a_15539_n2241.t5 530.01
R4093 a_15539_n2241.t0 a_15539_n2241.n5 421.021
R4094 a_15539_n2241.n0 a_15539_n2241.t3 337.142
R4095 a_15539_n2241.n3 a_15539_n2241.t1 280.223
R4096 a_15539_n2241.n4 a_15539_n2241.t4 263.173
R4097 a_15539_n2241.n4 a_15539_n2241.t6 227.826
R4098 a_15539_n2241.n0 a_15539_n2241.t2 199.762
R4099 a_15539_n2241.n2 a_15539_n2241.n1 170.81
R4100 a_15539_n2241.n2 a_15539_n2241.n0 167.321
R4101 a_15539_n2241.n5 a_15539_n2241.n4 152
R4102 a_15539_n2241.n1 a_15539_n2241.t7 141.923
R4103 a_15539_n2241.n3 a_15539_n2241.n2 10.8376
R4104 a_15539_n2241.n5 a_15539_n2241.n3 2.50485
R4105 a_16729_n1869.n0 a_16729_n1869.t1 68.3338
R4106 a_16729_n1869.n0 a_16729_n1869.t0 26.3935
R4107 a_16729_n1869.n1 a_16729_n1869.n0 14.4005
R4108 a_16055_n1869.n3 a_16055_n1869.n2 674.338
R4109 a_16055_n1869.n1 a_16055_n1869.t4 332.58
R4110 a_16055_n1869.n2 a_16055_n1869.n0 284.012
R4111 a_16055_n1869.n2 a_16055_n1869.n1 253.648
R4112 a_16055_n1869.n1 a_16055_n1869.t5 168.701
R4113 a_16055_n1869.t0 a_16055_n1869.n3 96.1553
R4114 a_16055_n1869.n3 a_16055_n1869.t2 65.6672
R4115 a_16055_n1869.n0 a_16055_n1869.t1 65.0005
R4116 a_16055_n1869.n0 a_16055_n1869.t3 45.0005
R4117 a_2132_n15258.t0 a_2132_n15258.t1 83.9223
R4118 a_18990_n2425.t0 a_18990_n2425.t1 126.644
R4119 a_24530_n19350.t0 a_24530_n19350.t1 81.9478
R4120 a_16163_n2247.t0 a_16163_n2247.n0 1327.82
R4121 a_16163_n2247.n0 a_16163_n2247.t2 194.655
R4122 a_16163_n2247.n0 a_16163_n2247.t1 63.3219
R4123 a_2132_n16918.t0 a_2132_n16918.t1 82.3314
R4124 a_18932_n17084.t0 a_18932_n17084.t1 83.5579
R4125 a_10620_n9334.t0 a_10620_n9334.t1 83.9243
R4126 a_3134_n13324.t0 a_3134_n13324.t1 83.9223
R4127 x7.x1.x2.Q x7.x1.x2.Q.t0 240.05
R4128 x7.x1.x2.Q x7.x1.x2.Q.t1 155.386
R4129 a_18932_n17748.t0 a_18932_n17748.t1 83.5579
R4130 a_18937_n2791.t0 a_18937_n2791.t1 94.7268
R4131 x3.out.n3 x3.out.t6 393.144
R4132 x3.out.n5 x3.out.t7 393.144
R4133 x3.out.n4 x3.out.t6 391.815
R4134 x3.out.t7 x3.out.n2 391.815
R4135 x3.out.n5 x3.out.t4 371.31
R4136 x3.out.t4 x3.out.n2 371.31
R4137 x3.out.t3 x3.out.n1 371.31
R4138 x3.out.n6 x3.out.t3 371.31
R4139 x3.out.n4 x3.out.t8 371.31
R4140 x3.out.t8 x3.out.n3 371.31
R4141 x3.out.n0 x3.out.t2 227.886
R4142 x3.out.n0 x3.out.n9 25.0903
R4143 x3.out.n1 x3.out.n5 21.8335
R4144 x3.out.n3 x3.out.n1 21.6959
R4145 x3.out.n6 x3.out.n4 20.5053
R4146 x3.out.n7 x3.out.n2 19.6003
R4147 x3.out.n0 x3.out.t5 12.7763
R4148 x3.out.n9 x3.out.t0 5.5105
R4149 x3.out.n9 x3.out.t1 5.5105
R4150 x3.out.n8 x3.out.n1 5.0449
R4151 x3.out.n8 x3.out.n7 2.71826
R4152 x3.out.n7 x3.out.n6 0.90555
R4153 x3.out x3.out.n8 0.88175
R4154 x3.out x3.out.n0 0.794875
R4155 a_17359_n2247.t0 a_17359_n2247.n1 386.31
R4156 a_17359_n2247.n1 a_17359_n2247.t1 249.956
R4157 a_17359_n2247.n0 a_17359_n2247.t2 239.04
R4158 a_17359_n2247.n1 a_17359_n2247.n0 175.661
R4159 a_17359_n2247.n0 a_17359_n2247.t3 166.739
R4160 a_24530_n22338.t0 a_24530_n22338.t1 81.9492
R4161 dout_filt.n0 dout_filt.t2 687.288
R4162 x7.clkout dout_filt.t0 229.845
R4163 dout_filt.n1 dout_filt.t1 223.571
R4164 dout_filt.n1 dout_filt.n0 139.672
R4165 dout_filt.n2 dout_filt.t4 97.4114
R4166 dout_filt.n2 dout_filt.t3 56.9639
R4167 x7.clkout x7.x5.Z 28.6323
R4168 x7.x5.Z x7.clkout 28.3622
R4169 x7.clkout dout_filt.n2 10.5187
R4170 x7.x5.Z dout_filt.n1 4.70638
R4171 x7.x5.Z dout_filt.n0 4.70638
R4172 x4.out_b.n0 x4.out_b.t0 227.887
R4173 x4.out_b.n0 x4.out_b.n1 25.0905
R4174 x4.out_b.n0 x4.out_b.t3 12.777
R4175 x4.out_b.n1 x4.out_b.t1 5.5105
R4176 x4.out_b.n1 x4.out_b.t2 5.5105
R4177 x4.out_b x4.out_b.n0 0.83175
R4178 a_15960_n1881.n1 a_15960_n1881.n0 926.024
R4179 a_15960_n1881.n0 a_15960_n1881.t3 82.0838
R4180 a_15960_n1881.n1 a_15960_n1881.t2 63.3338
R4181 a_15960_n1881.n0 a_15960_n1881.t1 63.3219
R4182 a_15960_n1881.t0 a_15960_n1881.n1 29.7268
R4183 a_20471_n2791.n3 a_20471_n2791.n2 674.338
R4184 a_20471_n2791.n1 a_20471_n2791.t5 332.58
R4185 a_20471_n2791.n2 a_20471_n2791.n0 284.012
R4186 a_20471_n2791.n2 a_20471_n2791.n1 253.648
R4187 a_20471_n2791.n1 a_20471_n2791.t4 168.701
R4188 a_20471_n2791.t0 a_20471_n2791.n3 96.1553
R4189 a_20471_n2791.n3 a_20471_n2791.t2 65.6672
R4190 a_20471_n2791.n0 a_20471_n2791.t1 65.0005
R4191 a_20471_n2791.n0 a_20471_n2791.t3 45.0005
R4192 a_24220_n9168.t0 a_24220_n9168.t1 83.56
R4193 a_21036_n2791.n3 a_21036_n2791.n2 636.953
R4194 a_21036_n2791.n1 a_21036_n2791.t5 366.856
R4195 a_21036_n2791.n2 a_21036_n2791.n0 300.2
R4196 a_21036_n2791.n2 a_21036_n2791.n1 225.036
R4197 a_21036_n2791.n1 a_21036_n2791.t4 174.056
R4198 a_21036_n2791.n0 a_21036_n2791.t3 70.0005
R4199 a_21036_n2791.t1 a_21036_n2791.n3 68.0124
R4200 a_21036_n2791.n3 a_21036_n2791.t2 63.3219
R4201 a_21036_n2791.n0 a_21036_n2791.t0 61.6672
R4202 a_18937_n1869.n0 a_18937_n1869.t0 68.3338
R4203 a_18937_n1869.n0 a_18937_n1869.t1 26.3935
R4204 a_18937_n1869.n1 a_18937_n1869.n0 14.4005
R4205 a_17747_n2791.n1 a_17747_n2791.t7 530.01
R4206 a_17747_n2791.t0 a_17747_n2791.n5 421.021
R4207 a_17747_n2791.n0 a_17747_n2791.t6 337.142
R4208 a_17747_n2791.n3 a_17747_n2791.t1 280.223
R4209 a_17747_n2791.n4 a_17747_n2791.t3 263.173
R4210 a_17747_n2791.n4 a_17747_n2791.t5 227.826
R4211 a_17747_n2791.n0 a_17747_n2791.t2 199.762
R4212 a_17747_n2791.n2 a_17747_n2791.n1 170.81
R4213 a_17747_n2791.n2 a_17747_n2791.n0 167.321
R4214 a_17747_n2791.n5 a_17747_n2791.n4 152
R4215 a_17747_n2791.n1 a_17747_n2791.t4 141.923
R4216 a_17747_n2791.n3 a_17747_n2791.n2 10.8376
R4217 a_17747_n2791.n5 a_17747_n2791.n3 2.50485
R4218 a_17359_n2791.t0 a_17359_n2791.n1 386.31
R4219 a_17359_n2791.n1 a_17359_n2791.t1 249.956
R4220 a_17359_n2791.n0 a_17359_n2791.t3 239.04
R4221 a_17359_n2791.n1 a_17359_n2791.n0 175.661
R4222 a_17359_n2791.n0 a_17359_n2791.t2 166.739
R4223 a_2130_n20512.t0 a_2130_n20512.t1 82.0028
R4224 a_18263_n2791.n3 a_18263_n2791.n2 674.338
R4225 a_18263_n2791.n1 a_18263_n2791.t4 332.58
R4226 a_18263_n2791.n2 a_18263_n2791.n0 284.012
R4227 a_18263_n2791.n2 a_18263_n2791.n1 253.648
R4228 a_18263_n2791.n1 a_18263_n2791.t5 168.701
R4229 a_18263_n2791.t1 a_18263_n2791.n3 96.1553
R4230 a_18263_n2791.n3 a_18263_n2791.t2 65.6672
R4231 a_18263_n2791.n0 a_18263_n2791.t0 65.0005
R4232 a_18263_n2791.n0 a_18263_n2791.t3 45.0005
R4233 a_2132_n14926.t0 a_2132_n14926.t1 83.9223
R4234 a_18932_n15092.t0 a_18932_n15092.t1 83.5579
R4235 a_14357_n2743.t0 a_14357_n2743.t1 64.6411
R4236 dout.n0 dout.t0 120.561
R4237 dout.n0 dout.t1 61.4115
R4238 dout dout.n0 3.88384
R4239 a_20376_n1881.n1 a_20376_n1881.n0 926.024
R4240 a_20376_n1881.n1 a_20376_n1881.t3 82.0838
R4241 a_20376_n1881.n0 a_20376_n1881.t0 63.3338
R4242 a_20376_n1881.t1 a_20376_n1881.n1 63.3219
R4243 a_20376_n1881.n0 a_20376_n1881.t2 29.7268
R4244 a_20471_n1869.n3 a_20471_n1869.n2 674.338
R4245 a_20471_n1869.n1 a_20471_n1869.t5 332.58
R4246 a_20471_n1869.n2 a_20471_n1869.n0 284.012
R4247 a_20471_n1869.n2 a_20471_n1869.n1 253.648
R4248 a_20471_n1869.n1 a_20471_n1869.t4 168.701
R4249 a_20471_n1869.t1 a_20471_n1869.n3 96.1553
R4250 a_20471_n1869.n3 a_20471_n1869.t3 65.6672
R4251 a_20471_n1869.n0 a_20471_n1869.t0 65.0005
R4252 a_20471_n1869.n0 a_20471_n1869.t2 45.0005
R4253 x7.x1.Qb1.n4 x7.x1.Qb1.t0 372.361
R4254 x7.x1.Qb1.n2 x7.x1.Qb1.t4 333.651
R4255 x7.x1.Qb1.n2 x7.x1.Qb1.t5 297.233
R4256 x7.x1.Qb1.n0 x7.x1.Qb1.t2 294.557
R4257 x7.x1.Qb1.n5 x7.x1.Qb1.t1 231.921
R4258 x7.x1.Qb1.n0 x7.x1.Qb1.t3 211.01
R4259 x7.x1.Qb1 x7.x1.Qb1.n2 195.701
R4260 x7.x1.Qb1.n1 x7.x1.Qb1.n0 152
R4261 x7.x1.Qb1.n5 x7.x1.Qb1.n1 41.5091
R4262 x7.x1.Qb1.n5 x7.x1.Qb1.n4 18.1966
R4263 x7.x1.Qb1.n4 x7.x1.Qb1.n3 9.35675
R4264 x7.x1.Qb1.n3 x7.x1.Qb1 6.49269
R4265 x7.x1.Qb1.n1 x7.x1.Qb1 4.20621
R4266 x7.x1.Qb1.n3 x7.x1.Qb1 3.52967
R4267 x7.x1.Qb1 x7.x1.Qb1.n5 2.5605
R4268 x7.x2.x2.Q x7.x2.x2.Q.t0 246.839
R4269 x7.x2.x2.Q x7.x2.x2.Q.t1 148.597
R4270 a_14035_n2743.t0 a_14035_n2743.t1 60.0005
R4271 a_24530_n20346.t0 a_24530_n20346.t1 81.9478
R4272 a_18932_n14760.t0 a_18932_n14760.t1 83.5579
R4273 x7.x1.x3.Q x7.x1.x3.Q.t0 240.05
R4274 x7.x1.x3.Q x7.x1.x3.Q.t1 155.386
R4275 a_2130_n19184.t0 a_2130_n19184.t1 82.0028
R4276 a_24530_n19018.t0 a_24530_n19018.t1 81.9478
R4277 a_10620_n9002.t0 a_10620_n9002.t1 83.9243
R4278 a_14035_n2281.t0 a_14035_n2281.t1 60.9236
R4279 a_24220_n8836.t0 a_24220_n8836.t1 83.56
R4280 a_2130_n20180.t0 a_2130_n20180.t1 82.0028
R4281 a_2130_n22172.t0 a_2130_n22172.t1 82.0028
R4282 a_24530_n22006.t0 a_24530_n22006.t1 81.9492
R4283 a_2130_n21840.t0 a_2130_n21840.t1 82.0028
R4284 a_2132_n16586.t0 a_2132_n16586.t1 83.9223
R4285 a_18932_n16420.t0 a_18932_n16420.t1 83.5579
R4286 a_10620_n8670.t0 a_10620_n8670.t1 83.9243
R4287 a_22601_n15524.t0 a_22601_n15524.t1 120.212
R4288 a_20579_n2425.t0 a_20579_n2425.n0 1327.82
R4289 a_20579_n2425.n0 a_20579_n2425.t1 194.655
R4290 a_20579_n2425.n0 a_20579_n2425.t2 63.3219
R4291 a_21198_n2247.t0 a_21198_n2247.t1 126.644
R4292 a_17747_n2241.n1 a_17747_n2241.t4 530.01
R4293 a_17747_n2241.t0 a_17747_n2241.n5 421.021
R4294 a_17747_n2241.n0 a_17747_n2241.t2 337.142
R4295 a_17747_n2241.n3 a_17747_n2241.t1 280.223
R4296 a_17747_n2241.n4 a_17747_n2241.t3 263.173
R4297 a_17747_n2241.n4 a_17747_n2241.t6 227.826
R4298 a_17747_n2241.n0 a_17747_n2241.t5 199.762
R4299 a_17747_n2241.n2 a_17747_n2241.n1 170.81
R4300 a_17747_n2241.n2 a_17747_n2241.n0 167.321
R4301 a_17747_n2241.n5 a_17747_n2241.n4 152
R4302 a_17747_n2241.n1 a_17747_n2241.t7 141.923
R4303 a_17747_n2241.n3 a_17747_n2241.n2 10.8376
R4304 a_17747_n2241.n5 a_17747_n2241.n3 2.50485
R4305 a_2132_n14594.t0 a_2132_n14594.t1 82.3314
R4306 a_18932_n14428.t0 a_18932_n14428.t1 83.5579
R4307 a_16163_n2425.n0 a_16163_n2425.t1 1327.82
R4308 a_16163_n2425.n0 a_16163_n2425.t2 194.655
R4309 a_16163_n2425.t0 a_16163_n2425.n0 63.3219
R4310 a_18371_n2247.t0 a_18371_n2247.n0 1327.82
R4311 a_18371_n2247.n0 a_18371_n2247.t2 194.655
R4312 a_18371_n2247.n0 a_18371_n2247.t1 63.3219
R4313 a_24220_n8504.t0 a_24220_n8504.t1 83.56
R4314 x7.x2.x4.Q x7.x2.x4.Q.t0 246.839
R4315 x7.x2.x4.Q x7.x2.x4.Q.t1 148.597
R4316 a_18932_n16752.t0 a_18932_n16752.t1 83.5579
R4317 a_2130_n21508.t0 a_2130_n21508.t1 82.0028
R4318 a_24530_n21674.t0 a_24530_n21674.t1 81.9478
R4319 a_21390_n2791.t0 a_21390_n2791.t1 87.1434
R4320 a_2130_n18852.t0 a_2130_n18852.t1 82.0028
R4321 a_21390_n1881.t0 a_21390_n1881.t1 87.1434
R4322 a_8268_n12482.t1 a_8268_n12482.t0 193.599
R4323 a_21145_n2791.t1 a_21145_n2791.t0 94.7268
R4324 a_16782_n2247.t0 a_16782_n2247.t1 126.644
R4325 x7.x2.x3.Q x7.x2.x3.Q.t0 246.839
R4326 x7.x2.x3.Q x7.x2.x3.Q.t1 148.597
R4327 a_10620_n8006.t0 a_10620_n8006.t1 83.9243
R4328 a_2132_n16254.t0 a_2132_n16254.t1 83.9053
R4329 a_16729_n2791.t0 a_16729_n2791.t1 94.7268
R4330 a_2132_n17914.t0 a_2132_n17914.t1 83.9223
R4331 a_21198_n2425.t0 a_21198_n2425.t1 126.644
R4332 a_18932_n16088.t0 a_18932_n16088.t1 83.5579
R4333 a_18371_n2425.n0 a_18371_n2425.t1 1327.82
R4334 a_18371_n2425.n0 a_18371_n2425.t2 194.655
R4335 a_18371_n2425.t0 a_18371_n2425.n0 63.3219
R4336 a_18990_n2247.t0 a_18990_n2247.t1 126.644
R4337 a_2132_n14262.t0 a_2132_n14262.t1 83.9053
R4338 a_2132_n15922.t0 a_2132_n15922.t1 83.9223
C0 x7.x2.x2.CLK x7.stby_done_b 0.055466f
C1 vn xout 0.039662f
C2 avdd_ip dvss_ip 20.735699f
C3 dvdd_ip avss_ip 2.2865f
C4 dvss_ip vrb 1.20334f
C5 x7.x1.x2.Q x7.ena_done_b 0.012057f
C6 vg1 xout 0.637062f
C7 inv_in xin 0.302115f
C8 vg1 vg2 1.36272f
C9 standby_33 dvdd 0.092308f
C10 dvdd x7.x2.x4.Q 0.118417f
C11 xin xout 12.4168f
C12 x7.x1.x4.Q x7.ena_done_b 0.061065f
C13 x4.out_b standby_33 0.696369f
C14 x7.x1.Qb1 x7.ena_done_b 0.095485f
C15 dvdd_ip dvdd 14.0307f
C16 dvss_ip x7.stby_done_b 1.50194f
C17 ibias_ip dvss_ip 20.300303f
C18 avdd_ip avss_ip 0.856941p
C19 avss_ip vrb 6.48162f
C20 x7.x2.Qb2 dvdd 1.2179f
C21 vg2 xin 6.28706f
C22 standby_33 ibias 1.10533f
C23 avdd standby_33 9.00234f
C24 dvss_ip ena_ip 0.012218f
C25 avdd dvdd_ip 0.061641f
C26 inv_in xout 1.1656f
C27 vbp tail 10.143401f
C28 x7.x2.Qb1 x7.stby_done_b 0.111333f
C29 inv_in vg2 0.137694f
C30 dvdd x7.x2.x2.CLK 0.367738f
C31 dvss_ip avss_ip 23.869501f
C32 vbp dvdd_ip 26.197498f
C33 vg2 xout 0.938912f
C34 standby_33 avss 1.55853f
C35 inv_in inv_m1 0.243271f
C36 x7.x1.x3.Q x7.ena_done_b 0.012117f
C37 standby_ip dvdd_ip 3.44007f
C38 dvdd_ip avss 0.031496f
C39 avdd avdd_ip 9.33419f
C40 vn tail 0.670061f
C41 dvdd_ip dout 1.66314f
C42 dvdd x7.stby_done_b 5.41509f
C43 ibias_ip dvdd 0.020082f
C44 dvss_ip dvdd 20.2555f
C45 x7.clk_disable x7.x2.x2.CLK 0.012819f
C46 vn dvdd_ip 1.05192f
C47 x7.x2.x2.Q x7.stby_done_b 0.012057f
C48 standby ena_ip 0.035742f
C49 x7.x1.x2.CLK x7.x2.x2.CLK 0.011009f
C50 dvdd ena_ip 7.78413f
C51 x7.x1.Qb2 x7.ena_done_b 0.095442f
C52 vg1 dvdd_ip 0.707385f
C53 ibias_ip ibias 0.846688f
C54 dvss_ip ibias 0.012666f
C55 avdd_ip avss 0.574893f
C56 tail xin 1.6128f
C57 dvdd x7.x2.Qb1 1.15446f
C58 ibias ena_ip 0.171255f
C59 dvdd_ip xin 4.32555f
C60 avdd ena_ip 0.711014f
C61 x7.clk_disable x7.stby_done_b 0.724301f
C62 vbp ibias_ip 1.36181f
C63 x7.x2.x2.Q x7.x2.Qb1 0.040893f
C64 vbp dvss_ip 1.28877f
C65 inv_m1 inv_m2 0.947856f
C66 inv_in tail 0.604094f
C67 vg1 avdd_ip 1.99589f
C68 x7.x1.Qb2 x7.x1.x3.Q 0.040893f
C69 inv_in standby_33 0.08455f
C70 vg1 vrb 0.454276f
C71 avdd avss_ip 2.34938f
C72 tail xout 1.23159f
C73 inv_in dvdd_ip 10.408401f
C74 dvdd_ip x7.ena_done_b 0.022633f
C75 x7.x1.x2.CLK ena_ip 0.073063f
C76 dvdd standby 0.386478f
C77 standby_ip ena_ip 4.63202f
C78 avss ena_ip 1.87755f
C79 dvdd_ip xout 4.80514f
C80 dvss_ip dout 6.66227f
C81 avdd_ip xin 6.74409f
C82 vn dvss_ip 6.6789f
C83 dvdd x7.x2.x2.Q 0.11753f
C84 dvdd_ip vg2 0.10449f
C85 x7.x2.x3.Q x7.x2.Qb2 0.040893f
C86 x3.out avdd_ip 0.010186f
C87 dvdd ibias 0.083154f
C88 vg1 dvss_ip 6.37401f
C89 avss_ip avss 7.31391f
C90 avdd dvdd 0.106948f
C91 x4.out_b avdd 7.47205f
C92 inv_m1 dvdd_ip 2.8465f
C93 inv_in avdd_ip 0.669037f
C94 x7.x1.x2.Q ena_ip 0.035311f
C95 avdd_ip xout 7.21813f
C96 dvss_ip xin 1.63056f
C97 x7.clk_disable dvdd 0.383458f
C98 standby_ip standby 0.045013f
C99 avdd_ip vg2 0.488655f
C100 x7.x1.x2.CLK dvdd 0.406962f
C101 vrb vg2 4.64006f
C102 standby_ip dvdd 10.280701f
C103 vg1 avss_ip 20.7774f
C104 dvdd avss 0.230567f
C105 x4.out_b standby_ip 0.931668f
C106 x4.out_b avss 1.60462f
C107 x7.stby_done_b x7.ena_done_b 1.61077f
C108 inv_in ibias_ip 0.023743f
C109 x7.x1.Qb1 ena_ip 0.347396f
C110 dvss_ip x7.ena_done_b 1.48709f
C111 inv_in dvss_ip 14.9291f
C112 inv_m2 dvdd_ip 1.90217f
C113 dvdd dout 0.550876f
C114 x7.x2.Qb2 x7.x1.Qb2 0.0262f
C115 standby_ip ibias 0.288163f
C116 avss_ip xin 73.1079f
C117 dvss_ip xout 14.2041f
C118 avdd standby_ip 0.690112f
C119 avdd avss 0.110507p
C120 x7.ena_done_b ena_ip 0.702741f
C121 x7.x2.x3.Q x7.stby_done_b 0.012117f
C122 x7.x1.Qb1 x7.x2.Qb1 0.0262f
C123 dvss_ip vg2 3.9276f
C124 x3.out avss_ip 2.42141f
C125 x7.x1.x2.Q dvdd 0.116301f
C126 tail dvdd_ip 3.21426f
C127 inv_in avss_ip 1.9489f
C128 inv_m1 dvss_ip 3.10099f
C129 standby_33 dvdd_ip 3.26892f
C130 standby_ip avss 1.86774f
C131 avss_ip xout 26.396301f
C132 x7.x1.x3.Q ena_ip 0.035311f
C133 x7.x1.x4.Q dvdd 0.118427f
C134 x7.x1.Qb1 dvdd 1.22948f
C135 ena ena_ip 0.081602f
C136 avss_ip vg2 0.156017p
C137 inv_in dvdd 0.696511f
C138 dvdd x7.ena_done_b 6.16668f
C139 inv_m2 dvss_ip 1.69963f
C140 dvss_ip x7.x1.Qb2 0.069883f
C141 x3.out avdd 9.26841f
C142 dvdd_ip avdd_ip 3.59467f
C143 dvdd_ip vrb 0.182588f
C144 x7.x2.x3.Q dvdd 0.112734f
C145 inv_in avdd 0.025173f
C146 x7.x1.Qb2 ena_ip 0.347451f
C147 ena standby 0.095384f
C148 tail ibias_ip 0.011037f
C149 dvdd x7.x1.x3.Q 0.112744f
C150 tail dvss_ip 0.416372f
C151 vbp inv_in 0.265485f
C152 dvdd ena 0.377442f
C153 standby_33 ibias_ip 0.621612f
C154 x7.x2.x4.Q x7.stby_done_b 0.061065f
C155 x3.out avss 5.85073f
C156 standby_33 dvss_ip 3.27772f
C157 x7.x1.x2.CLK x7.ena_done_b 0.044383f
C158 ibias_ip dvdd_ip 1.46921f
C159 dvdd_ip x7.stby_done_b 0.02481f
C160 vn xin 3.09633f
C161 dvdd_ip dvss_ip 0.502455p
C162 standby_ip x7.ena_done_b 0.121215f
C163 x7.x2.Qb2 x7.stby_done_b 0.099468f
C164 inv_in avss 0.144174f
C165 x7.x2.Qb2 dvss_ip 0.07326f
C166 avdd ena 0.026781f
C167 vg1 xin 0.215332p
C168 x7.x1.Qb1 x7.x1.x2.Q 0.040893f
C169 dvdd x7.x1.Qb2 1.22125f
C170 vn inv_in 0.137437f
C171 xout dvss 4.260475f
C172 xin dvss 11.878201f
C173 dout dvss 6.13496f
C174 standby dvss 1.31628f
C175 ena dvss 1.29685f
C176 avss dvss 11.55251f
C177 ibias dvss 6.38685f
C178 dvdd dvss 0.140297p
C179 avdd dvss 95.102425f
C180 vg1 dvss -0.243245f
C181 vrb dvss 0.16284f
C182 vg2 dvss 4.397135f
C183 tail dvss 12.477897f
C184 inv_m2 dvss 0.562228f
C185 inv_m1 dvss 1.142152f
C186 inv_in dvss 6.596221f
C187 vn dvss 7.77323f
C188 vbp dvss 24.51475f
C189 x4.out_b dvss 1.061455f
C190 x3.out dvss 2.07027f
C191 x7.x2.x4.Q dvss 0.099773f
C192 x7.x2.x3.Q dvss 0.092032f
C193 x7.x2.Qb2 dvss 0.510929f
C194 x7.x2.x2.Q dvss 0.092454f
C195 x7.x2.Qb1 dvss 0.540099f
C196 x7.x2.x2.CLK dvss 0.389657f
C197 x7.clk_disable dvss 4.60726f
C198 x7.x1.x4.Q dvss 0.099773f
C199 x7.x1.x3.Q dvss 0.092032f
C200 x7.x1.x2.Q dvss 0.092454f
C201 x7.stby_done_b dvss 3.876771f
C202 ibias_ip dvss 13.1769f
C203 standby_33 dvss 13.62504f
C204 x7.x1.Qb2 dvss 0.510897f
C205 x7.x1.Qb1 dvss 0.528095f
C206 x7.x1.x2.CLK dvss 0.38222f
C207 x7.ena_done_b dvss 5.912164f
C208 standby_ip dvss 26.074802f
C209 ena_ip dvss 26.648424f
C210 avss_ip dvss 29.749199f
C211 dvss_ip dvss 41.9846f
C212 avdd_ip dvss 0.98484p
C213 dvdd_ip dvss 0.377434p
C214 a_8268_n12482.t1 dvss 0.033931f
C215 a_8268_n12482.t0 dvss 3.56607f
C216 a_22601_n15524.t1 dvss 1.2f
C217 a_22601_n15524.t0 dvss 1.2f
C218 dout.t0 dvss 0.040138f
C219 dout.t1 dvss 0.223213f
C220 dout.n0 dvss 3.29562f
C221 x4.out_b.n0 dvss 5.53652f
C222 x4.out_b.t3 dvss 1.30743f
C223 x4.out_b.t1 dvss 0.044437f
C224 x4.out_b.t2 dvss 0.044437f
C225 x4.out_b.n1 dvss 0.140668f
C226 x4.out_b.t0 dvss 0.055178f
C227 x7.clkout dvss 5.76435f
C228 dout_filt.t2 dvss 0.033084f
C229 dout_filt.n0 dvss 0.063466f
C230 dout_filt.t1 dvss 0.020119f
C231 dout_filt.n1 dvss 0.064349f
C232 x7.x5.Z dvss 0.084653f
C233 dout_filt.t0 dvss 0.028544f
C234 dout_filt.t3 dvss 0.296603f
C235 dout_filt.t4 dvss 0.738515f
C236 dout_filt.n2 dvss 6.50632f
C237 x3.out.n0 dvss 7.39524f
C238 x3.out.n1 dvss 0.893601f
C239 x3.out.n2 dvss 0.392503f
C240 x3.out.t6 dvss 0.479128f
C241 x3.out.n3 dvss 0.382459f
C242 x3.out.t8 dvss 0.458669f
C243 x3.out.n4 dvss 0.394877f
C244 x3.out.t7 dvss 0.479113f
C245 x3.out.t4 dvss 0.458669f
C246 x3.out.n5 dvss 0.382543f
C247 x3.out.t3 dvss 0.458669f
C248 x3.out.n6 dvss 0.161457f
C249 x3.out.n7 dvss 0.521199f
C250 x3.out.n8 dvss 1.69978f
C251 x3.out.t5 dvss 1.7568f
C252 x3.out.t0 dvss 0.059712f
C253 x3.out.t1 dvss 0.059712f
C254 x3.out.n9 dvss 0.188953f
C255 x3.out.t2 dvss 0.074144f
C256 vn.n0 dvss 0.636215f
C257 vn.n1 dvss 0.311146f
C258 vn.t7 dvss 0.039422f
C259 vn.t5 dvss 0.039422f
C260 vn.n2 dvss 0.106375f
C261 vn.t6 dvss 0.171883f
C262 vn.n3 dvss 0.444704f
C263 vn.t8 dvss 0.871134f
C264 vn.t9 dvss 1.02426f
C265 vn.n4 dvss 0.591267f
C266 vn.n5 dvss 0.320978f
C267 vn.t2 dvss 0.973785f
C268 vn.t1 dvss 0.039422f
C269 vn.t3 dvss 0.039422f
C270 vn.n6 dvss 0.078843f
C271 vn.t4 dvss 0.133384f
C272 vn.n7 dvss 0.489753f
C273 vn.n8 dvss 0.299827f
C274 vn.t0 dvss 0.871134f
C275 vn.n9 dvss 0.296493f
C276 vrb.t2 dvss 0.274519f
C277 vrb.t4 dvss 0.33602f
C278 vrb.n0 dvss 3.02505f
C279 vrb.t3 dvss 0.274548f
C280 vrb.t1 dvss 0.333171f
C281 vrb.n1 dvss 3.02989f
C282 vrb.t0 dvss 0.080693f
C283 vrb.n2 dvss 2.40037f
C284 vrb.n3 dvss 1.30448f
C285 vg2.n0 dvss 0.282949f
C286 vg2.n1 dvss 0.261019f
C287 vg2.t9 dvss 0.640509f
C288 vg2.n2 dvss 1.17147f
C289 vg2.n3 dvss 0.244906f
C290 vg2.n4 dvss 0.522037f
C291 vg2.t6 dvss 0.628646f
C292 vg2.n5 dvss 0.314177f
C293 vg2.n6 dvss 0.32051f
C294 vg2.n7 dvss 0.282949f
C295 vg2.n8 dvss 0.261019f
C296 vg2.t5 dvss 0.640544f
C297 vg2.n9 dvss 1.17258f
C298 vg2.n10 dvss 0.244906f
C299 vg2.n11 dvss 0.522037f
C300 vg2.t7 dvss 0.628646f
C301 vg2.n12 dvss 0.313029f
C302 vg2.n13 dvss 0.32051f
C303 vg2.n14 dvss 0.051368f
C304 vg2.t4 dvss 0.031316f
C305 vg2.t8 dvss 0.505469f
C306 vg2.t1 dvss 39.125f
C307 vg2.t0 dvss 39.3426f
C308 vg2.t3 dvss 39.3426f
C309 vg2.t2 dvss 39.11f
C310 vg2.n15 dvss 9.00528f
C311 vg2.n16 dvss 2.91513f
C312 xin.t21 dvss 0.023968f
C313 xin.t8 dvss 0.023338f
C314 xin.n0 dvss 0.172822f
C315 xin.n1 dvss 0.096776f
C316 xin.n2 dvss 0.096776f
C317 xin.n3 dvss 0.096776f
C318 xin.n4 dvss 0.096776f
C319 xin.n5 dvss 0.184148f
C320 xin.t18 dvss 0.1922f
C321 xin.t15 dvss 0.19211f
C322 xin.n6 dvss 0.184148f
C323 xin.n7 dvss 0.096776f
C324 xin.t13 dvss 0.19211f
C325 xin.n8 dvss 0.096776f
C326 xin.t19 dvss 0.19211f
C327 xin.n9 dvss 0.096776f
C328 xin.n10 dvss 0.096776f
C329 xin.t16 dvss 0.19211f
C330 xin.n11 dvss 0.096776f
C331 xin.t11 dvss 0.19211f
C332 xin.n12 dvss 0.096776f
C333 xin.n13 dvss 0.096776f
C334 xin.t10 dvss 0.19211f
C335 xin.n14 dvss 0.096776f
C336 xin.t17 dvss 0.19211f
C337 xin.n15 dvss 0.096776f
C338 xin.n16 dvss 0.096776f
C339 xin.t14 dvss 0.19211f
C340 xin.n17 dvss 0.096776f
C341 xin.t12 dvss 0.19211f
C342 xin.n18 dvss 0.096776f
C343 xin.n19 dvss 0.096776f
C344 xin.t9 dvss 0.19211f
C345 xin.n20 dvss 0.096776f
C346 xin.t6 dvss 0.19211f
C347 xin.n21 dvss 0.175223f
C348 xin.n22 dvss 0.784969f
C349 xin.n23 dvss 0.308623f
C350 xin.n24 dvss 0.374761f
C351 xin.t20 dvss 0.828066f
C352 xin.t7 dvss 0.796281f
C353 xin.n25 dvss 0.514f
C354 xin.n26 dvss 0.386948f
C355 xin.n27 dvss 3.79487f
C356 xin.n28 dvss 4.5191f
C357 xin.n29 dvss 3.61279f
C358 xin.t2 dvss 57.0239f
C359 xin.t4 dvss 44.1862f
C360 xin.t1 dvss 44.012f
C361 xin.t0 dvss 0.124226f
C362 xin.n30 dvss 4.7746f
C363 xin.n31 dvss 27.2736f
C364 xin.t5 dvss 31.1925f
C365 xin.n32 dvss 27.266699f
C366 xin.t3 dvss 31.1614f
C367 xin.n33 dvss 27.270199f
C368 xin.n34 dvss 3.77704f
C369 xin.n35 dvss 1.85671f
C370 xin.n36 dvss 0.500575f
C371 vg1.t3 dvss 0.056949f
C372 vg1.n0 dvss 0.44953f
C373 vg1.t8 dvss 46.057503f
C374 vg1.t9 dvss 46.8352f
C375 vg1.t4 dvss 23.996801f
C376 vg1.n1 dvss 23.9575f
C377 vg1.t7 dvss 23.996801f
C378 vg1.n2 dvss 23.4861f
C379 vg1.t6 dvss 23.996801f
C380 vg1.n3 dvss 12.9859f
C381 vg1.n4 dvss 15.228601f
C382 vg1.t0 dvss 0.01371f
C383 vg1.n5 dvss 3.04049f
C384 vg1.n6 dvss 1.50262f
C385 vg1.t1 dvss 0.271659f
C386 vg1.t5 dvss 0.353472f
C387 vg1.n7 dvss 0.229145f
C388 vg1.n8 dvss 0.08087f
C389 vg1.t2 dvss 0.049005f
C390 vg1.n9 dvss 0.281876f
C391 vg1.n10 dvss 0.146945f
C392 vg1.n11 dvss 0.153437f
C393 vg1.n12 dvss 0.372304f
C394 x3.out_b.t6 dvss 0.402581f
C395 x3.out_b.n0 dvss 0.790285f
C396 x3.out_b.n1 dvss 1.5584f
C397 x3.out_b.n2 dvss 6.60541f
C398 x3.out_b.t4 dvss 0.420289f
C399 x3.out_b.n3 dvss 0.339622f
C400 x3.out_b.t7 dvss 0.402581f
C401 x3.out_b.n4 dvss 0.342378f
C402 x3.out_b.t8 dvss 0.420331f
C403 x3.out_b.n5 dvss 0.338349f
C404 x3.out_b.t3 dvss 0.402581f
C405 x3.out_b.n6 dvss 0.345348f
C406 x3.out_b.n7 dvss 0.58218f
C407 x3.out_b.t5 dvss 1.5189f
C408 x3.out_b.t1 dvss 0.051624f
C409 x3.out_b.t2 dvss 0.051624f
C410 x3.out_b.n8 dvss 0.163419f
C411 x3.out_b.t0 dvss 0.064102f
C412 avdd.n0 dvss 0.492818f
C413 avdd.t6 dvss 0.034087f
C414 avdd.n1 dvss 1.6981f
C415 avdd.n2 dvss 0.060856f
C416 avdd.n3 dvss 0.056499f
C417 avdd.n4 dvss 0.266474f
C418 avdd.n5 dvss 0.585389f
C419 avdd.n6 dvss 1.03476f
C420 avdd.n7 dvss 1.03476f
C421 avdd.t4 dvss 0.894926f
C422 avdd.t9 dvss 0.702496f
C423 avdd.t18 dvss 0.894926f
C424 avdd.t15 dvss 0.702496f
C425 avdd.n8 dvss 0.46232f
C426 avdd.t12 dvss 7.53658f
C427 avdd.n9 dvss 7.5153f
C428 avdd.t11 dvss 9.12027f
C429 avdd.t14 dvss 7.25381f
C430 avdd.n10 dvss 7.71793f
C431 avdd.t13 dvss 9.163919f
C432 avdd.n11 dvss 3.68652f
C433 avdd.n12 dvss 0.768588f
C434 avdd.n13 dvss 0.579746f
C435 avdd.n14 dvss 0.560241f
C436 avdd.n15 dvss 0.353066f
C437 avdd.n16 dvss 0.487874f
C438 avdd.n17 dvss 3.7478f
C439 avdd.n18 dvss 0.731215f
C440 avdd.t16 dvss 0.036998f
C441 avdd.t19 dvss 0.036998f
C442 avdd.n19 dvss 0.090684f
C443 avdd.t10 dvss 0.036998f
C444 avdd.t8 dvss 0.036998f
C445 avdd.n20 dvss 0.090684f
C446 avdd.n21 dvss 1.93441f
C447 avdd.n22 dvss 0.967373f
C448 avdd.t5 dvss 0.135207f
C449 avdd.n23 dvss 0.34342f
C450 avdd.n24 dvss 5.68989f
C451 avdd.n25 dvss 1.05169f
C452 avdd.n26 dvss 1.1887f
C453 avdd.n27 dvss 1.1887f
C454 avdd.n28 dvss 4.46094f
C455 avdd.n29 dvss 1.35368f
C456 avdd.n30 dvss 0.090671f
C457 avdd.n31 dvss 0.071983f
C458 avdd.n32 dvss 0.548551f
C459 avdd.n33 dvss 1.56238f
C460 avdd.t1 dvss 0.034087f
C461 avdd.n34 dvss 1.46595f
C462 avdd.n35 dvss 0.107384f
C463 avdd.n36 dvss 0.107943f
C464 avdd.n37 dvss 0.158157f
C465 avdd.t0 dvss 2.51038f
C466 avdd.n38 dvss 0.071983f
C467 avdd.n39 dvss 0.10415f
C468 avdd.n40 dvss 0.107943f
C469 avdd.n41 dvss 0.559667f
C470 avdd.t17 dvss 0.034087f
C471 avdd.n42 dvss 0.023315f
C472 avdd.n43 dvss 0.687088f
C473 avdd.n44 dvss 1.48367f
C474 avdd.n45 dvss 1.13727f
C475 avdd.n46 dvss 0.744579f
C476 avdd.n47 dvss 2.46523f
C477 avdd.n48 dvss 3.43088f
C478 avdd.n49 dvss 1.15288f
C479 avdd.n50 dvss 0.362301f
C480 avdd.n51 dvss 0.321745f
C481 avdd.n52 dvss 0.106191f
C482 avdd.n53 dvss 1.67879f
C483 avdd.n54 dvss 0.106191f
C484 avdd.n55 dvss 0.158157f
C485 avdd.n56 dvss 0.090671f
C486 avdd.n57 dvss 0.062903f
C487 avdd.n58 dvss 0.106191f
C488 avdd.n59 dvss 1.67879f
C489 avdd.n60 dvss 0.106191f
C490 avdd.n61 dvss 0.060856f
C491 avdd.n62 dvss 0.116928f
C492 avdd.n63 dvss 0.719248f
C493 avdd.n64 dvss 1.37927f
C494 avdd.n65 dvss 1.47231f
C495 avdd.t3 dvss 0.034087f
C496 avdd.n66 dvss 1.45902f
C497 avdd.n67 dvss 0.366507f
C498 avdd.n68 dvss 0.107943f
C499 avdd.n69 dvss 0.158157f
C500 avdd.t2 dvss 2.51038f
C501 avdd.n70 dvss 0.10415f
C502 avdd.n71 dvss 0.107943f
C503 avdd.n72 dvss 0.107384f
C504 avdd.n73 dvss 0.062903f
C505 avdd.n74 dvss 0.106191f
C506 avdd.n75 dvss 1.67879f
C507 avdd.n76 dvss 0.106191f
C508 avdd.n77 dvss 0.158157f
C509 avdd.n78 dvss 0.106191f
C510 avdd.n79 dvss 1.67879f
C511 avdd.n80 dvss 0.106191f
C512 avdd.n81 dvss 0.319178f
C513 avdd.n82 dvss 0.73302f
C514 avdd.n83 dvss 1.95073f
C515 avdd.n84 dvss 4.13419f
C516 avdd.n85 dvss 0.707422f
C517 avdd.n86 dvss 0.479606f
C518 avdd.n87 dvss 1.32047f
C519 avdd.n88 dvss 1.35617f
C520 avdd.n89 dvss 0.536684f
C521 avdd.n90 dvss 1.19042f
C522 avdd.n91 dvss 4.48227f
C523 avdd.n92 dvss 4.46094f
C524 avdd.n93 dvss 4.48227f
C525 avdd.n94 dvss 1.19042f
C526 avdd.n95 dvss 0.66577f
C527 avdd.n96 dvss 3.27742f
C528 avdd.n97 dvss 0.20944f
C529 avdd.t7 dvss 0.702496f
C530 avdd.n98 dvss 0.20944f
C531 avdd.n99 dvss 0.731637f
C532 avdd.n100 dvss 0.757787f
C533 avdd.n101 dvss 0.146948f
C534 avdd.n102 dvss 0.057614f
C535 avdd.n103 dvss 0.303016f
C536 avss.n0 dvss 0.274689f
C537 avss.n1 dvss 0.256432f
C538 avss.t7 dvss 0.062902f
C539 avss.n2 dvss 0.199691f
C540 avss.n3 dvss 0.027139f
C541 avss.n4 dvss 0.10291f
C542 avss.n5 dvss 0.092262f
C543 avss.n6 dvss 0.092262f
C544 avss.t6 dvss 0.441575f
C545 avss.t4 dvss 0.441575f
C546 avss.n7 dvss 0.044347f
C547 avss.n8 dvss 0.078584f
C548 avss.t5 dvss 0.063155f
C549 avss.t21 dvss 0.063155f
C550 avss.n9 dvss 0.832446f
C551 avss.n10 dvss 0.117588f
C552 avss.t11 dvss 0.062902f
C553 avss.t23 dvss 0.062902f
C554 avss.n11 dvss 0.501337f
C555 avss.n12 dvss 0.044307f
C556 avss.n13 dvss 0.093826f
C557 avss.n14 dvss 0.093826f
C558 avss.n15 dvss 0.506602f
C559 avss.n16 dvss 0.092262f
C560 avss.n17 dvss 0.506602f
C561 avss.t20 dvss 0.441575f
C562 avss.n18 dvss 0.238935f
C563 avss.t22 dvss 0.441575f
C564 avss.n19 dvss 3.28532f
C565 avss.n20 dvss 7.3481f
C566 avss.t10 dvss 0.441575f
C567 avss.n21 dvss 0.093826f
C568 avss.n22 dvss 0.093826f
C569 avss.n23 dvss 0.078584f
C570 avss.n24 dvss 0.152326f
C571 avss.n25 dvss 0.092262f
C572 avss.n26 dvss 0.092262f
C573 avss.n27 dvss 0.238935f
C574 avss.t12 dvss 0.441575f
C575 avss.n28 dvss 0.092262f
C576 avss.n29 dvss 0.506602f
C577 avss.n30 dvss 0.506602f
C578 avss.t0 dvss 0.441575f
C579 avss.t2 dvss 0.441575f
C580 avss.n31 dvss 0.044347f
C581 avss.t13 dvss 0.063155f
C582 avss.t1 dvss 0.063155f
C583 avss.t3 dvss 0.062902f
C584 avss.t15 dvss 0.080794f
C585 avss.n32 dvss 0.370586f
C586 avss.n33 dvss 0.325025f
C587 avss.n34 dvss 0.132878f
C588 avss.n35 dvss 0.404741f
C589 avss.n36 dvss 2.98049f
C590 avss.t24 dvss 0.860518f
C591 avss.t18 dvss 0.732948f
C592 avss.n37 dvss 2.16357f
C593 avss.n38 dvss 1.84584f
C594 avss.t14 dvss 0.841962f
C595 avss.t16 dvss 0.732948f
C596 avss.n39 dvss 0.3741f
C597 avss.n40 dvss 0.133098f
C598 avss.t8 dvss 0.732948f
C599 avss.n41 dvss 0.133098f
C600 avss.n42 dvss 1.68799f
C601 avss.n43 dvss 0.462717f
C602 avss.t9 dvss 0.023705f
C603 avss.t17 dvss 0.023705f
C604 avss.n44 dvss 0.079436f
C605 avss.t25 dvss 0.023705f
C606 avss.t19 dvss 0.023705f
C607 avss.n45 dvss 0.086235f
C608 avss.n46 dvss 1.36147f
C609 avss.n47 dvss 1.03577f
C610 avss.t26 dvss 8.17429f
C611 avss.n48 dvss 7.701231f
C612 avss.t29 dvss 8.17429f
C613 avss.n49 dvss 8.01034f
C614 avss.t28 dvss 8.17429f
C615 avss.n50 dvss 7.90618f
C616 avss.n51 dvss 4.01706f
C617 avss.t27 dvss 8.17429f
C618 avss.n52 dvss 2.18128f
C619 avss.n53 dvss 4.97729f
C620 avss.n54 dvss 1.85282f
C621 avss.n55 dvss 1.94389f
C622 avss.n56 dvss 1.85115f
C623 avss.n57 dvss 0.09532f
C624 avss.n58 dvss 0.227287f
C625 avss.n59 dvss 0.265186f
C626 avss.n60 dvss 0.643717f
C627 avss.n61 dvss 0.274689f
C628 avss.n62 dvss 0.354568f
C629 avss.n63 dvss 0.078584f
C630 avss.n64 dvss 0.102951f
C631 avss.n65 dvss 0.027139f
C632 avss.n66 dvss 0.036993f
C633 avss.n67 dvss 0.093826f
C634 avss.n68 dvss 0.238935f
C635 avss.n69 dvss 0.093826f
C636 avss.n70 dvss 0.036957f
C637 avss.n71 dvss 0.10291f
C638 avss.n72 dvss 0.044307f
C639 avss.n73 dvss 0.117505f
C640 avss.n74 dvss 0.092262f
C641 avss.n75 dvss 0.79544f
C642 avss.n76 dvss 1.9882f
C643 avss.n77 dvss 0.79544f
C644 avss.n78 dvss 0.092262f
C645 avss.n79 dvss 0.117505f
C646 avss.n80 dvss 0.117588f
C647 avss.n81 dvss 0.455799f
C648 avss.n82 dvss 1.20688f
C649 avss.n83 dvss 0.606761f
C650 avss.n84 dvss 0.354568f
C651 avss.n85 dvss 0.078584f
C652 avss.n86 dvss 0.102951f
C653 avss.n87 dvss 0.036993f
C654 avss.n88 dvss 0.093826f
C655 avss.n89 dvss 0.238935f
C656 avss.n90 dvss 0.093826f
C657 avss.n91 dvss 0.036957f
C658 avss.n92 dvss 0.152326f
C659 avss.n93 dvss 0.088692f
C660 avss.n94 dvss 0.162188f
C661 avss.n95 dvss 0.241706f
C662 standby_ip.n0 dvss 0.437228f
C663 standby_ip.n1 dvss 2.91743f
C664 standby_ip.n2 dvss 0.095599f
C665 standby_ip.t0 dvss 0.020325f
C666 standby_ip.t1 dvss 0.029229f
C667 standby_ip.t3 dvss 0.018853f
C668 standby_ip.t14 dvss 0.011782f
C669 standby_ip.n4 dvss 0.033754f
C670 standby_ip.n5 dvss 0.059774f
C671 standby_ip.t10 dvss 0.927569f
C672 standby_ip.n6 dvss 0.640216f
C673 standby_ip.n7 dvss 0.111584f
C674 standby_ip.n8 dvss 0.207294f
C675 standby_ip.t15 dvss 0.300607f
C676 standby_ip.t9 dvss 0.285452f
C677 standby_ip.n9 dvss 0.207294f
C678 standby_ip.n10 dvss 0.111584f
C679 standby_ip.t8 dvss 0.285452f
C680 standby_ip.n11 dvss 0.111584f
C681 standby_ip.t12 dvss 0.285452f
C682 standby_ip.n12 dvss 0.111584f
C683 standby_ip.n13 dvss 0.101714f
C684 standby_ip.t11 dvss 0.285452f
C685 standby_ip.n14 dvss 0.101714f
C686 standby_ip.n15 dvss 0.111584f
C687 standby_ip.n16 dvss 0.212597f
C688 standby_ip.t4 dvss 0.301362f
C689 standby_ip.t6 dvss 0.285452f
C690 standby_ip.n17 dvss 0.211536f
C691 standby_ip.n18 dvss 0.111584f
C692 standby_ip.t17 dvss 0.285452f
C693 standby_ip.n19 dvss 0.111584f
C694 standby_ip.t18 dvss 0.285452f
C695 standby_ip.n20 dvss 0.111584f
C696 standby_ip.n21 dvss 0.098853f
C697 standby_ip.t5 dvss 0.285452f
C698 standby_ip.n22 dvss 0.098853f
C699 standby_ip.t2 dvss 0.261318f
C700 standby_ip.n23 dvss 0.226201f
C701 standby_ip.t13 dvss 0.236298f
C702 standby_ip.t7 dvss 0.236114f
C703 standby_ip.n24 dvss 0.198459f
C704 standby_ip.n25 dvss 0.912751f
C705 standby_ip.t16 dvss 0.270102f
C706 standby_ip.n26 dvss 0.12259f
C707 xin_buf.t3 dvss 0.205358p
C708 xin_buf.t0 dvss 0.22283f
C709 xin_buf.t1 dvss 0.075836f
C710 xin_buf.n0 dvss 0.129036f
C711 xin_buf.t2 dvss 0.263405f
C712 xin_buf.t4 dvss 0.089459f
C713 xin_buf.n1 dvss 0.161326f
C714 x7.x1.x1.A dvss 0.017818f
C715 x7.x1.clkin dvss 0.290534f
C716 x7.x2.x1.A dvss 0.017818f
C717 x7.x2.clkin dvss 0.174689f
C718 x7.x5.A dvss 0.084584f
C719 dout_ip.n0 dvss 3.72627f
C720 x7.clkin dvss 5.05976f
C721 dout_ip.t9 dvss 0.01616f
C722 dout_ip.n1 dvss 0.038785f
C723 dout_ip.t6 dvss 0.012534f
C724 dout_ip.n2 dvss 0.033243f
C725 dout_ip.n3 dvss 0.027616f
C726 dout_ip.n4 dvss 0.027616f
C727 dout_ip.t5 dvss 0.012534f
C728 dout_ip.n5 dvss 0.033243f
C729 dout_ip.n6 dvss 0.35872f
C730 dout_ip.n7 dvss 0.352547f
C731 dout_ip.t2 dvss 0.022644f
C732 dout_ip.t3 dvss 0.022607f
C733 dout_ip.t1 dvss 0.021945f
C734 dout_ip.t0 dvss 0.021852f
C735 inv_m1.t0 dvss 0.045634f
C736 inv_m1.n0 dvss 1.05525f
C737 inv_m1.n1 dvss 0.129812f
C738 inv_m1.t5 dvss 0.363826f
C739 inv_m1.t2 dvss 0.363827f
C740 inv_m1.n2 dvss 0.117923f
C741 inv_m1.t4 dvss 0.341649f
C742 inv_m1.t3 dvss 0.34165f
C743 inv_m1.n3 dvss 2.65565f
C744 inv_m1.t1 dvss 0.046767f
C745 inv_in.t3 dvss 0.657711f
C746 inv_in.t11 dvss 5.68012f
C747 inv_in.n0 dvss 5.17707f
C748 inv_in.t5 dvss 5.52894f
C749 inv_in.n1 dvss 2.62426f
C750 inv_in.t6 dvss 5.52894f
C751 inv_in.n2 dvss 2.66147f
C752 inv_in.n3 dvss 2.79669f
C753 inv_in.t14 dvss 5.52894f
C754 inv_in.n4 dvss 5.29306f
C755 inv_in.t12 dvss 5.55261f
C756 inv_in.n5 dvss 5.28615f
C757 inv_in.t13 dvss 5.52894f
C758 inv_in.n6 dvss 2.66147f
C759 inv_in.t9 dvss 5.5836f
C760 inv_in.n7 dvss 5.39875f
C761 inv_in.t10 dvss 5.5836f
C762 inv_in.t2 dvss 5.5836f
C763 inv_in.n8 dvss 5.26653f
C764 inv_in.n9 dvss 5.40864f
C765 inv_in.t4 dvss 5.52894f
C766 inv_in.n10 dvss 2.66147f
C767 inv_in.n11 dvss 2.90209f
C768 inv_in.n12 dvss 2.75998f
C769 inv_in.t8 dvss 5.52894f
C770 inv_in.n13 dvss 2.62426f
C771 inv_in.n14 dvss 2.76492f
C772 inv_in.n15 dvss 2.76492f
C773 inv_in.n16 dvss 2.76201f
C774 inv_in.t7 dvss 5.52894f
C775 inv_in.n17 dvss 5.4592f
C776 inv_in.n18 dvss 0.82306f
C777 inv_in.t0 dvss 0.104143f
C778 inv_in.t1 dvss 0.647866f
C779 inv_in.n19 dvss 2.16816f
C780 xout.t26 dvss 0.047347f
C781 xout.t24 dvss 0.048657f
C782 xout.t22 dvss 0.243993f
C783 xout.t20 dvss 0.243993f
C784 xout.n0 dvss 2.4243f
C785 xout.t21 dvss 0.243993f
C786 xout.t19 dvss 0.243993f
C787 xout.n1 dvss 1.60432f
C788 xout.n2 dvss 6.32987f
C789 xout.t18 dvss 0.256529f
C790 xout.t11 dvss 0.243993f
C791 xout.n3 dvss 1.22843f
C792 xout.t16 dvss 0.256529f
C793 xout.t12 dvss 0.243993f
C794 xout.n4 dvss 1.23308f
C795 xout.n5 dvss 2.18555f
C796 xout.n6 dvss 8.527769f
C797 xout.n7 dvss 3.77761f
C798 xout.t13 dvss 0.243993f
C799 xout.t14 dvss 0.243993f
C800 xout.n8 dvss 1.27442f
C801 xout.n9 dvss 1.83376f
C802 xout.t15 dvss 0.243993f
C803 xout.t17 dvss 0.243993f
C804 xout.n10 dvss 1.43377f
C805 xout.n11 dvss 1.68066f
C806 xout.n12 dvss 1.24537f
C807 xout.t1 dvss 0.066767f
C808 xout.t7 dvss 0.066767f
C809 xout.n13 dvss 0.227228f
C810 xout.t0 dvss 0.066767f
C811 xout.t4 dvss 0.066767f
C812 xout.n14 dvss 0.217681f
C813 xout.t8 dvss 0.066767f
C814 xout.t2 dvss 0.066767f
C815 xout.n15 dvss 0.229174f
C816 xout.n16 dvss 4.49086f
C817 xout.t6 dvss 0.066767f
C818 xout.t10 dvss 0.066767f
C819 xout.n17 dvss 0.217681f
C820 xout.t9 dvss 0.066767f
C821 xout.t5 dvss 0.066767f
C822 xout.n18 dvss 0.149204f
C823 xout.n19 dvss 2.97025f
C824 xout.n20 dvss 3.47714f
C825 xout.n21 dvss 4.15788f
C826 xout.t3 dvss 0.091048f
C827 xout.n22 dvss 4.02374f
C828 xout.n23 dvss 0.626416f
C829 xout.n24 dvss 0.760656f
C830 xout.t25 dvss 1.61622f
C831 xout.t23 dvss 1.68073f
C832 xout.n25 dvss 1.04327f
C833 xout.n26 dvss 0.785936f
C834 xout.n27 dvss 8.087669f
C835 xout.n28 dvss 9.65943f
C836 xout.n29 dvss 1.9924f
C837 avdd_ip.t1 dvss 0.074663f
C838 avdd_ip.t4 dvss 0.074663f
C839 avdd_ip.n0 dvss 0.183001f
C840 avdd_ip.t0 dvss 0.074663f
C841 avdd_ip.t2 dvss 0.074663f
C842 avdd_ip.n1 dvss 0.193101f
C843 avdd_ip.t6 dvss 0.312571f
C844 avdd_ip.n2 dvss 25.687199f
C845 avdd_ip.t33 dvss 0.201546p
C846 avdd_ip.n3 dvss 42.3367f
C847 avdd_ip.n4 dvss 31.209301f
C848 avdd_ip.t30 dvss 12.6155f
C849 avdd_ip.n5 dvss 8.054391f
C850 avdd_ip.t31 dvss 12.6155f
C851 avdd_ip.n6 dvss 7.765079f
C852 avdd_ip.n7 dvss 10.2323f
C853 avdd_ip.t29 dvss 12.6155f
C854 avdd_ip.n8 dvss 11.3223f
C855 avdd_ip.t32 dvss 12.6155f
C856 avdd_ip.n9 dvss 11.2988f
C857 avdd_ip.n10 dvss 11.0453f
C858 avdd_ip.n11 dvss 25.8585f
C859 avdd_ip.n12 dvss 11.8125f
C860 avdd_ip.n13 dvss 15.647901f
C861 avdd_ip.t21 dvss 0.272851f
C862 avdd_ip.n14 dvss 0.353227f
C863 avdd_ip.t24 dvss 0.272851f
C864 avdd_ip.n15 dvss 1.24555f
C865 avdd_ip.t25 dvss 0.272851f
C866 avdd_ip.n16 dvss 1.36471f
C867 avdd_ip.t23 dvss 0.284354f
C868 avdd_ip.n17 dvss 1.00481f
C869 avdd_ip.n18 dvss 1.60279f
C870 avdd_ip.n19 dvss 0.908877f
C871 avdd_ip.n20 dvss 0.312041f
C872 avdd_ip.t26 dvss 0.272851f
C873 avdd_ip.n21 dvss 0.511759f
C874 avdd_ip.n22 dvss 1.0293f
C875 avdd_ip.n23 dvss 1.19091f
C876 avdd_ip.t20 dvss 0.272851f
C877 avdd_ip.n24 dvss 1.06873f
C878 avdd_ip.n25 dvss 4.33929f
C879 avdd_ip.n26 dvss 15.187299f
C880 avdd_ip.n27 dvss 15.187299f
C881 avdd_ip.t7 dvss 19.331099f
C882 avdd_ip.n28 dvss 1.61496f
C883 avdd_ip.t12 dvss 0.272851f
C884 avdd_ip.n29 dvss 5.41016f
C885 avdd_ip.t17 dvss 0.272851f
C886 avdd_ip.t18 dvss 0.272851f
C887 avdd_ip.n30 dvss 2.76186f
C888 avdd_ip.t14 dvss 0.272851f
C889 avdd_ip.t16 dvss 0.272851f
C890 avdd_ip.n31 dvss 1.60468f
C891 avdd_ip.n32 dvss 2.4602f
C892 avdd_ip.n33 dvss 6.7614f
C893 avdd_ip.n34 dvss 0.081048f
C894 avdd_ip.n35 dvss 0.056209f
C895 avdd_ip.n36 dvss 0.056638f
C896 avdd_ip.n37 dvss 0.056638f
C897 avdd_ip.n38 dvss 0.065474f
C898 avdd_ip.n39 dvss 0.058077f
C899 avdd_ip.n40 dvss 0.275331f
C900 avdd_ip.t3 dvss 0.366056f
C901 avdd_ip.n42 dvss -24.5529f
C902 avdd_ip.n43 dvss 24.8309f
C903 avdd_ip.n44 dvss 0.057159f
C904 avdd_ip.n45 dvss 0.06457f
C905 avdd_ip.n46 dvss 0.060147f
C906 avdd_ip.n47 dvss 2.63147f
C907 avdd_ip.n48 dvss 0.07741f
C908 avdd_ip.n49 dvss 0.056204f
C909 avdd_ip.n50 dvss 0.056638f
C910 avdd_ip.t5 dvss 0.425863f
C911 avdd_ip.n52 dvss 0.066326f
C912 avdd_ip.n53 dvss 0.05862f
C913 avdd_ip.n54 dvss 0.275331f
C914 avdd_ip.n55 dvss 0.056638f
C915 avdd_ip.n57 dvss 0.275331f
C916 avdd_ip.n58 dvss 0.06457f
C917 avdd_ip.n59 dvss 0.060147f
C918 avdd_ip.n60 dvss 2.34174f
C919 avdd_ip.n61 dvss 3.08369f
C920 avdd_ip.n62 dvss 7.458549f
C921 avdd_ip.t8 dvss 0.272851f
C922 avdd_ip.t9 dvss 0.272851f
C923 avdd_ip.t10 dvss 0.272851f
C924 avdd_ip.n63 dvss 2.28083f
C925 avdd_ip.t22 dvss 0.272851f
C926 avdd_ip.t28 dvss 0.272851f
C927 avdd_ip.n64 dvss 2.68748f
C928 avdd_ip.t19 dvss 0.272851f
C929 avdd_ip.t27 dvss 0.272851f
C930 avdd_ip.n65 dvss 1.60335f
C931 avdd_ip.n66 dvss 2.5326f
C932 avdd_ip.n67 dvss 6.54556f
C933 avdd_ip.n68 dvss 5.37955f
C934 avdd_ip.n69 dvss 12.5401f
C935 avdd_ip.n70 dvss 7.683919f
C936 avdd_ip.n71 dvss 8.52327f
C937 avdd_ip.n72 dvss 8.52327f
C938 avdd_ip.n73 dvss 32.6198f
C939 avdd_ip.n74 dvss 7.0648f
C940 avdd_ip.n75 dvss 2.67542f
C941 avdd_ip.n76 dvss 5.79729f
C942 avdd_ip.n77 dvss 37.3139f
C943 avdd_ip.n78 dvss 13.6449f
C944 avdd_ip.n79 dvss 32.799896f
C945 avdd_ip.n80 dvss 32.6198f
C946 avdd_ip.n81 dvss 32.799896f
C947 avdd_ip.n82 dvss 8.53496f
C948 avdd_ip.n83 dvss 8.47481f
C949 avdd_ip.n84 dvss 3.99638f
C950 avdd_ip.n85 dvss 32.939102f
C951 avdd_ip.n86 dvss 7.89575f
C952 avdd_ip.n87 dvss 2.20458f
C953 avdd_ip.n88 dvss 5.76955f
C954 avdd_ip.t13 dvss 0.272851f
C955 avdd_ip.t15 dvss 0.272851f
C956 avdd_ip.n89 dvss 2.2737f
C957 avdd_ip.n90 dvss 0.777352f
C958 avdd_ip.n91 dvss 1.40119f
C959 avdd_ip.t11 dvss 19.331099f
C960 avdd_ip.n92 dvss 16.5454f
C961 avdd_ip.n93 dvss 1.40119f
C962 avdd_ip.n94 dvss 2.89538f
C963 avdd_ip.n95 dvss 1.66736f
C964 avdd_ip.n96 dvss 7.11433f
C965 avdd_ip.n97 dvss 23.7224f
C966 ibias_ip.n0 dvss 4.75326f
C967 ibias_ip.n1 dvss 0.974101f
C968 ibias_ip.t13 dvss 0.653909f
C969 ibias_ip.t2 dvss 0.646782f
C970 ibias_ip.t3 dvss 0.082653f
C971 ibias_ip.t7 dvss 0.081898f
C972 ibias_ip.t6 dvss 0.644915f
C973 ibias_ip.t1 dvss 0.077591f
C974 ibias_ip.t0 dvss 0.650434f
C975 ibias_ip.t4 dvss 0.647233f
C976 ibias_ip.t11 dvss 0.653916f
C977 ibias_ip.t5 dvss 0.082116f
C978 ibias_ip.t9 dvss 0.082367f
C979 ibias_ip.t8 dvss 0.645067f
C980 ibias_ip.t12 dvss 0.646314f
C981 ibias_ip.t10 dvss 0.184945f
C982 standby_33.n0 dvss 7.3102f
C983 standby_33.t3 dvss 0.80334f
C984 standby_33.t4 dvss 1.62318f
C985 standby_33.t2 dvss 0.05517f
C986 standby_33.t1 dvss 0.05517f
C987 standby_33.n1 dvss 0.174581f
C988 standby_33.t0 dvss 0.068505f
C989 x7.ena_done_b.t1 dvss 0.054284f
C990 x7.ena_done_b.t0 dvss 0.068732f
C991 x7.ena_done_b.t3 dvss 0.033951f
C992 x7.ena_done_b.t2 dvss 0.02132f
C993 x7.ena_done_b.n0 dvss 0.045927f
C994 x7.ena_done_b.n1 dvss 0.058447f
C995 x7.ena_done_b.t4 dvss 0.018591f
C996 x7.ena_done_b.n2 dvss 0.053311f
C997 x7.ena_done_b.t7 dvss 0.018802f
C998 x7.ena_done_b.n3 dvss 0.05789f
C999 x7.ena_done_b.n4 dvss 0.011573f
C1000 x7.ena_done_b.n5 dvss 0.060019f
C1001 x7.ena_done_b.t6 dvss 0.025304f
C1002 x7.ena_done_b.t5 dvss 0.027855f
C1003 x7.ena_done_b.n6 dvss 0.079658f
C1004 x7.ena_done_b.n7 dvss 1.96309f
C1005 x7.ena_done_b.n8 dvss 0.077694f
C1006 a_9120_n9346.t1 dvss 0.036089f
C1007 a_9120_n9346.t0 dvss 1.47746f
C1008 a_9120_n9346.n0 dvss 3.32132f
C1009 a_9120_n9346.t2 dvss 1.67898f
C1010 a_9120_n9346.t3 dvss 0.027167f
C1011 a_9120_n9346.n1 dvss 2.97825f
C1012 a_9120_n9346.n2 dvss 1.80939f
C1013 a_9120_n9346.t4 dvss 0.071336f
C1014 x7.x2.x4.RESET_B dvss 1.471743f
C1015 x7.x3.A1 dvss 0.02912f
C1016 standby_b.n0 dvss 0.153287f
C1017 x4.in_b dvss 2.69011f
C1018 x7.x2.x2.RESET_B dvss 0.028793f
C1019 x7.x2.x3.RESET_B dvss 0.028793f
C1020 standby_b.n1 dvss 3.12348f
C1021 x7.stby_b dvss 1.34845f
C1022 standby_b.t12 dvss 0.182513f
C1023 standby_b.t4 dvss 0.182371f
C1024 standby_b.n2 dvss 0.084915f
C1025 standby_b.n3 dvss 0.157601f
C1026 standby_b.t19 dvss 0.228815f
C1027 standby_b.t17 dvss 0.217171f
C1028 standby_b.n4 dvss 0.157601f
C1029 standby_b.n5 dvss 0.084915f
C1030 standby_b.t7 dvss 0.217171f
C1031 standby_b.n6 dvss 0.084915f
C1032 standby_b.t23 dvss 0.217171f
C1033 standby_b.n7 dvss 0.084915f
C1034 standby_b.n8 dvss 0.077844f
C1035 standby_b.t21 dvss 0.217171f
C1036 standby_b.n9 dvss 0.077734f
C1037 standby_b.n10 dvss 0.084915f
C1038 standby_b.n11 dvss 0.162102f
C1039 standby_b.t6 dvss 0.229503f
C1040 standby_b.t16 dvss 0.217171f
C1041 standby_b.n12 dvss 0.161693f
C1042 standby_b.n13 dvss 0.084915f
C1043 standby_b.t18 dvss 0.217171f
C1044 standby_b.n14 dvss 0.084915f
C1045 standby_b.t0 dvss 0.217171f
C1046 standby_b.n15 dvss 0.084915f
C1047 standby_b.n16 dvss 0.074529f
C1048 standby_b.t3 dvss 0.217171f
C1049 standby_b.n17 dvss 0.07464f
C1050 standby_b.t14 dvss 0.014102f
C1051 standby_b.n18 dvss 0.025012f
C1052 standby_b.t25 dvss 0.014102f
C1053 standby_b.n20 dvss 0.025012f
C1054 standby_b.t11 dvss 0.014102f
C1055 standby_b.n22 dvss 0.025012f
C1056 standby_b.t2 dvss 0.012275f
C1057 standby_b.n24 dvss 0.023944f
C1058 standby_b.t15 dvss 0.012275f
C1059 standby_b.n25 dvss 0.023944f
C1060 standby_b.t13 dvss 0.012275f
C1061 standby_b.n26 dvss 0.023944f
C1062 standby_b.t24 dvss 0.014675f
C1063 standby_b.n27 dvss 0.022499f
C1064 tail.n0 dvss 0.76343f
C1065 tail.n1 dvss 2.82244f
C1066 tail.n2 dvss 0.753923f
C1067 tail.t11 dvss 0.054705f
C1068 tail.t10 dvss 0.054705f
C1069 tail.n3 dvss 0.119757f
C1070 tail.t0 dvss 0.102772f
C1071 tail.t5 dvss 0.102893f
C1072 tail.t7 dvss 0.102832f
C1073 tail.t2 dvss 0.102832f
C1074 tail.t4 dvss 0.103102f
C1075 tail.t9 dvss 0.102562f
C1076 tail.t3 dvss 0.103102f
C1077 tail.t8 dvss 0.102562f
C1078 tail.t6 dvss 0.102998f
C1079 tail.t1 dvss 0.102668f
C1080 dvdd_ip.n0 dvss 1.69476f
C1081 dvdd_ip.n1 dvss 9.839379f
C1082 dvdd_ip.n2 dvss 1.74378f
C1083 dvdd_ip.n3 dvss 0.433764f
C1084 dvdd_ip.n4 dvss 6.83399f
C1085 dvdd_ip.n5 dvss 0.511649f
C1086 dvdd_ip.n6 dvss 16.4905f
C1087 dvdd_ip.n7 dvss 5.38562f
C1088 dvdd_ip.n8 dvss 0.857057f
C1089 dvdd_ip.n9 dvss 0.547208f
C1090 dvdd_ip.n10 dvss 0.059815f
C1091 dvdd_ip.t56 dvss 0.407697p
C1092 dvdd_ip.n11 dvss 0.923193f
C1093 dvdd_ip.n12 dvss 0.626219f
C1094 dvdd_ip.n13 dvss 2.12711f
C1095 dvdd_ip.n14 dvss 1.11074f
C1096 dvdd_ip.n15 dvss 6.764f
C1097 dvdd_ip.n16 dvss 0.540653f
C1098 dvdd_ip.n17 dvss 1.29089f
C1099 dvdd_ip.n18 dvss 0.411041f
C1100 dvdd_ip.n19 dvss 0.257042f
C1101 dvdd_ip.n20 dvss 12.777401f
C1102 dvdd_ip.n21 dvss 2.28119f
C1103 dvdd_ip.n22 dvss 0.852694f
C1104 dvdd_ip.n23 dvss 0.753119f
C1105 dvdd_ip.n24 dvss 1.71693f
C1106 dvdd_ip.n25 dvss 0.719725f
C1107 dvdd_ip.n26 dvss 0.855677f
C1108 dvdd_ip.t24 dvss 0.08138f
C1109 dvdd_ip.t25 dvss 0.051814f
C1110 dvdd_ip.n27 dvss 0.496394f
C1111 dvdd_ip.t29 dvss 0.053882f
C1112 dvdd_ip.t33 dvss 0.051814f
C1113 dvdd_ip.t9 dvss 0.051814f
C1114 dvdd_ip.t27 dvss 0.054424f
C1115 dvdd_ip.t11 dvss 0.051814f
C1116 dvdd_ip.n28 dvss 0.366042f
C1117 dvdd_ip.t12 dvss 0.051814f
C1118 dvdd_ip.n29 dvss 0.278999f
C1119 dvdd_ip.n30 dvss 1.14823f
C1120 dvdd_ip.t18 dvss 0.054424f
C1121 dvdd_ip.t30 dvss 0.051814f
C1122 dvdd_ip.n31 dvss 0.366042f
C1123 dvdd_ip.t31 dvss 0.051814f
C1124 dvdd_ip.n32 dvss 0.278999f
C1125 dvdd_ip.n33 dvss 0.889286f
C1126 dvdd_ip.n34 dvss 0.249013f
C1127 dvdd_ip.t28 dvss 0.054363f
C1128 dvdd_ip.t22 dvss 0.051814f
C1129 dvdd_ip.n35 dvss 0.364127f
C1130 dvdd_ip.t21 dvss 0.051814f
C1131 dvdd_ip.n36 dvss 0.278999f
C1132 dvdd_ip.t20 dvss 0.054424f
C1133 dvdd_ip.t7 dvss 0.051814f
C1134 dvdd_ip.n37 dvss 0.366042f
C1135 dvdd_ip.t6 dvss 0.051814f
C1136 dvdd_ip.n38 dvss 0.278999f
C1137 dvdd_ip.n39 dvss 0.04435f
C1138 dvdd_ip.n40 dvss 0.332493f
C1139 dvdd_ip.n41 dvss 0.673943f
C1140 dvdd_ip.n42 dvss 0.776442f
C1141 dvdd_ip.n43 dvss 0.776442f
C1142 dvdd_ip.n44 dvss 0.45776f
C1143 dvdd_ip.n45 dvss 0.033319f
C1144 dvdd_ip.t37 dvss 0.01337f
C1145 dvdd_ip.n46 dvss 0.077263f
C1146 dvdd_ip.n49 dvss 0.505719f
C1147 dvdd_ip.n50 dvss 0.540653f
C1148 dvdd_ip.n51 dvss 0.975669f
C1149 dvdd_ip.n52 dvss 2.06088f
C1150 dvdd_ip.n53 dvss 2.06088f
C1151 dvdd_ip.n54 dvss 7.83078f
C1152 dvdd_ip.n55 dvss 0.821534f
C1153 dvdd_ip.n56 dvss 0.088522f
C1154 dvdd_ip.n57 dvss 0.835542f
C1155 dvdd_ip.n58 dvss 0.835542f
C1156 dvdd_ip.n59 dvss 0.638491f
C1157 dvdd_ip.n60 dvss 0.105906f
C1158 dvdd_ip.n61 dvss 0.098224f
C1159 dvdd_ip.n62 dvss 0.098224f
C1160 dvdd_ip.t45 dvss 1.169f
C1161 dvdd_ip.n65 dvss 0.098224f
C1162 dvdd_ip.n66 dvss 0.16276f
C1163 dvdd_ip.t46 dvss 0.01337f
C1164 dvdd_ip.t44 dvss 0.028653f
C1165 dvdd_ip.t51 dvss 0.028653f
C1166 dvdd_ip.n68 dvss 0.068717f
C1167 dvdd_ip.t55 dvss 0.028653f
C1168 dvdd_ip.t48 dvss 0.028653f
C1169 dvdd_ip.n69 dvss 0.068738f
C1170 dvdd_ip.t34 dvss 0.028653f
C1171 dvdd_ip.t47 dvss 0.028653f
C1172 dvdd_ip.n70 dvss 0.068717f
C1173 dvdd_ip.t43 dvss 0.028653f
C1174 dvdd_ip.t40 dvss 0.028653f
C1175 dvdd_ip.n71 dvss 0.068717f
C1176 dvdd_ip.t50 dvss 0.028653f
C1177 dvdd_ip.t39 dvss 0.028653f
C1178 dvdd_ip.n72 dvss 0.068738f
C1179 dvdd_ip.n73 dvss 1.79527f
C1180 dvdd_ip.n74 dvss 2.06716f
C1181 dvdd_ip.n75 dvss 7.9286f
C1182 dvdd_ip.n76 dvss 7.83078f
C1183 dvdd_ip.n77 dvss 7.9286f
C1184 dvdd_ip.n78 dvss 2.06716f
C1185 dvdd_ip.n79 dvss 1.53964f
C1186 dvdd_ip.n80 dvss 0.568083f
C1187 dvdd_ip.n81 dvss 0.067329f
C1188 dvdd_ip.t2 dvss 0.86612f
C1189 dvdd_ip.n84 dvss 0.067329f
C1190 dvdd_ip.t3 dvss 0.104436f
C1191 dvdd_ip.n85 dvss 0.362629f
C1192 dvdd_ip.n86 dvss 0.362629f
C1193 dvdd_ip.t0 dvss 0.378548f
C1194 dvdd_ip.t35 dvss 0.378548f
C1195 dvdd_ip.n87 dvss 0.058833f
C1196 dvdd_ip.n88 dvss 0.244079f
C1197 dvdd_ip.n89 dvss 0.058833f
C1198 dvdd_ip.n90 dvss 0.300628f
C1199 dvdd_ip.n91 dvss 0.242337f
C1200 dvdd_ip.n92 dvss 0.35259f
C1201 dvdd_ip.n93 dvss 0.659441f
C1202 dvdd_ip.n94 dvss 0.754876f
C1203 dvdd_ip.n95 dvss 0.092315f
C1204 dvdd_ip.n96 dvss 1.14476f
C1205 dvdd_ip.n97 dvss 1.14476f
C1206 dvdd_ip.t52 dvss 1.45869f
C1207 dvdd_ip.t54 dvss 1.18277f
C1208 dvdd_ip.n98 dvss 0.235453f
C1209 dvdd_ip.t49 dvss 1.45869f
C1210 dvdd_ip.t38 dvss 1.18277f
C1211 dvdd_ip.n99 dvss 0.788516f
C1212 dvdd_ip.n100 dvss 0.235453f
C1213 dvdd_ip.n101 dvss 0.303409f
C1214 dvdd_ip.t42 dvss 0.01337f
C1215 dvdd_ip.n102 dvss 0.105974f
C1216 dvdd_ip.n104 dvss 0.50155f
C1217 dvdd_ip.t41 dvss 1.29083f
C1218 dvdd_ip.n107 dvss 0.096406f
C1219 dvdd_ip.n108 dvss 0.462744f
C1220 dvdd_ip.t32 dvss 0.053882f
C1221 dvdd_ip.t16 dvss 0.053836f
C1222 dvdd_ip.t14 dvss 0.053947f
C1223 dvdd_ip.t26 dvss 0.053774f
C1224 dvdd_ip.n109 dvss 0.974626f
C1225 dvdd_ip.t5 dvss 1.57869f
C1226 dvdd_ip.t19 dvss 1.93001f
C1227 dvdd_ip.t13 dvss 1.93001f
C1228 dvdd_ip.t15 dvss 1.44751f
C1229 dvdd_ip.n110 dvss 0.965004f
C1230 dvdd_ip.t23 dvss 1.44751f
C1231 dvdd_ip.t8 dvss 1.93001f
C1232 dvdd_ip.t17 dvss 1.93001f
C1233 dvdd_ip.t10 dvss 1.57869f
C1234 dvdd_ip.n111 dvss 0.97316f
C1235 vbp.n0 dvss 0.600345f
C1236 vbp.t11 dvss 0.764244f
C1237 vbp.n1 dvss 0.609664f
C1238 vbp.n2 dvss 0.707943f
C1239 vbp.t4 dvss 0.742966f
C1240 vbp.t6 dvss 0.742966f
C1241 vbp.n3 dvss 0.569145f
C1242 vbp.t3 dvss 0.760583f
C1243 vbp.n4 dvss 0.593784f
C1244 vbp.t13 dvss 0.895585f
C1245 vbp.n5 dvss 0.569145f
C1246 vbp.t14 dvss 0.742966f
C1247 vbp.t8 dvss 0.742966f
C1248 vbp.n6 dvss 0.569145f
C1249 vbp.t1 dvss 0.742966f
C1250 vbp.t5 dvss 0.742966f
C1251 vbp.n7 dvss 0.569145f
C1252 vbp.t10 dvss 0.742966f
C1253 vbp.t15 dvss 0.760684f
C1254 vbp.n8 dvss 0.594226f
C1255 vbp.t9 dvss 0.896467f
C1256 vbp.t12 dvss 0.742966f
C1257 vbp.n9 dvss 0.569145f
C1258 vbp.t2 dvss 0.742966f
C1259 vbp.t0 dvss 0.742966f
C1260 vbp.t7 dvss 0.742966f
C1261 vbp.n10 dvss 0.569145f
C1262 vbreg.n0 dvss 3.5606f
C1263 vbreg.n1 dvss 0.713613f
C1264 vbreg.n2 dvss 0.583542f
C1265 vbreg.n3 dvss 3.65749f
C1266 vbreg.n4 dvss 1.34473f
C1267 vbreg.n5 dvss 3.556f
C1268 vbreg.n6 dvss 0.687636f
C1269 vbreg.n7 dvss 0.582626f
C1270 vbreg.n8 dvss 1.213f
C1271 vbreg.n9 dvss 2.841f
C1272 vbreg.n10 dvss 0.583359f
C1273 vbreg.n11 dvss 2.61721f
C1274 vbreg.n12 dvss 0.592924f
C1275 vbreg.n14 dvss 0.594449f
C1276 vbreg.n15 dvss 0.931401f
C1277 vbreg.n16 dvss 0.93305f
C1278 vbreg.n17 dvss 0.404251f
C1279 vbreg.n18 dvss 0.93305f
C1280 vbreg.t11 dvss 1.20117f
C1281 vbreg.n19 dvss 0.931401f
C1282 vbreg.t8 dvss 0.23921f
C1283 vbreg.n20 dvss 1.79539f
C1284 vbreg.n21 dvss 12.184299f
C1285 vbreg.t4 dvss 0.228907f
C1286 vbreg.n22 dvss 1.25884f
C1287 vbreg.n23 dvss 0.616431f
C1288 vbreg.t6 dvss 1.20117f
C1289 vbreg.n24 dvss 0.662505f
C1290 vbreg.t19 dvss 1.20117f
C1291 vbreg.n25 dvss 0.404251f
C1292 vbreg.n26 dvss 0.400957f
C1293 vbreg.t20 dvss 1.20117f
C1294 vbreg.t18 dvss 1.20117f
C1295 vbreg.t15 dvss 1.20117f
C1296 vbreg.n27 dvss 1.00001f
C1297 vbreg.t16 dvss 1.20117f
C1298 vbreg.n28 dvss 0.685977f
C1299 vbreg.n29 dvss 0.530447f
C1300 vbreg.n30 dvss 0.404251f
C1301 vbreg.n31 dvss 0.710976f
C1302 vbreg.t10 dvss 1.21612f
C1303 vbreg.t13 dvss 1.20117f
C1304 vbreg.n32 dvss 1.00001f
C1305 vbreg.n33 dvss 0.085368f
C1306 vbreg.t12 dvss 1.20117f
C1307 vbreg.n34 dvss 1.00001f
C1308 vbreg.t14 dvss 1.20117f
C1309 vbreg.n35 dvss 0.692695f
C1310 vbreg.n36 dvss 1.00001f
C1311 vbreg.t9 dvss 1.20117f
C1312 vbreg.n37 dvss 0.530447f
C1313 vbreg.n38 dvss 0.661796f
C1314 vbreg.t17 dvss 1.20117f
C1315 vbreg.n39 dvss 1.00001f
C1316 vbreg.n40 dvss 0.168268f
C1317 vbreg.n41 dvss 1.00001f
C1318 vbreg.t7 dvss 0.228404f
C1319 vbreg.n42 dvss 0.815331f
C1320 vbreg.n43 dvss 0.528798f
C1321 vbreg.n44 dvss 0.404251f
C1322 vbreg.n45 dvss 1.00001f
C1323 vbreg.t22 dvss 1.20117f
C1324 vbreg.t24 dvss 1.20117f
C1325 vbreg.t25 dvss 1.20117f
C1326 vbreg.n46 dvss 1.00001f
C1327 vbreg.t21 dvss 1.20117f
C1328 vbreg.n47 dvss 0.531546f
C1329 vbreg.t23 dvss 1.21618f
C1330 vbreg.n48 dvss 1.00001f
C1331 vbreg.n49 dvss 0.085917f
C1332 vbreg.n50 dvss 1.30967f
C1333 vbreg.n51 dvss 0.705366f
C1334 vbreg.n52 dvss 0.531546f
C1335 vbreg.n53 dvss 0.404251f
C1336 vbreg.n54 dvss 0.527699f
C1337 vbreg.n55 dvss 0.527699f
C1338 vbreg.n56 dvss 0.404251f
C1339 vbreg.n57 dvss 0.55298f
C1340 vbreg.t1 dvss 0.214967f
C1341 vbreg.t3 dvss 0.228223f
C1342 vbreg.t2 dvss 0.268952f
C1343 vbreg.t0 dvss 0.218294f
C1344 vbreg.t5 dvss 0.138373f
C1345 icnode.t0 dvss 80.4574f
C1346 icnode.t1 dvss 0.042604f
C1347 ena_ip.n0 dvss 0.052729f
C1348 ena_ip.t1 dvss 0.038646f
C1349 ena_ip.n1 dvss 0.299073f
C1350 ena_ip.t14 dvss 0.312422f
C1351 ena_ip.t17 dvss 0.312179f
C1352 ena_ip.n2 dvss 0.262394f
C1353 ena_ip.n3 dvss 1.2068f
C1354 ena_ip.t2 dvss 0.357117f
C1355 ena_ip.t12 dvss 0.343909f
C1356 ena_ip.t18 dvss 0.013233f
C1357 ena_ip.t16 dvss 0.021012f
C1358 ena_ip.n4 dvss 0.040986f
C1359 ena_ip.t15 dvss 0.010303f
C1360 ena_ip.t4 dvss 0.024139f
C1361 ena_ip.n7 dvss 0.042815f
C1362 ena_ip.t10 dvss 0.013233f
C1363 ena_ip.t8 dvss 0.021012f
C1364 ena_ip.n8 dvss 0.040986f
C1365 ena_ip.t5 dvss 0.010303f
C1366 ena_ip.t13 dvss 0.024139f
C1367 ena_ip.n11 dvss 0.042815f
C1368 ena_ip.t9 dvss 0.013233f
C1369 ena_ip.t6 dvss 0.021012f
C1370 ena_ip.n12 dvss 0.040986f
C1371 ena_ip.t3 dvss 0.010303f
C1372 ena_ip.t7 dvss 0.024139f
C1373 ena_ip.n15 dvss 0.042815f
C1374 ena_ip.t19 dvss 0.025235f
C1375 ena_ip.t11 dvss 0.015832f
C1376 ena_ip.n16 dvss 0.036079f
C1377 ena_ip.n17 dvss 0.024525f
C1378 ena_ip.n18 dvss 0.153572f
C1379 ena_ip.t0 dvss 0.026873f
C1380 dvdd.t5 dvss 0.010219f
C1381 dvdd.t79 dvss 0.010219f
C1382 dvdd.n0 dvss 0.231928f
C1383 dvdd.n1 dvss 0.072142f
C1384 dvdd.n3 dvss 0.016591f
C1385 dvdd.n4 dvss 0.114981f
C1386 dvdd.n5 dvss 0.114981f
C1387 dvdd.t82 dvss 0.054184f
C1388 dvdd.t156 dvss 0.018317f
C1389 dvdd.n9 dvss 0.01366f
C1390 dvdd.n11 dvss 0.044846f
C1391 dvdd.n14 dvss 0.023491f
C1392 dvdd.n15 dvss 0.02799f
C1393 dvdd.n16 dvss 0.018549f
C1394 dvdd.t152 dvss 0.054184f
C1395 dvdd.t37 dvss 0.018317f
C1396 dvdd.n18 dvss 0.044846f
C1397 dvdd.n23 dvss 0.01366f
C1398 dvdd.n25 dvss 0.028887f
C1399 dvdd.n26 dvss 0.011759f
C1400 dvdd.n27 dvss 0.114981f
C1401 dvdd.n28 dvss 0.016591f
C1402 dvdd.n29 dvss 0.114981f
C1403 dvdd.n30 dvss 0.016604f
C1404 dvdd.t78 dvss 0.165457f
C1405 dvdd.n33 dvss 0.016604f
C1406 dvdd.n34 dvss 0.011759f
C1407 dvdd.n38 dvss 0.47343f
C1408 dvdd.n39 dvss 0.249961f
C1409 dvdd.n41 dvss 0.011759f
C1410 dvdd.n42 dvss 0.016604f
C1411 dvdd.t4 dvss 0.165457f
C1412 dvdd.n45 dvss 0.016604f
C1413 dvdd.n46 dvss 0.011759f
C1414 dvdd.n48 dvss 0.09794f
C1415 dvdd.n49 dvss 1.8472f
C1416 dvdd.t175 dvss 3.83628f
C1417 dvdd.n50 dvss 3.2293f
C1418 dvdd.n51 dvss 1.13209f
C1419 dvdd.n53 dvss 0.031923f
C1420 dvdd.n54 dvss 0.031923f
C1421 dvdd.n55 dvss 0.031923f
C1422 dvdd.n56 dvss 0.013356f
C1423 dvdd.n69 dvss 0.018557f
C1424 dvdd.n73 dvss 0.01242f
C1425 dvdd.n90 dvss 0.018557f
C1426 dvdd.n94 dvss 0.01242f
C1427 dvdd.n111 dvss 0.018557f
C1428 dvdd.n115 dvss 0.01242f
C1429 dvdd.n125 dvss 0.01532f
C1430 dvdd.n131 dvss 0.025945f
C1431 dvdd.n144 dvss 0.013253f
C1432 dvdd.n151 dvss 0.013028f
C1433 dvdd.n156 dvss 0.016464f
C1434 dvdd.n163 dvss 0.01532f
C1435 dvdd.n169 dvss 0.025945f
C1436 dvdd.n182 dvss 0.013253f
C1437 dvdd.n189 dvss 0.013028f
C1438 dvdd.n194 dvss 0.016464f
C1439 dvdd.n201 dvss 0.01532f
C1440 dvdd.n207 dvss 0.025945f
C1441 dvdd.n220 dvss 0.013253f
C1442 dvdd.n227 dvss 0.013028f
C1443 dvdd.n232 dvss 0.016464f
C1444 dvdd.n239 dvss 0.03748f
C1445 dvdd.t134 dvss 0.052336f
C1446 dvdd.t51 dvss 0.026937f
C1447 dvdd.t53 dvss 0.021088f
C1448 dvdd.t86 dvss 0.038944f
C1449 dvdd.t13 dvss 0.029092f
C1450 dvdd.t24 dvss 0.043716f
C1451 dvdd.t155 dvss 0.041869f
C1452 dvdd.t160 dvss 0.02586f
C1453 dvdd.t43 dvss 0.017548f
C1454 dvdd.n246 dvss 0.045043f
C1455 dvdd.n247 dvss 0.024385f
C1456 dvdd.n255 dvss 0.010777f
C1457 dvdd.n258 dvss 0.013019f
C1458 dvdd.n266 dvss 0.01321f
C1459 dvdd.n268 dvss 0.032777f
C1460 dvdd.n270 dvss 0.0709f
C1461 dvdd.t113 dvss 0.045327f
C1462 dvdd.t15 dvss 0.065683f
C1463 dvdd.t33 dvss 0.084139f
C1464 dvdd.n271 dvss 0.072054f
C1465 dvdd.t109 dvss 0.040441f
C1466 dvdd.t55 dvss 0.095267f
C1467 dvdd.t41 dvss 0.097439f
C1468 dvdd.t150 dvss 0.051841f
C1469 dvdd.t132 dvss 0.064869f
C1470 dvdd.t84 dvss 0.064326f
C1471 dvdd.t72 dvss 0.079797f
C1472 dvdd.t88 dvss 0.080339f
C1473 dvdd.t131 dvss 0.050212f
C1474 dvdd.t57 dvss 0.046141f
C1475 dvdd.t28 dvss 0.052112f
C1476 dvdd.t126 dvss 0.052112f
C1477 dvdd.t11 dvss 0.067311f
C1478 dvdd.t98 dvss 0.103953f
C1479 dvdd.t65 dvss 0.085768f
C1480 dvdd.t0 dvss 0.067311f
C1481 dvdd.n272 dvss 0.070697f
C1482 dvdd.t122 dvss 0.040441f
C1483 dvdd.t164 dvss 0.095267f
C1484 dvdd.t22 dvss 0.097439f
C1485 dvdd.t30 dvss 0.051841f
C1486 dvdd.t19 dvss 0.064869f
C1487 dvdd.t63 dvss 0.064326f
C1488 dvdd.t26 dvss 0.079797f
C1489 dvdd.t76 dvss 0.080339f
C1490 dvdd.t119 dvss 0.050212f
C1491 dvdd.t104 dvss 0.046141f
C1492 dvdd.t68 dvss 0.052112f
C1493 dvdd.t74 dvss 0.052112f
C1494 dvdd.t39 dvss 0.067311f
C1495 dvdd.t44 dvss 0.103953f
C1496 dvdd.t120 dvss 0.085768f
C1497 dvdd.t146 dvss 0.067311f
C1498 dvdd.n273 dvss 0.070697f
C1499 dvdd.t111 dvss 0.040441f
C1500 dvdd.t20 dvss 0.095267f
C1501 dvdd.t17 dvss 0.097439f
C1502 dvdd.t141 dvss 0.051841f
C1503 dvdd.t174 dvss 0.064869f
C1504 dvdd.t2 dvss 0.064326f
C1505 dvdd.t47 dvss 0.079797f
C1506 dvdd.t6 dvss 0.080339f
C1507 dvdd.t70 dvss 0.050212f
C1508 dvdd.t10 dvss 0.046141f
C1509 dvdd.t137 dvss 0.052112f
C1510 dvdd.t105 dvss 0.052112f
C1511 dvdd.t8 dvss 0.067311f
C1512 dvdd.t102 dvss 0.103953f
C1513 dvdd.t31 dvss 0.085768f
C1514 dvdd.t58 dvss 0.095709f
C1515 dvdd.n274 dvss 0.097883f
C1516 dvdd.n275 dvss 6.53977f
C1517 dvdd.n276 dvss 9.40408f
C1518 dvdd.t178 dvss 3.83628f
C1519 dvdd.n277 dvss 6.79779f
C1520 dvdd.t177 dvss 3.83628f
C1521 dvdd.n278 dvss 3.72992f
C1522 dvdd.t176 dvss 3.83628f
C1523 dvdd.n279 dvss 3.60793f
C1524 dvdd.n280 dvss 2.57602f
C1525 dvdd.n281 dvss 0.390563f
C1526 dvdd.t118 dvss 0.011125f
C1527 dvdd.t93 dvss 0.011125f
C1528 dvdd.n282 dvss 0.026681f
C1529 dvdd.t81 dvss 0.011125f
C1530 dvdd.t36 dvss 0.011125f
C1531 dvdd.n283 dvss 0.026681f
C1532 dvdd.n284 dvss 0.05226f
C1533 dvdd.t116 dvss 0.04055f
C1534 dvdd.n285 dvss 0.047939f
C1535 dvdd.n286 dvss 0.047799f
C1536 dvdd.n287 dvss 0.047799f
C1537 dvdd.t95 dvss 0.04055f
C1538 dvdd.t145 dvss 0.011125f
C1539 dvdd.t143 dvss 0.011125f
C1540 dvdd.n288 dvss 0.026681f
C1541 dvdd.t50 dvss 0.011125f
C1542 dvdd.t170 dvss 0.011125f
C1543 dvdd.n289 dvss 0.026681f
C1544 dvdd.n290 dvss 0.466107f
C1545 dvdd.n291 dvss 0.869136f
C1546 dvdd.n292 dvss 0.243102f
C1547 dvdd.n293 dvss 0.211035f
C1548 dvdd.t94 dvss 0.222917f
C1549 dvdd.t144 dvss 0.187598f
C1550 dvdd.t142 dvss 0.187598f
C1551 dvdd.t49 dvss 0.187598f
C1552 dvdd.t169 dvss 0.140698f
C1553 dvdd.n294 dvss 0.093799f
C1554 dvdd.t117 dvss 0.140698f
C1555 dvdd.t92 dvss 0.187598f
C1556 dvdd.t80 dvss 0.187598f
C1557 dvdd.t35 dvss 0.187598f
C1558 dvdd.t115 dvss 0.222917f
C1559 dvdd.n295 dvss 0.211035f
C1560 dvdd.n296 dvss 0.255981f
C1561 dvdd.n297 dvss 0.773905f
C1562 dvdd.n298 dvss 0.37474f
C1563 dvdd.n299 dvss 0.088468f
C1564 x7.stby_done_b.t0 dvss 0.057884f
C1565 x7.stby_done_b.n0 dvss 1.92933f
C1566 x7.stby_done_b.t5 dvss 0.028593f
C1567 x7.stby_done_b.t7 dvss 0.017955f
C1568 x7.stby_done_b.n1 dvss 0.038437f
C1569 x7.stby_done_b.n2 dvss 0.05998f
C1570 x7.stby_done_b.t4 dvss 0.015834f
C1571 x7.stby_done_b.n3 dvss 0.048959f
C1572 x7.stby_done_b.t3 dvss 0.015657f
C1573 x7.stby_done_b.n4 dvss 0.044896f
C1574 x7.stby_done_b.n5 dvss 0.047435f
C1575 x7.stby_done_b.t2 dvss 0.02131f
C1576 x7.stby_done_b.t6 dvss 0.023458f
C1577 x7.stby_done_b.n6 dvss 0.067085f
C1578 x7.stby_done_b.n7 dvss 1.67028f
C1579 x7.stby_done_b.n8 dvss 0.069954f
C1580 x7.stby_done_b.t1 dvss 0.043534f
.ends

