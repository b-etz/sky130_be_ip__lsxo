magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< pwell >>
rect -4268 -5782 4268 5782
<< psubdiff >>
rect -4232 5712 -4136 5746
rect 4136 5712 4232 5746
rect -4232 5650 -4198 5712
rect 4198 5650 4232 5712
rect -4232 -5712 -4198 -5650
rect 4198 -5712 4232 -5650
rect -4232 -5746 -4136 -5712
rect 4136 -5746 4232 -5712
<< psubdiffcont >>
rect -4136 5712 4136 5746
rect -4232 -5650 -4198 5650
rect 4198 -5650 4232 5650
rect -4136 -5746 4136 -5712
<< xpolycontact >>
rect -4102 5184 -4032 5616
rect -4102 -5616 -4032 -5184
rect -3936 5184 -3866 5616
rect -3936 -5616 -3866 -5184
rect -3770 5184 -3700 5616
rect -3770 -5616 -3700 -5184
rect -3604 5184 -3534 5616
rect -3604 -5616 -3534 -5184
rect -3438 5184 -3368 5616
rect -3438 -5616 -3368 -5184
rect -3272 5184 -3202 5616
rect -3272 -5616 -3202 -5184
rect -3106 5184 -3036 5616
rect -3106 -5616 -3036 -5184
rect -2940 5184 -2870 5616
rect -2940 -5616 -2870 -5184
rect -2774 5184 -2704 5616
rect -2774 -5616 -2704 -5184
rect -2608 5184 -2538 5616
rect -2608 -5616 -2538 -5184
rect -2442 5184 -2372 5616
rect -2442 -5616 -2372 -5184
rect -2276 5184 -2206 5616
rect -2276 -5616 -2206 -5184
rect -2110 5184 -2040 5616
rect -2110 -5616 -2040 -5184
rect -1944 5184 -1874 5616
rect -1944 -5616 -1874 -5184
rect -1778 5184 -1708 5616
rect -1778 -5616 -1708 -5184
rect -1612 5184 -1542 5616
rect -1612 -5616 -1542 -5184
rect -1446 5184 -1376 5616
rect -1446 -5616 -1376 -5184
rect -1280 5184 -1210 5616
rect -1280 -5616 -1210 -5184
rect -1114 5184 -1044 5616
rect -1114 -5616 -1044 -5184
rect -948 5184 -878 5616
rect -948 -5616 -878 -5184
rect -782 5184 -712 5616
rect -782 -5616 -712 -5184
rect -616 5184 -546 5616
rect -616 -5616 -546 -5184
rect -450 5184 -380 5616
rect -450 -5616 -380 -5184
rect -284 5184 -214 5616
rect -284 -5616 -214 -5184
rect -118 5184 -48 5616
rect -118 -5616 -48 -5184
rect 48 5184 118 5616
rect 48 -5616 118 -5184
rect 214 5184 284 5616
rect 214 -5616 284 -5184
rect 380 5184 450 5616
rect 380 -5616 450 -5184
rect 546 5184 616 5616
rect 546 -5616 616 -5184
rect 712 5184 782 5616
rect 712 -5616 782 -5184
rect 878 5184 948 5616
rect 878 -5616 948 -5184
rect 1044 5184 1114 5616
rect 1044 -5616 1114 -5184
rect 1210 5184 1280 5616
rect 1210 -5616 1280 -5184
rect 1376 5184 1446 5616
rect 1376 -5616 1446 -5184
rect 1542 5184 1612 5616
rect 1542 -5616 1612 -5184
rect 1708 5184 1778 5616
rect 1708 -5616 1778 -5184
rect 1874 5184 1944 5616
rect 1874 -5616 1944 -5184
rect 2040 5184 2110 5616
rect 2040 -5616 2110 -5184
rect 2206 5184 2276 5616
rect 2206 -5616 2276 -5184
rect 2372 5184 2442 5616
rect 2372 -5616 2442 -5184
rect 2538 5184 2608 5616
rect 2538 -5616 2608 -5184
rect 2704 5184 2774 5616
rect 2704 -5616 2774 -5184
rect 2870 5184 2940 5616
rect 2870 -5616 2940 -5184
rect 3036 5184 3106 5616
rect 3036 -5616 3106 -5184
rect 3202 5184 3272 5616
rect 3202 -5616 3272 -5184
rect 3368 5184 3438 5616
rect 3368 -5616 3438 -5184
rect 3534 5184 3604 5616
rect 3534 -5616 3604 -5184
rect 3700 5184 3770 5616
rect 3700 -5616 3770 -5184
rect 3866 5184 3936 5616
rect 3866 -5616 3936 -5184
rect 4032 5184 4102 5616
rect 4032 -5616 4102 -5184
<< xpolyres >>
rect -4102 -5184 -4032 5184
rect -3936 -5184 -3866 5184
rect -3770 -5184 -3700 5184
rect -3604 -5184 -3534 5184
rect -3438 -5184 -3368 5184
rect -3272 -5184 -3202 5184
rect -3106 -5184 -3036 5184
rect -2940 -5184 -2870 5184
rect -2774 -5184 -2704 5184
rect -2608 -5184 -2538 5184
rect -2442 -5184 -2372 5184
rect -2276 -5184 -2206 5184
rect -2110 -5184 -2040 5184
rect -1944 -5184 -1874 5184
rect -1778 -5184 -1708 5184
rect -1612 -5184 -1542 5184
rect -1446 -5184 -1376 5184
rect -1280 -5184 -1210 5184
rect -1114 -5184 -1044 5184
rect -948 -5184 -878 5184
rect -782 -5184 -712 5184
rect -616 -5184 -546 5184
rect -450 -5184 -380 5184
rect -284 -5184 -214 5184
rect -118 -5184 -48 5184
rect 48 -5184 118 5184
rect 214 -5184 284 5184
rect 380 -5184 450 5184
rect 546 -5184 616 5184
rect 712 -5184 782 5184
rect 878 -5184 948 5184
rect 1044 -5184 1114 5184
rect 1210 -5184 1280 5184
rect 1376 -5184 1446 5184
rect 1542 -5184 1612 5184
rect 1708 -5184 1778 5184
rect 1874 -5184 1944 5184
rect 2040 -5184 2110 5184
rect 2206 -5184 2276 5184
rect 2372 -5184 2442 5184
rect 2538 -5184 2608 5184
rect 2704 -5184 2774 5184
rect 2870 -5184 2940 5184
rect 3036 -5184 3106 5184
rect 3202 -5184 3272 5184
rect 3368 -5184 3438 5184
rect 3534 -5184 3604 5184
rect 3700 -5184 3770 5184
rect 3866 -5184 3936 5184
rect 4032 -5184 4102 5184
<< locali >>
rect -4232 5712 -4136 5746
rect 4136 5712 4232 5746
rect -4232 5650 -4198 5712
rect 4198 5650 4232 5712
rect -4232 -5712 -4198 -5650
rect 4198 -5712 4232 -5650
rect -4232 -5746 -4136 -5712
rect 4136 -5746 4232 -5712
<< viali >>
rect -4086 5201 -4048 5598
rect -3920 5201 -3882 5598
rect -3754 5201 -3716 5598
rect -3588 5201 -3550 5598
rect -3422 5201 -3384 5598
rect -3256 5201 -3218 5598
rect -3090 5201 -3052 5598
rect -2924 5201 -2886 5598
rect -2758 5201 -2720 5598
rect -2592 5201 -2554 5598
rect -2426 5201 -2388 5598
rect -2260 5201 -2222 5598
rect -2094 5201 -2056 5598
rect -1928 5201 -1890 5598
rect -1762 5201 -1724 5598
rect -1596 5201 -1558 5598
rect -1430 5201 -1392 5598
rect -1264 5201 -1226 5598
rect -1098 5201 -1060 5598
rect -932 5201 -894 5598
rect -766 5201 -728 5598
rect -600 5201 -562 5598
rect -434 5201 -396 5598
rect -268 5201 -230 5598
rect -102 5201 -64 5598
rect 64 5201 102 5598
rect 230 5201 268 5598
rect 396 5201 434 5598
rect 562 5201 600 5598
rect 728 5201 766 5598
rect 894 5201 932 5598
rect 1060 5201 1098 5598
rect 1226 5201 1264 5598
rect 1392 5201 1430 5598
rect 1558 5201 1596 5598
rect 1724 5201 1762 5598
rect 1890 5201 1928 5598
rect 2056 5201 2094 5598
rect 2222 5201 2260 5598
rect 2388 5201 2426 5598
rect 2554 5201 2592 5598
rect 2720 5201 2758 5598
rect 2886 5201 2924 5598
rect 3052 5201 3090 5598
rect 3218 5201 3256 5598
rect 3384 5201 3422 5598
rect 3550 5201 3588 5598
rect 3716 5201 3754 5598
rect 3882 5201 3920 5598
rect 4048 5201 4086 5598
rect -4086 -5598 -4048 -5201
rect -3920 -5598 -3882 -5201
rect -3754 -5598 -3716 -5201
rect -3588 -5598 -3550 -5201
rect -3422 -5598 -3384 -5201
rect -3256 -5598 -3218 -5201
rect -3090 -5598 -3052 -5201
rect -2924 -5598 -2886 -5201
rect -2758 -5598 -2720 -5201
rect -2592 -5598 -2554 -5201
rect -2426 -5598 -2388 -5201
rect -2260 -5598 -2222 -5201
rect -2094 -5598 -2056 -5201
rect -1928 -5598 -1890 -5201
rect -1762 -5598 -1724 -5201
rect -1596 -5598 -1558 -5201
rect -1430 -5598 -1392 -5201
rect -1264 -5598 -1226 -5201
rect -1098 -5598 -1060 -5201
rect -932 -5598 -894 -5201
rect -766 -5598 -728 -5201
rect -600 -5598 -562 -5201
rect -434 -5598 -396 -5201
rect -268 -5598 -230 -5201
rect -102 -5598 -64 -5201
rect 64 -5598 102 -5201
rect 230 -5598 268 -5201
rect 396 -5598 434 -5201
rect 562 -5598 600 -5201
rect 728 -5598 766 -5201
rect 894 -5598 932 -5201
rect 1060 -5598 1098 -5201
rect 1226 -5598 1264 -5201
rect 1392 -5598 1430 -5201
rect 1558 -5598 1596 -5201
rect 1724 -5598 1762 -5201
rect 1890 -5598 1928 -5201
rect 2056 -5598 2094 -5201
rect 2222 -5598 2260 -5201
rect 2388 -5598 2426 -5201
rect 2554 -5598 2592 -5201
rect 2720 -5598 2758 -5201
rect 2886 -5598 2924 -5201
rect 3052 -5598 3090 -5201
rect 3218 -5598 3256 -5201
rect 3384 -5598 3422 -5201
rect 3550 -5598 3588 -5201
rect 3716 -5598 3754 -5201
rect 3882 -5598 3920 -5201
rect 4048 -5598 4086 -5201
<< metal1 >>
rect -4092 5598 -4042 5610
rect -4092 5201 -4086 5598
rect -4048 5201 -4042 5598
rect -4092 5189 -4042 5201
rect -3926 5598 -3876 5610
rect -3926 5201 -3920 5598
rect -3882 5201 -3876 5598
rect -3926 5189 -3876 5201
rect -3760 5598 -3710 5610
rect -3760 5201 -3754 5598
rect -3716 5201 -3710 5598
rect -3760 5189 -3710 5201
rect -3594 5598 -3544 5610
rect -3594 5201 -3588 5598
rect -3550 5201 -3544 5598
rect -3594 5189 -3544 5201
rect -3428 5598 -3378 5610
rect -3428 5201 -3422 5598
rect -3384 5201 -3378 5598
rect -3428 5189 -3378 5201
rect -3262 5598 -3212 5610
rect -3262 5201 -3256 5598
rect -3218 5201 -3212 5598
rect -3262 5189 -3212 5201
rect -3096 5598 -3046 5610
rect -3096 5201 -3090 5598
rect -3052 5201 -3046 5598
rect -3096 5189 -3046 5201
rect -2930 5598 -2880 5610
rect -2930 5201 -2924 5598
rect -2886 5201 -2880 5598
rect -2930 5189 -2880 5201
rect -2764 5598 -2714 5610
rect -2764 5201 -2758 5598
rect -2720 5201 -2714 5598
rect -2764 5189 -2714 5201
rect -2598 5598 -2548 5610
rect -2598 5201 -2592 5598
rect -2554 5201 -2548 5598
rect -2598 5189 -2548 5201
rect -2432 5598 -2382 5610
rect -2432 5201 -2426 5598
rect -2388 5201 -2382 5598
rect -2432 5189 -2382 5201
rect -2266 5598 -2216 5610
rect -2266 5201 -2260 5598
rect -2222 5201 -2216 5598
rect -2266 5189 -2216 5201
rect -2100 5598 -2050 5610
rect -2100 5201 -2094 5598
rect -2056 5201 -2050 5598
rect -2100 5189 -2050 5201
rect -1934 5598 -1884 5610
rect -1934 5201 -1928 5598
rect -1890 5201 -1884 5598
rect -1934 5189 -1884 5201
rect -1768 5598 -1718 5610
rect -1768 5201 -1762 5598
rect -1724 5201 -1718 5598
rect -1768 5189 -1718 5201
rect -1602 5598 -1552 5610
rect -1602 5201 -1596 5598
rect -1558 5201 -1552 5598
rect -1602 5189 -1552 5201
rect -1436 5598 -1386 5610
rect -1436 5201 -1430 5598
rect -1392 5201 -1386 5598
rect -1436 5189 -1386 5201
rect -1270 5598 -1220 5610
rect -1270 5201 -1264 5598
rect -1226 5201 -1220 5598
rect -1270 5189 -1220 5201
rect -1104 5598 -1054 5610
rect -1104 5201 -1098 5598
rect -1060 5201 -1054 5598
rect -1104 5189 -1054 5201
rect -938 5598 -888 5610
rect -938 5201 -932 5598
rect -894 5201 -888 5598
rect -938 5189 -888 5201
rect -772 5598 -722 5610
rect -772 5201 -766 5598
rect -728 5201 -722 5598
rect -772 5189 -722 5201
rect -606 5598 -556 5610
rect -606 5201 -600 5598
rect -562 5201 -556 5598
rect -606 5189 -556 5201
rect -440 5598 -390 5610
rect -440 5201 -434 5598
rect -396 5201 -390 5598
rect -440 5189 -390 5201
rect -274 5598 -224 5610
rect -274 5201 -268 5598
rect -230 5201 -224 5598
rect -274 5189 -224 5201
rect -108 5598 -58 5610
rect -108 5201 -102 5598
rect -64 5201 -58 5598
rect -108 5189 -58 5201
rect 58 5598 108 5610
rect 58 5201 64 5598
rect 102 5201 108 5598
rect 58 5189 108 5201
rect 224 5598 274 5610
rect 224 5201 230 5598
rect 268 5201 274 5598
rect 224 5189 274 5201
rect 390 5598 440 5610
rect 390 5201 396 5598
rect 434 5201 440 5598
rect 390 5189 440 5201
rect 556 5598 606 5610
rect 556 5201 562 5598
rect 600 5201 606 5598
rect 556 5189 606 5201
rect 722 5598 772 5610
rect 722 5201 728 5598
rect 766 5201 772 5598
rect 722 5189 772 5201
rect 888 5598 938 5610
rect 888 5201 894 5598
rect 932 5201 938 5598
rect 888 5189 938 5201
rect 1054 5598 1104 5610
rect 1054 5201 1060 5598
rect 1098 5201 1104 5598
rect 1054 5189 1104 5201
rect 1220 5598 1270 5610
rect 1220 5201 1226 5598
rect 1264 5201 1270 5598
rect 1220 5189 1270 5201
rect 1386 5598 1436 5610
rect 1386 5201 1392 5598
rect 1430 5201 1436 5598
rect 1386 5189 1436 5201
rect 1552 5598 1602 5610
rect 1552 5201 1558 5598
rect 1596 5201 1602 5598
rect 1552 5189 1602 5201
rect 1718 5598 1768 5610
rect 1718 5201 1724 5598
rect 1762 5201 1768 5598
rect 1718 5189 1768 5201
rect 1884 5598 1934 5610
rect 1884 5201 1890 5598
rect 1928 5201 1934 5598
rect 1884 5189 1934 5201
rect 2050 5598 2100 5610
rect 2050 5201 2056 5598
rect 2094 5201 2100 5598
rect 2050 5189 2100 5201
rect 2216 5598 2266 5610
rect 2216 5201 2222 5598
rect 2260 5201 2266 5598
rect 2216 5189 2266 5201
rect 2382 5598 2432 5610
rect 2382 5201 2388 5598
rect 2426 5201 2432 5598
rect 2382 5189 2432 5201
rect 2548 5598 2598 5610
rect 2548 5201 2554 5598
rect 2592 5201 2598 5598
rect 2548 5189 2598 5201
rect 2714 5598 2764 5610
rect 2714 5201 2720 5598
rect 2758 5201 2764 5598
rect 2714 5189 2764 5201
rect 2880 5598 2930 5610
rect 2880 5201 2886 5598
rect 2924 5201 2930 5598
rect 2880 5189 2930 5201
rect 3046 5598 3096 5610
rect 3046 5201 3052 5598
rect 3090 5201 3096 5598
rect 3046 5189 3096 5201
rect 3212 5598 3262 5610
rect 3212 5201 3218 5598
rect 3256 5201 3262 5598
rect 3212 5189 3262 5201
rect 3378 5598 3428 5610
rect 3378 5201 3384 5598
rect 3422 5201 3428 5598
rect 3378 5189 3428 5201
rect 3544 5598 3594 5610
rect 3544 5201 3550 5598
rect 3588 5201 3594 5598
rect 3544 5189 3594 5201
rect 3710 5598 3760 5610
rect 3710 5201 3716 5598
rect 3754 5201 3760 5598
rect 3710 5189 3760 5201
rect 3876 5598 3926 5610
rect 3876 5201 3882 5598
rect 3920 5201 3926 5598
rect 3876 5189 3926 5201
rect 4042 5598 4092 5610
rect 4042 5201 4048 5598
rect 4086 5201 4092 5598
rect 4042 5189 4092 5201
rect -4092 -5201 -4042 -5189
rect -4092 -5598 -4086 -5201
rect -4048 -5598 -4042 -5201
rect -4092 -5610 -4042 -5598
rect -3926 -5201 -3876 -5189
rect -3926 -5598 -3920 -5201
rect -3882 -5598 -3876 -5201
rect -3926 -5610 -3876 -5598
rect -3760 -5201 -3710 -5189
rect -3760 -5598 -3754 -5201
rect -3716 -5598 -3710 -5201
rect -3760 -5610 -3710 -5598
rect -3594 -5201 -3544 -5189
rect -3594 -5598 -3588 -5201
rect -3550 -5598 -3544 -5201
rect -3594 -5610 -3544 -5598
rect -3428 -5201 -3378 -5189
rect -3428 -5598 -3422 -5201
rect -3384 -5598 -3378 -5201
rect -3428 -5610 -3378 -5598
rect -3262 -5201 -3212 -5189
rect -3262 -5598 -3256 -5201
rect -3218 -5598 -3212 -5201
rect -3262 -5610 -3212 -5598
rect -3096 -5201 -3046 -5189
rect -3096 -5598 -3090 -5201
rect -3052 -5598 -3046 -5201
rect -3096 -5610 -3046 -5598
rect -2930 -5201 -2880 -5189
rect -2930 -5598 -2924 -5201
rect -2886 -5598 -2880 -5201
rect -2930 -5610 -2880 -5598
rect -2764 -5201 -2714 -5189
rect -2764 -5598 -2758 -5201
rect -2720 -5598 -2714 -5201
rect -2764 -5610 -2714 -5598
rect -2598 -5201 -2548 -5189
rect -2598 -5598 -2592 -5201
rect -2554 -5598 -2548 -5201
rect -2598 -5610 -2548 -5598
rect -2432 -5201 -2382 -5189
rect -2432 -5598 -2426 -5201
rect -2388 -5598 -2382 -5201
rect -2432 -5610 -2382 -5598
rect -2266 -5201 -2216 -5189
rect -2266 -5598 -2260 -5201
rect -2222 -5598 -2216 -5201
rect -2266 -5610 -2216 -5598
rect -2100 -5201 -2050 -5189
rect -2100 -5598 -2094 -5201
rect -2056 -5598 -2050 -5201
rect -2100 -5610 -2050 -5598
rect -1934 -5201 -1884 -5189
rect -1934 -5598 -1928 -5201
rect -1890 -5598 -1884 -5201
rect -1934 -5610 -1884 -5598
rect -1768 -5201 -1718 -5189
rect -1768 -5598 -1762 -5201
rect -1724 -5598 -1718 -5201
rect -1768 -5610 -1718 -5598
rect -1602 -5201 -1552 -5189
rect -1602 -5598 -1596 -5201
rect -1558 -5598 -1552 -5201
rect -1602 -5610 -1552 -5598
rect -1436 -5201 -1386 -5189
rect -1436 -5598 -1430 -5201
rect -1392 -5598 -1386 -5201
rect -1436 -5610 -1386 -5598
rect -1270 -5201 -1220 -5189
rect -1270 -5598 -1264 -5201
rect -1226 -5598 -1220 -5201
rect -1270 -5610 -1220 -5598
rect -1104 -5201 -1054 -5189
rect -1104 -5598 -1098 -5201
rect -1060 -5598 -1054 -5201
rect -1104 -5610 -1054 -5598
rect -938 -5201 -888 -5189
rect -938 -5598 -932 -5201
rect -894 -5598 -888 -5201
rect -938 -5610 -888 -5598
rect -772 -5201 -722 -5189
rect -772 -5598 -766 -5201
rect -728 -5598 -722 -5201
rect -772 -5610 -722 -5598
rect -606 -5201 -556 -5189
rect -606 -5598 -600 -5201
rect -562 -5598 -556 -5201
rect -606 -5610 -556 -5598
rect -440 -5201 -390 -5189
rect -440 -5598 -434 -5201
rect -396 -5598 -390 -5201
rect -440 -5610 -390 -5598
rect -274 -5201 -224 -5189
rect -274 -5598 -268 -5201
rect -230 -5598 -224 -5201
rect -274 -5610 -224 -5598
rect -108 -5201 -58 -5189
rect -108 -5598 -102 -5201
rect -64 -5598 -58 -5201
rect -108 -5610 -58 -5598
rect 58 -5201 108 -5189
rect 58 -5598 64 -5201
rect 102 -5598 108 -5201
rect 58 -5610 108 -5598
rect 224 -5201 274 -5189
rect 224 -5598 230 -5201
rect 268 -5598 274 -5201
rect 224 -5610 274 -5598
rect 390 -5201 440 -5189
rect 390 -5598 396 -5201
rect 434 -5598 440 -5201
rect 390 -5610 440 -5598
rect 556 -5201 606 -5189
rect 556 -5598 562 -5201
rect 600 -5598 606 -5201
rect 556 -5610 606 -5598
rect 722 -5201 772 -5189
rect 722 -5598 728 -5201
rect 766 -5598 772 -5201
rect 722 -5610 772 -5598
rect 888 -5201 938 -5189
rect 888 -5598 894 -5201
rect 932 -5598 938 -5201
rect 888 -5610 938 -5598
rect 1054 -5201 1104 -5189
rect 1054 -5598 1060 -5201
rect 1098 -5598 1104 -5201
rect 1054 -5610 1104 -5598
rect 1220 -5201 1270 -5189
rect 1220 -5598 1226 -5201
rect 1264 -5598 1270 -5201
rect 1220 -5610 1270 -5598
rect 1386 -5201 1436 -5189
rect 1386 -5598 1392 -5201
rect 1430 -5598 1436 -5201
rect 1386 -5610 1436 -5598
rect 1552 -5201 1602 -5189
rect 1552 -5598 1558 -5201
rect 1596 -5598 1602 -5201
rect 1552 -5610 1602 -5598
rect 1718 -5201 1768 -5189
rect 1718 -5598 1724 -5201
rect 1762 -5598 1768 -5201
rect 1718 -5610 1768 -5598
rect 1884 -5201 1934 -5189
rect 1884 -5598 1890 -5201
rect 1928 -5598 1934 -5201
rect 1884 -5610 1934 -5598
rect 2050 -5201 2100 -5189
rect 2050 -5598 2056 -5201
rect 2094 -5598 2100 -5201
rect 2050 -5610 2100 -5598
rect 2216 -5201 2266 -5189
rect 2216 -5598 2222 -5201
rect 2260 -5598 2266 -5201
rect 2216 -5610 2266 -5598
rect 2382 -5201 2432 -5189
rect 2382 -5598 2388 -5201
rect 2426 -5598 2432 -5201
rect 2382 -5610 2432 -5598
rect 2548 -5201 2598 -5189
rect 2548 -5598 2554 -5201
rect 2592 -5598 2598 -5201
rect 2548 -5610 2598 -5598
rect 2714 -5201 2764 -5189
rect 2714 -5598 2720 -5201
rect 2758 -5598 2764 -5201
rect 2714 -5610 2764 -5598
rect 2880 -5201 2930 -5189
rect 2880 -5598 2886 -5201
rect 2924 -5598 2930 -5201
rect 2880 -5610 2930 -5598
rect 3046 -5201 3096 -5189
rect 3046 -5598 3052 -5201
rect 3090 -5598 3096 -5201
rect 3046 -5610 3096 -5598
rect 3212 -5201 3262 -5189
rect 3212 -5598 3218 -5201
rect 3256 -5598 3262 -5201
rect 3212 -5610 3262 -5598
rect 3378 -5201 3428 -5189
rect 3378 -5598 3384 -5201
rect 3422 -5598 3428 -5201
rect 3378 -5610 3428 -5598
rect 3544 -5201 3594 -5189
rect 3544 -5598 3550 -5201
rect 3588 -5598 3594 -5201
rect 3544 -5610 3594 -5598
rect 3710 -5201 3760 -5189
rect 3710 -5598 3716 -5201
rect 3754 -5598 3760 -5201
rect 3710 -5610 3760 -5598
rect 3876 -5201 3926 -5189
rect 3876 -5598 3882 -5201
rect 3920 -5598 3926 -5201
rect 3876 -5610 3926 -5598
rect 4042 -5201 4092 -5189
rect 4042 -5598 4048 -5201
rect 4086 -5598 4092 -5201
rect 4042 -5610 4092 -5598
<< properties >>
string FIXED_BBOX -4215 -5729 4215 5729
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 52.0 m 1 nx 50 wmin 0.350 lmin 0.50 rho 2000 val 298.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
