magic
tech sky130A
magscale 1 2
timestamp 1712853061
use sky130_fd_pr__cap_mim_m3_1_4MNTN9  XC1
timestamp 1712853061
transform 0 1 3490 -1 0 -8940
box -2492 -6960 2492 6960
use sky130_fd_pr__nfet_g5v0d10v5_LNU7CV  XM1_2
timestamp 1712853061
transform 1 0 2845 0 1 -1484
box -2031 -458 2031 458
use sky130_fd_pr__nfet_01v8_ZWWV9A  XM4_18
timestamp 1712853061
transform 1 0 7787 0 1 -5736
box -1083 -610 1083 610
use sky130_fd_pr__pfet_g5v0d10v5_47BKFH  XM5
timestamp 1712782684
transform 1 0 7743 0 1 -3749
box -1145 -697 1145 697
use sky130_fd_pr__pfet_01v8_CQSSVD  XM6
timestamp 1712071977
transform 1 0 13800 0 1 -10163
box -996 -269 996 269
use sky130_fd_pr__nfet_01v8_FMHZDY  XM7
timestamp 1712071977
transform 1 0 13798 0 1 -10738
box -996 -260 996 260
use sky130_fd_pr__pfet_01v8_CQSSVD  XM8
timestamp 1712071977
transform 1 0 11914 0 1 -10163
box -996 -269 996 269
use sky130_fd_pr__nfet_01v8_FMHZDY  XM9
timestamp 1712071977
transform 1 0 11912 0 1 -10738
box -996 -260 996 260
use sky130_fd_pr__pfet_01v8_FQSSVM  XM10
timestamp 1712071977
transform 1 0 15786 0 1 -10173
box -296 -269 296 269
use sky130_fd_pr__nfet_01v8_FMMQLY  XM11
timestamp 1712071977
transform 1 0 15772 0 1 -11240
box -296 -260 296 260
use sky130_fd_pr__pfet_01v8_3HMWVM  XM12
timestamp 1712071977
transform 1 0 16686 0 1 -10039
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_69TQ3K  XM13
timestamp 1712071977
transform 1 0 16672 0 1 -10976
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_ZMTD9P  XM16_17
timestamp 1712853061
transform 1 0 2843 0 1 -2755
box -1999 -683 1999 683
use sky130_fd_pr__res_xhigh_po_0p35_TYV4QT  XR1
timestamp 1712071977
transform 1 0 13097 0 1 -5190
box -2193 -4582 2193 4582
<< end >>
