magic
tech sky130A
magscale 1 2
timestamp 1712930846
<< nwell >>
rect -2061 -761 2061 761
<< mvpmos >>
rect -1803 64 -1403 464
rect -1345 64 -945 464
rect -887 64 -487 464
rect -429 64 -29 464
rect 29 64 429 464
rect 487 64 887 464
rect 945 64 1345 464
rect 1403 64 1803 464
rect -1803 -464 -1403 -64
rect -1345 -464 -945 -64
rect -887 -464 -487 -64
rect -429 -464 -29 -64
rect 29 -464 429 -64
rect 487 -464 887 -64
rect 945 -464 1345 -64
rect 1403 -464 1803 -64
<< mvpdiff >>
rect -1861 452 -1803 464
rect -1861 76 -1849 452
rect -1815 76 -1803 452
rect -1861 64 -1803 76
rect -1403 452 -1345 464
rect -1403 76 -1391 452
rect -1357 76 -1345 452
rect -1403 64 -1345 76
rect -945 452 -887 464
rect -945 76 -933 452
rect -899 76 -887 452
rect -945 64 -887 76
rect -487 452 -429 464
rect -487 76 -475 452
rect -441 76 -429 452
rect -487 64 -429 76
rect -29 452 29 464
rect -29 76 -17 452
rect 17 76 29 452
rect -29 64 29 76
rect 429 452 487 464
rect 429 76 441 452
rect 475 76 487 452
rect 429 64 487 76
rect 887 452 945 464
rect 887 76 899 452
rect 933 76 945 452
rect 887 64 945 76
rect 1345 452 1403 464
rect 1345 76 1357 452
rect 1391 76 1403 452
rect 1345 64 1403 76
rect 1803 452 1861 464
rect 1803 76 1815 452
rect 1849 76 1861 452
rect 1803 64 1861 76
rect -1861 -76 -1803 -64
rect -1861 -452 -1849 -76
rect -1815 -452 -1803 -76
rect -1861 -464 -1803 -452
rect -1403 -76 -1345 -64
rect -1403 -452 -1391 -76
rect -1357 -452 -1345 -76
rect -1403 -464 -1345 -452
rect -945 -76 -887 -64
rect -945 -452 -933 -76
rect -899 -452 -887 -76
rect -945 -464 -887 -452
rect -487 -76 -429 -64
rect -487 -452 -475 -76
rect -441 -452 -429 -76
rect -487 -464 -429 -452
rect -29 -76 29 -64
rect -29 -452 -17 -76
rect 17 -452 29 -76
rect -29 -464 29 -452
rect 429 -76 487 -64
rect 429 -452 441 -76
rect 475 -452 487 -76
rect 429 -464 487 -452
rect 887 -76 945 -64
rect 887 -452 899 -76
rect 933 -452 945 -76
rect 887 -464 945 -452
rect 1345 -76 1403 -64
rect 1345 -452 1357 -76
rect 1391 -452 1403 -76
rect 1345 -464 1403 -452
rect 1803 -76 1861 -64
rect 1803 -452 1815 -76
rect 1849 -452 1861 -76
rect 1803 -464 1861 -452
<< mvpdiffc >>
rect -1849 76 -1815 452
rect -1391 76 -1357 452
rect -933 76 -899 452
rect -475 76 -441 452
rect -17 76 17 452
rect 441 76 475 452
rect 899 76 933 452
rect 1357 76 1391 452
rect 1815 76 1849 452
rect -1849 -452 -1815 -76
rect -1391 -452 -1357 -76
rect -933 -452 -899 -76
rect -475 -452 -441 -76
rect -17 -452 17 -76
rect 441 -452 475 -76
rect 899 -452 933 -76
rect 1357 -452 1391 -76
rect 1815 -452 1849 -76
<< mvnsubdiff >>
rect -1995 683 1995 695
rect -1995 649 -1887 683
rect 1887 649 1995 683
rect -1995 637 1995 649
rect -1995 587 -1937 637
rect -1995 -587 -1983 587
rect -1949 -587 -1937 587
rect 1937 587 1995 637
rect -1995 -637 -1937 -587
rect 1937 -587 1949 587
rect 1983 -587 1995 587
rect 1937 -637 1995 -587
rect -1995 -649 1995 -637
rect -1995 -683 -1887 -649
rect 1887 -683 1995 -649
rect -1995 -695 1995 -683
<< mvnsubdiffcont >>
rect -1887 649 1887 683
rect -1983 -587 -1949 587
rect 1949 -587 1983 587
rect -1887 -683 1887 -649
<< poly >>
rect -1803 545 -1403 561
rect -1803 511 -1787 545
rect -1419 511 -1403 545
rect -1803 464 -1403 511
rect -1345 545 -945 561
rect -1345 511 -1329 545
rect -961 511 -945 545
rect -1345 464 -945 511
rect -887 545 -487 561
rect -887 511 -871 545
rect -503 511 -487 545
rect -887 464 -487 511
rect -429 545 -29 561
rect -429 511 -413 545
rect -45 511 -29 545
rect -429 464 -29 511
rect 29 545 429 561
rect 29 511 45 545
rect 413 511 429 545
rect 29 464 429 511
rect 487 545 887 561
rect 487 511 503 545
rect 871 511 887 545
rect 487 464 887 511
rect 945 545 1345 561
rect 945 511 961 545
rect 1329 511 1345 545
rect 945 464 1345 511
rect 1403 545 1803 561
rect 1403 511 1419 545
rect 1787 511 1803 545
rect 1403 464 1803 511
rect -1803 17 -1403 64
rect -1803 -17 -1787 17
rect -1419 -17 -1403 17
rect -1803 -64 -1403 -17
rect -1345 17 -945 64
rect -1345 -17 -1329 17
rect -961 -17 -945 17
rect -1345 -64 -945 -17
rect -887 17 -487 64
rect -887 -17 -871 17
rect -503 -17 -487 17
rect -887 -64 -487 -17
rect -429 17 -29 64
rect -429 -17 -413 17
rect -45 -17 -29 17
rect -429 -64 -29 -17
rect 29 17 429 64
rect 29 -17 45 17
rect 413 -17 429 17
rect 29 -64 429 -17
rect 487 17 887 64
rect 487 -17 503 17
rect 871 -17 887 17
rect 487 -64 887 -17
rect 945 17 1345 64
rect 945 -17 961 17
rect 1329 -17 1345 17
rect 945 -64 1345 -17
rect 1403 17 1803 64
rect 1403 -17 1419 17
rect 1787 -17 1803 17
rect 1403 -64 1803 -17
rect -1803 -511 -1403 -464
rect -1803 -545 -1787 -511
rect -1419 -545 -1403 -511
rect -1803 -561 -1403 -545
rect -1345 -511 -945 -464
rect -1345 -545 -1329 -511
rect -961 -545 -945 -511
rect -1345 -561 -945 -545
rect -887 -511 -487 -464
rect -887 -545 -871 -511
rect -503 -545 -487 -511
rect -887 -561 -487 -545
rect -429 -511 -29 -464
rect -429 -545 -413 -511
rect -45 -545 -29 -511
rect -429 -561 -29 -545
rect 29 -511 429 -464
rect 29 -545 45 -511
rect 413 -545 429 -511
rect 29 -561 429 -545
rect 487 -511 887 -464
rect 487 -545 503 -511
rect 871 -545 887 -511
rect 487 -561 887 -545
rect 945 -511 1345 -464
rect 945 -545 961 -511
rect 1329 -545 1345 -511
rect 945 -561 1345 -545
rect 1403 -511 1803 -464
rect 1403 -545 1419 -511
rect 1787 -545 1803 -511
rect 1403 -561 1803 -545
<< polycont >>
rect -1787 511 -1419 545
rect -1329 511 -961 545
rect -871 511 -503 545
rect -413 511 -45 545
rect 45 511 413 545
rect 503 511 871 545
rect 961 511 1329 545
rect 1419 511 1787 545
rect -1787 -17 -1419 17
rect -1329 -17 -961 17
rect -871 -17 -503 17
rect -413 -17 -45 17
rect 45 -17 413 17
rect 503 -17 871 17
rect 961 -17 1329 17
rect 1419 -17 1787 17
rect -1787 -545 -1419 -511
rect -1329 -545 -961 -511
rect -871 -545 -503 -511
rect -413 -545 -45 -511
rect 45 -545 413 -511
rect 503 -545 871 -511
rect 961 -545 1329 -511
rect 1419 -545 1787 -511
<< locali >>
rect -1983 649 -1887 683
rect 1887 649 1983 683
rect -1983 587 -1949 649
rect 1949 587 1983 649
rect -1803 511 -1787 545
rect -1419 511 -1403 545
rect -1345 511 -1329 545
rect -961 511 -945 545
rect -887 511 -871 545
rect -503 511 -487 545
rect -429 511 -413 545
rect -45 511 -29 545
rect 29 511 45 545
rect 413 511 429 545
rect 487 511 503 545
rect 871 511 887 545
rect 945 511 961 545
rect 1329 511 1345 545
rect 1403 511 1419 545
rect 1787 511 1803 545
rect -1849 452 -1815 468
rect -1849 60 -1815 76
rect -1391 452 -1357 468
rect -1391 60 -1357 76
rect -933 452 -899 468
rect -933 60 -899 76
rect -475 452 -441 468
rect -475 60 -441 76
rect -17 452 17 468
rect -17 60 17 76
rect 441 452 475 468
rect 441 60 475 76
rect 899 452 933 468
rect 899 60 933 76
rect 1357 452 1391 468
rect 1357 60 1391 76
rect 1815 452 1849 468
rect 1815 60 1849 76
rect -1803 -17 -1787 17
rect -1419 -17 -1403 17
rect -1345 -17 -1329 17
rect -961 -17 -945 17
rect -887 -17 -871 17
rect -503 -17 -487 17
rect -429 -17 -413 17
rect -45 -17 -29 17
rect 29 -17 45 17
rect 413 -17 429 17
rect 487 -17 503 17
rect 871 -17 887 17
rect 945 -17 961 17
rect 1329 -17 1345 17
rect 1403 -17 1419 17
rect 1787 -17 1803 17
rect -1849 -76 -1815 -60
rect -1849 -468 -1815 -452
rect -1391 -76 -1357 -60
rect -1391 -468 -1357 -452
rect -933 -76 -899 -60
rect -933 -468 -899 -452
rect -475 -76 -441 -60
rect -475 -468 -441 -452
rect -17 -76 17 -60
rect -17 -468 17 -452
rect 441 -76 475 -60
rect 441 -468 475 -452
rect 899 -76 933 -60
rect 899 -468 933 -452
rect 1357 -76 1391 -60
rect 1357 -468 1391 -452
rect 1815 -76 1849 -60
rect 1815 -468 1849 -452
rect -1803 -545 -1787 -511
rect -1419 -545 -1403 -511
rect -1345 -545 -1329 -511
rect -961 -545 -945 -511
rect -887 -545 -871 -511
rect -503 -545 -487 -511
rect -429 -545 -413 -511
rect -45 -545 -29 -511
rect 29 -545 45 -511
rect 413 -545 429 -511
rect 487 -545 503 -511
rect 871 -545 887 -511
rect 945 -545 961 -511
rect 1329 -545 1345 -511
rect 1403 -545 1419 -511
rect 1787 -545 1803 -511
rect -1983 -649 -1949 -587
rect 1949 -649 1983 -587
rect -1983 -683 -1887 -649
rect 1887 -683 1983 -649
<< viali >>
rect -1787 511 -1419 545
rect -1329 511 -961 545
rect -871 511 -503 545
rect -413 511 -45 545
rect 45 511 413 545
rect 503 511 871 545
rect 961 511 1329 545
rect 1419 511 1787 545
rect -1849 76 -1815 452
rect -1391 76 -1357 452
rect -933 76 -899 452
rect -475 76 -441 452
rect -17 76 17 452
rect 441 76 475 452
rect 899 76 933 452
rect 1357 76 1391 452
rect 1815 76 1849 452
rect -1787 -17 -1419 17
rect -1329 -17 -961 17
rect -871 -17 -503 17
rect -413 -17 -45 17
rect 45 -17 413 17
rect 503 -17 871 17
rect 961 -17 1329 17
rect 1419 -17 1787 17
rect -1849 -452 -1815 -76
rect -1391 -452 -1357 -76
rect -933 -452 -899 -76
rect -475 -452 -441 -76
rect -17 -452 17 -76
rect 441 -452 475 -76
rect 899 -452 933 -76
rect 1357 -452 1391 -76
rect 1815 -452 1849 -76
rect -1787 -545 -1419 -511
rect -1329 -545 -961 -511
rect -871 -545 -503 -511
rect -413 -545 -45 -511
rect 45 -545 413 -511
rect 503 -545 871 -511
rect 961 -545 1329 -511
rect 1419 -545 1787 -511
<< metal1 >>
rect -1799 545 -1407 551
rect -1799 511 -1787 545
rect -1419 511 -1407 545
rect -1799 505 -1407 511
rect -1341 545 -949 551
rect -1341 511 -1329 545
rect -961 511 -949 545
rect -1341 505 -949 511
rect -883 545 -491 551
rect -883 511 -871 545
rect -503 511 -491 545
rect -883 505 -491 511
rect -425 545 -33 551
rect -425 511 -413 545
rect -45 511 -33 545
rect -425 505 -33 511
rect 33 545 425 551
rect 33 511 45 545
rect 413 511 425 545
rect 33 505 425 511
rect 491 545 883 551
rect 491 511 503 545
rect 871 511 883 545
rect 491 505 883 511
rect 949 545 1341 551
rect 949 511 961 545
rect 1329 511 1341 545
rect 949 505 1341 511
rect 1407 545 1799 551
rect 1407 511 1419 545
rect 1787 511 1799 545
rect 1407 505 1799 511
rect -1855 452 -1809 464
rect -1855 76 -1849 452
rect -1815 76 -1809 452
rect -1855 64 -1809 76
rect -1397 452 -1351 464
rect -1397 76 -1391 452
rect -1357 76 -1351 452
rect -1397 64 -1351 76
rect -939 452 -893 464
rect -939 76 -933 452
rect -899 76 -893 452
rect -939 64 -893 76
rect -481 452 -435 464
rect -481 76 -475 452
rect -441 76 -435 452
rect -481 64 -435 76
rect -23 452 23 464
rect -23 76 -17 452
rect 17 76 23 452
rect -23 64 23 76
rect 435 452 481 464
rect 435 76 441 452
rect 475 76 481 452
rect 435 64 481 76
rect 893 452 939 464
rect 893 76 899 452
rect 933 76 939 452
rect 893 64 939 76
rect 1351 452 1397 464
rect 1351 76 1357 452
rect 1391 76 1397 452
rect 1351 64 1397 76
rect 1809 452 1855 464
rect 1809 76 1815 452
rect 1849 76 1855 452
rect 1809 64 1855 76
rect -1799 17 -1407 23
rect -1799 -17 -1787 17
rect -1419 -17 -1407 17
rect -1799 -23 -1407 -17
rect -1341 17 -949 23
rect -1341 -17 -1329 17
rect -961 -17 -949 17
rect -1341 -23 -949 -17
rect -883 17 -491 23
rect -883 -17 -871 17
rect -503 -17 -491 17
rect -883 -23 -491 -17
rect -425 17 -33 23
rect -425 -17 -413 17
rect -45 -17 -33 17
rect -425 -23 -33 -17
rect 33 17 425 23
rect 33 -17 45 17
rect 413 -17 425 17
rect 33 -23 425 -17
rect 491 17 883 23
rect 491 -17 503 17
rect 871 -17 883 17
rect 491 -23 883 -17
rect 949 17 1341 23
rect 949 -17 961 17
rect 1329 -17 1341 17
rect 949 -23 1341 -17
rect 1407 17 1799 23
rect 1407 -17 1419 17
rect 1787 -17 1799 17
rect 1407 -23 1799 -17
rect -1855 -76 -1809 -64
rect -1855 -452 -1849 -76
rect -1815 -452 -1809 -76
rect -1855 -464 -1809 -452
rect -1397 -76 -1351 -64
rect -1397 -452 -1391 -76
rect -1357 -452 -1351 -76
rect -1397 -464 -1351 -452
rect -939 -76 -893 -64
rect -939 -452 -933 -76
rect -899 -452 -893 -76
rect -939 -464 -893 -452
rect -481 -76 -435 -64
rect -481 -452 -475 -76
rect -441 -452 -435 -76
rect -481 -464 -435 -452
rect -23 -76 23 -64
rect -23 -452 -17 -76
rect 17 -452 23 -76
rect -23 -464 23 -452
rect 435 -76 481 -64
rect 435 -452 441 -76
rect 475 -452 481 -76
rect 435 -464 481 -452
rect 893 -76 939 -64
rect 893 -452 899 -76
rect 933 -452 939 -76
rect 893 -464 939 -452
rect 1351 -76 1397 -64
rect 1351 -452 1357 -76
rect 1391 -452 1397 -76
rect 1351 -464 1397 -452
rect 1809 -76 1855 -64
rect 1809 -452 1815 -76
rect 1849 -452 1855 -76
rect 1809 -464 1855 -452
rect -1799 -511 -1407 -505
rect -1799 -545 -1787 -511
rect -1419 -545 -1407 -511
rect -1799 -551 -1407 -545
rect -1341 -511 -949 -505
rect -1341 -545 -1329 -511
rect -961 -545 -949 -511
rect -1341 -551 -949 -545
rect -883 -511 -491 -505
rect -883 -545 -871 -511
rect -503 -545 -491 -511
rect -883 -551 -491 -545
rect -425 -511 -33 -505
rect -425 -545 -413 -511
rect -45 -545 -33 -511
rect -425 -551 -33 -545
rect 33 -511 425 -505
rect 33 -545 45 -511
rect 413 -545 425 -511
rect 33 -551 425 -545
rect 491 -511 883 -505
rect 491 -545 503 -511
rect 871 -545 883 -511
rect 491 -551 883 -545
rect 949 -511 1341 -505
rect 949 -545 961 -511
rect 1329 -545 1341 -511
rect 949 -551 1341 -545
rect 1407 -511 1799 -505
rect 1407 -545 1419 -511
rect 1787 -545 1799 -511
rect 1407 -551 1799 -545
<< properties >>
string FIXED_BBOX -1966 -666 1966 666
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 2 m 2 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
