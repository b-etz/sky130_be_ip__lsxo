magic
tech sky130A
magscale 1 2
timestamp 1712250795
<< metal3 >>
rect -8304 1812 -4332 1840
rect -8304 -1812 -4416 1812
rect -4352 -1812 -4332 1812
rect -8304 -1840 -4332 -1812
rect -4092 1812 -120 1840
rect -4092 -1812 -204 1812
rect -140 -1812 -120 1812
rect -4092 -1840 -120 -1812
rect 120 1812 4092 1840
rect 120 -1812 4008 1812
rect 4072 -1812 4092 1812
rect 120 -1840 4092 -1812
rect 4332 1812 8304 1840
rect 4332 -1812 8220 1812
rect 8284 -1812 8304 1812
rect 4332 -1840 8304 -1812
<< via3 >>
rect -4416 -1812 -4352 1812
rect -204 -1812 -140 1812
rect 4008 -1812 4072 1812
rect 8220 -1812 8284 1812
<< mimcap >>
rect -8264 1760 -4664 1800
rect -8264 -1760 -8224 1760
rect -4704 -1760 -4664 1760
rect -8264 -1800 -4664 -1760
rect -4052 1760 -452 1800
rect -4052 -1760 -4012 1760
rect -492 -1760 -452 1760
rect -4052 -1800 -452 -1760
rect 160 1760 3760 1800
rect 160 -1760 200 1760
rect 3720 -1760 3760 1760
rect 160 -1800 3760 -1760
rect 4372 1760 7972 1800
rect 4372 -1760 4412 1760
rect 7932 -1760 7972 1760
rect 4372 -1800 7972 -1760
<< mimcapcontact >>
rect -8224 -1760 -4704 1760
rect -4012 -1760 -492 1760
rect 200 -1760 3720 1760
rect 4412 -1760 7932 1760
<< metal4 >>
rect -4432 1812 -4336 1828
rect -8225 1760 -4703 1761
rect -8225 -1760 -8224 1760
rect -4704 -1760 -4703 1760
rect -8225 -1761 -4703 -1760
rect -4432 -1812 -4416 1812
rect -4352 -1812 -4336 1812
rect -220 1812 -124 1828
rect -4013 1760 -491 1761
rect -4013 -1760 -4012 1760
rect -492 -1760 -491 1760
rect -4013 -1761 -491 -1760
rect -4432 -1828 -4336 -1812
rect -220 -1812 -204 1812
rect -140 -1812 -124 1812
rect 3992 1812 4088 1828
rect 199 1760 3721 1761
rect 199 -1760 200 1760
rect 3720 -1760 3721 1760
rect 199 -1761 3721 -1760
rect -220 -1828 -124 -1812
rect 3992 -1812 4008 1812
rect 4072 -1812 4088 1812
rect 8204 1812 8300 1828
rect 4411 1760 7933 1761
rect 4411 -1760 4412 1760
rect 7932 -1760 7933 1760
rect 4411 -1761 7933 -1760
rect 3992 -1828 4088 -1812
rect 8204 -1812 8220 1812
rect 8284 -1812 8300 1812
rect 8204 -1828 8300 -1812
<< properties >>
string FIXED_BBOX 4332 -1840 8012 1840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 18 l 18 val 661.68 carea 2.00 cperi 0.19 nx 4 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
