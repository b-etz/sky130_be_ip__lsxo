magic
tech sky130A
magscale 1 2
timestamp 1713220443
<< metal3 >>
rect -1986 4040 1700 7720
rect -1986 120 1700 3800
rect -1986 -3800 1700 -120
rect -1986 -7720 1700 -4040
<< mimcap >>
rect -1946 7640 1654 7680
rect -1946 4120 -1906 7640
rect 1614 4120 1654 7640
rect -1946 4080 1654 4120
rect -1946 3720 1654 3760
rect -1946 200 -1906 3720
rect 1614 200 1654 3720
rect -1946 160 1654 200
rect -1946 -200 1654 -160
rect -1946 -3720 -1906 -200
rect 1614 -3720 1654 -200
rect -1946 -3760 1654 -3720
rect -1946 -4120 1654 -4080
rect -1946 -7640 -1906 -4120
rect 1614 -7640 1654 -4120
rect -1946 -7680 1654 -7640
<< mimcapcontact >>
rect -1906 4120 1614 7640
rect -1906 200 1614 3720
rect -1906 -3720 1614 -200
rect -1906 -7640 1614 -4120
<< metal4 >>
rect -198 7641 -94 7724
rect -1907 7640 1615 7641
rect -1907 4120 -1906 7640
rect 1614 4120 1615 7640
rect -1907 4119 1615 4120
rect -198 3721 -94 4119
rect -1907 3720 1615 3721
rect -1907 200 -1906 3720
rect 1614 200 1615 3720
rect -1907 199 1615 200
rect -198 -199 -94 199
rect -1907 -200 1615 -199
rect -1907 -3720 -1906 -200
rect 1614 -3720 1615 -200
rect -1907 -3721 1615 -3720
rect -198 -4119 -94 -3721
rect -1907 -4120 1615 -4119
rect -1907 -7640 -1906 -4120
rect 1614 -7640 1615 -4120
rect -1907 -7641 1615 -7640
rect -198 -7722 -94 -7641
<< properties >>
string FIXED_BBOX -1986 4040 1694 7720
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 18 l 18 val 661.68 carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
