magic
tech sky130A
magscale 1 2
timestamp 1713224120
<< psubdiff >>
rect 472 -1694 532 -1670
rect 472 -1778 532 -1754
<< psubdiffcont >>
rect 472 -1754 532 -1694
<< locali >>
rect 216 -520 798 -506
rect 216 -692 230 -520
rect 402 -556 798 -520
rect 402 -692 416 -556
rect 216 -706 416 -692
rect 758 -776 798 -556
rect 742 -1412 886 -1390
rect 742 -1460 762 -1412
rect 862 -1460 886 -1412
rect 472 -1694 532 -1678
rect 472 -1770 532 -1754
rect 594 -1828 660 -1660
rect 594 -1842 694 -1828
rect 766 -1956 866 -1728
rect 968 -1828 1034 -1660
rect 968 -1842 1068 -1828
rect 1214 -1956 1314 -952
rect 490 -2056 1314 -1956
rect 490 -2068 690 -2056
rect 490 -2400 504 -2068
rect 676 -2400 690 -2068
rect 490 -2416 690 -2400
<< viali >>
rect 230 -692 402 -520
rect 758 -900 796 -812
rect 692 -1014 784 -980
rect 690 -1130 782 -1096
rect 758 -1268 796 -1190
rect 762 -1512 862 -1412
rect 594 -1922 694 -1842
rect 968 -1922 1068 -1842
rect 504 -2400 676 -2068
<< metal1 >>
rect 468 -220 1522 -120
rect 216 -516 416 -506
rect 216 -696 226 -516
rect 406 -696 416 -516
rect 468 -689 564 -220
rect 624 -302 1336 -290
rect 624 -478 636 -302
rect 1324 -478 1336 -302
rect 624 -482 1336 -478
rect 1038 -690 1134 -482
rect 1422 -642 1522 -220
rect 216 -706 416 -696
rect 8690 -738 9016 -642
rect 742 -812 990 -798
rect 742 -904 756 -812
rect 976 -904 990 -812
rect 742 -918 990 -904
rect 678 -964 798 -958
rect 678 -1016 686 -964
rect 792 -1016 798 -964
rect 678 -1022 798 -1016
rect 678 -1090 798 -1084
rect 678 -1142 686 -1090
rect 792 -1142 798 -1090
rect 678 -1148 798 -1142
rect 740 -1190 988 -1184
rect 740 -1198 758 -1190
rect 796 -1198 988 -1190
rect 740 -1290 754 -1198
rect 974 -1290 988 -1198
rect 1086 -1282 1434 -1186
rect 740 -1304 988 -1290
rect 740 -1412 886 -1390
rect 740 -1512 762 -1412
rect 862 -1512 886 -1412
rect 740 -1556 886 -1512
rect 740 -1688 820 -1556
rect 8690 -1674 8700 -794
rect 8842 -1674 8854 -794
rect 740 -1756 746 -1688
rect 814 -1756 820 -1688
rect 8916 -1730 9016 -738
rect 740 -1762 820 -1756
rect 576 -1842 1086 -1826
rect 576 -1922 594 -1842
rect 694 -1922 968 -1842
rect 1068 -1922 1086 -1842
rect 576 -1938 1086 -1922
rect 490 -2068 690 -2056
rect 490 -2400 504 -2068
rect 676 -2400 690 -2068
rect 490 -2416 690 -2400
rect 886 -2106 1086 -1938
rect 1714 -1988 2504 -1976
rect 1714 -2066 1726 -1988
rect 2492 -2066 2504 -1988
rect 1714 -2074 2504 -2066
rect 2606 -2106 2706 -1792
rect 8690 -1826 9016 -1730
rect 886 -2206 1704 -2106
rect 2516 -2206 2706 -2106
rect 886 -2416 1086 -2206
<< via1 >>
rect 226 -520 406 -516
rect 226 -692 230 -520
rect 230 -692 402 -520
rect 402 -692 406 -520
rect 226 -696 406 -692
rect 636 -478 1324 -302
rect 756 -900 758 -812
rect 758 -900 796 -812
rect 796 -900 976 -812
rect 756 -904 976 -900
rect 686 -980 792 -964
rect 686 -1014 692 -980
rect 692 -1014 784 -980
rect 784 -1014 792 -980
rect 686 -1016 792 -1014
rect 686 -1096 792 -1090
rect 686 -1130 690 -1096
rect 690 -1130 782 -1096
rect 782 -1130 792 -1096
rect 686 -1142 792 -1130
rect 754 -1268 758 -1198
rect 758 -1268 796 -1198
rect 796 -1268 974 -1198
rect 754 -1290 974 -1268
rect 8700 -1674 8842 -794
rect 746 -1756 814 -1688
rect 1726 -2066 2492 -1988
<< metal2 >>
rect 624 -302 1336 -290
rect 624 -478 636 -302
rect 1324 -478 1336 -302
rect 624 -482 1336 -478
rect 216 -516 416 -506
rect 216 -696 226 -516
rect 406 -696 416 -516
rect 216 -706 416 -696
rect 910 -642 1798 -542
rect 910 -798 990 -642
rect 742 -812 990 -798
rect 216 -950 416 -830
rect 742 -904 756 -812
rect 976 -904 990 -812
rect 742 -918 990 -904
rect 1280 -950 1360 -868
rect 1698 -912 1798 -642
rect 216 -964 1360 -950
rect 216 -1016 686 -964
rect 792 -1016 1360 -964
rect 216 -1030 1360 -1016
rect 216 -1090 1360 -1076
rect 216 -1142 686 -1090
rect 792 -1142 1360 -1090
rect 216 -1156 1360 -1142
rect 216 -1276 416 -1156
rect 740 -1198 988 -1184
rect 740 -1290 754 -1198
rect 974 -1290 988 -1198
rect 740 -1304 988 -1290
rect 740 -1688 820 -1682
rect 740 -1756 746 -1688
rect 814 -1756 820 -1688
rect 740 -1978 820 -1756
rect 908 -1826 988 -1304
rect 1280 -1608 1360 -1156
rect 1698 -1826 1798 -1556
rect 8690 -1674 8700 -794
rect 8842 -1674 8854 -794
rect 908 -1926 1798 -1826
rect 740 -1988 2504 -1978
rect 740 -2038 1726 -1988
rect 1714 -2066 1726 -2038
rect 2492 -2066 2504 -1988
rect 1714 -2074 2504 -2066
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1713224120
transform 0 1 542 -1 0 -598
box -38 -48 130 592
use ripple_dly_4  x1
timestamp 1713224120
transform 1 0 1378 0 -1 -1870
box -98 -1228 7350 -588
use ripple_dly_4  x2
timestamp 1713224120
transform 1 0 1378 0 1 -598
box -98 -1228 7350 -588
use sky130_fd_sc_hd__a221o_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1713224120
transform 0 1 542 -1 0 -690
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_0  x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1713224120
transform 0 1 542 -1 0 -1426
box -38 -48 406 592
use sky130_fd_pr__nfet_01v8_AHZR5K  XM3
timestamp 1713224120
transform 1 0 2110 0 1 -2156
box -596 -260 596 260
<< labels >>
flabel space 624 -490 1336 -290 0 FreeSans 800 0 0 0 dvdd
port 1 nsew
flabel metal1 490 -2416 690 -2056 0 FreeSans 800 0 0 0 clkin
port 3 nsew
flabel metal1 886 -2416 1086 -2206 0 FreeSans 800 0 0 0 clkout
port 4 nsew
flabel metal2 216 -1030 416 -830 0 FreeSans 800 0 0 0 ena
port 5 nsew
flabel metal2 216 -706 416 -506 0 FreeSans 800 0 0 0 stby
port 6 nsew
flabel metal2 216 -1276 416 -1076 0 FreeSans 800 0 0 0 stby_b
port 7 nsew
flabel metal2 740 -2038 1726 -1978 0 FreeSans 400 0 0 0 clk_disable
flabel metal1 494 -220 1470 -120 0 FreeSans 800 0 0 0 dvss
port 2 nsew
flabel metal2 910 -642 1798 -542 0 FreeSans 400 0 0 0 ena_done_b
flabel metal2 908 -1926 1798 -1826 0 FreeSans 400 0 0 0 stby_done_b
<< end >>
