magic
tech sky130A
magscale 1 2
timestamp 1712851378
<< pwell >>
rect -367 -15582 367 15582
<< psubdiff >>
rect -331 15512 -235 15546
rect 235 15512 331 15546
rect -331 15450 -297 15512
rect 297 15450 331 15512
rect -331 -15512 -297 -15450
rect 297 -15512 331 -15450
rect -331 -15546 -235 -15512
rect 235 -15546 331 -15512
<< psubdiffcont >>
rect -235 15512 235 15546
rect -331 -15450 -297 15450
rect 297 -15450 331 15450
rect -235 -15546 235 -15512
<< xpolycontact >>
rect -201 14984 -131 15416
rect -201 -15416 -131 -14984
rect -35 14984 35 15416
rect -35 -15416 35 -14984
rect 131 14984 201 15416
rect 131 -15416 201 -14984
<< xpolyres >>
rect -201 -14984 -131 14984
rect -35 -14984 35 14984
rect 131 -14984 201 14984
<< locali >>
rect -331 15512 -235 15546
rect 235 15512 331 15546
rect -331 15450 -297 15512
rect 297 15450 331 15512
rect -331 -15512 -297 -15450
rect 297 -15512 331 -15450
rect -331 -15546 -235 -15512
rect 235 -15546 331 -15512
<< viali >>
rect -185 15001 -147 15398
rect -19 15001 19 15398
rect 147 15001 185 15398
rect -185 -15398 -147 -15001
rect -19 -15398 19 -15001
rect 147 -15398 185 -15001
<< metal1 >>
rect -191 15398 -141 15410
rect -191 15001 -185 15398
rect -147 15001 -141 15398
rect -191 14989 -141 15001
rect -25 15398 25 15410
rect -25 15001 -19 15398
rect 19 15001 25 15398
rect -25 14989 25 15001
rect 141 15398 191 15410
rect 141 15001 147 15398
rect 185 15001 191 15398
rect 141 14989 191 15001
rect -191 -15001 -141 -14989
rect -191 -15398 -185 -15001
rect -147 -15398 -141 -15001
rect -191 -15410 -141 -15398
rect -25 -15001 25 -14989
rect -25 -15398 -19 -15001
rect 19 -15398 25 -15001
rect -25 -15410 25 -15398
rect 141 -15001 191 -14989
rect 141 -15398 147 -15001
rect 185 -15398 191 -15001
rect 141 -15410 191 -15398
<< properties >>
string FIXED_BBOX -314 -15529 314 15529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 150 m 1 nx 3 wmin 0.350 lmin 0.50 rho 2000 val 858.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
