magic
tech sky130A
magscale 1 2
timestamp 1712087189
<< nwell >>
rect -562 -1137 562 1137
<< pmos >>
rect -366 118 -266 918
rect -208 118 -108 918
rect -50 118 50 918
rect 108 118 208 918
rect 266 118 366 918
rect -366 -918 -266 -118
rect -208 -918 -108 -118
rect -50 -918 50 -118
rect 108 -918 208 -118
rect 266 -918 366 -118
<< pdiff >>
rect -424 906 -366 918
rect -424 130 -412 906
rect -378 130 -366 906
rect -424 118 -366 130
rect -266 906 -208 918
rect -266 130 -254 906
rect -220 130 -208 906
rect -266 118 -208 130
rect -108 906 -50 918
rect -108 130 -96 906
rect -62 130 -50 906
rect -108 118 -50 130
rect 50 906 108 918
rect 50 130 62 906
rect 96 130 108 906
rect 50 118 108 130
rect 208 906 266 918
rect 208 130 220 906
rect 254 130 266 906
rect 208 118 266 130
rect 366 906 424 918
rect 366 130 378 906
rect 412 130 424 906
rect 366 118 424 130
rect -424 -130 -366 -118
rect -424 -906 -412 -130
rect -378 -906 -366 -130
rect -424 -918 -366 -906
rect -266 -130 -208 -118
rect -266 -906 -254 -130
rect -220 -906 -208 -130
rect -266 -918 -208 -906
rect -108 -130 -50 -118
rect -108 -906 -96 -130
rect -62 -906 -50 -130
rect -108 -918 -50 -906
rect 50 -130 108 -118
rect 50 -906 62 -130
rect 96 -906 108 -130
rect 50 -918 108 -906
rect 208 -130 266 -118
rect 208 -906 220 -130
rect 254 -906 266 -130
rect 208 -918 266 -906
rect 366 -130 424 -118
rect 366 -906 378 -130
rect 412 -906 424 -130
rect 366 -918 424 -906
<< pdiffc >>
rect -412 130 -378 906
rect -254 130 -220 906
rect -96 130 -62 906
rect 62 130 96 906
rect 220 130 254 906
rect 378 130 412 906
rect -412 -906 -378 -130
rect -254 -906 -220 -130
rect -96 -906 -62 -130
rect 62 -906 96 -130
rect 220 -906 254 -130
rect 378 -906 412 -130
<< nsubdiff >>
rect -526 1067 -430 1101
rect 430 1067 526 1101
rect -526 1005 -492 1067
rect 492 1005 526 1067
rect -526 -1067 -492 -1005
rect 492 -1067 526 -1005
rect -526 -1101 -430 -1067
rect 430 -1101 526 -1067
<< nsubdiffcont >>
rect -430 1067 430 1101
rect -526 -1005 -492 1005
rect 492 -1005 526 1005
rect -430 -1101 430 -1067
<< poly >>
rect -366 999 -266 1015
rect -366 965 -350 999
rect -282 965 -266 999
rect -366 918 -266 965
rect -208 999 -108 1015
rect -208 965 -192 999
rect -124 965 -108 999
rect -208 918 -108 965
rect -50 999 50 1015
rect -50 965 -34 999
rect 34 965 50 999
rect -50 918 50 965
rect 108 999 208 1015
rect 108 965 124 999
rect 192 965 208 999
rect 108 918 208 965
rect 266 999 366 1015
rect 266 965 282 999
rect 350 965 366 999
rect 266 918 366 965
rect -366 71 -266 118
rect -366 37 -350 71
rect -282 37 -266 71
rect -366 21 -266 37
rect -208 71 -108 118
rect -208 37 -192 71
rect -124 37 -108 71
rect -208 21 -108 37
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect 108 71 208 118
rect 108 37 124 71
rect 192 37 208 71
rect 108 21 208 37
rect 266 71 366 118
rect 266 37 282 71
rect 350 37 366 71
rect 266 21 366 37
rect -366 -37 -266 -21
rect -366 -71 -350 -37
rect -282 -71 -266 -37
rect -366 -118 -266 -71
rect -208 -37 -108 -21
rect -208 -71 -192 -37
rect -124 -71 -108 -37
rect -208 -118 -108 -71
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect 108 -37 208 -21
rect 108 -71 124 -37
rect 192 -71 208 -37
rect 108 -118 208 -71
rect 266 -37 366 -21
rect 266 -71 282 -37
rect 350 -71 366 -37
rect 266 -118 366 -71
rect -366 -965 -266 -918
rect -366 -999 -350 -965
rect -282 -999 -266 -965
rect -366 -1015 -266 -999
rect -208 -965 -108 -918
rect -208 -999 -192 -965
rect -124 -999 -108 -965
rect -208 -1015 -108 -999
rect -50 -965 50 -918
rect -50 -999 -34 -965
rect 34 -999 50 -965
rect -50 -1015 50 -999
rect 108 -965 208 -918
rect 108 -999 124 -965
rect 192 -999 208 -965
rect 108 -1015 208 -999
rect 266 -965 366 -918
rect 266 -999 282 -965
rect 350 -999 366 -965
rect 266 -1015 366 -999
<< polycont >>
rect -350 965 -282 999
rect -192 965 -124 999
rect -34 965 34 999
rect 124 965 192 999
rect 282 965 350 999
rect -350 37 -282 71
rect -192 37 -124 71
rect -34 37 34 71
rect 124 37 192 71
rect 282 37 350 71
rect -350 -71 -282 -37
rect -192 -71 -124 -37
rect -34 -71 34 -37
rect 124 -71 192 -37
rect 282 -71 350 -37
rect -350 -999 -282 -965
rect -192 -999 -124 -965
rect -34 -999 34 -965
rect 124 -999 192 -965
rect 282 -999 350 -965
<< locali >>
rect -526 1067 -430 1101
rect 430 1067 526 1101
rect -526 1005 -492 1067
rect 492 1005 526 1067
rect -366 965 -350 999
rect -282 965 -266 999
rect -208 965 -192 999
rect -124 965 -108 999
rect -50 965 -34 999
rect 34 965 50 999
rect 108 965 124 999
rect 192 965 208 999
rect 266 965 282 999
rect 350 965 366 999
rect -412 906 -378 922
rect -412 114 -378 130
rect -254 906 -220 922
rect -254 114 -220 130
rect -96 906 -62 922
rect -96 114 -62 130
rect 62 906 96 922
rect 62 114 96 130
rect 220 906 254 922
rect 220 114 254 130
rect 378 906 412 922
rect 378 114 412 130
rect -366 37 -350 71
rect -282 37 -266 71
rect -208 37 -192 71
rect -124 37 -108 71
rect -50 37 -34 71
rect 34 37 50 71
rect 108 37 124 71
rect 192 37 208 71
rect 266 37 282 71
rect 350 37 366 71
rect -366 -71 -350 -37
rect -282 -71 -266 -37
rect -208 -71 -192 -37
rect -124 -71 -108 -37
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect 108 -71 124 -37
rect 192 -71 208 -37
rect 266 -71 282 -37
rect 350 -71 366 -37
rect -412 -130 -378 -114
rect -412 -922 -378 -906
rect -254 -130 -220 -114
rect -254 -922 -220 -906
rect -96 -130 -62 -114
rect -96 -922 -62 -906
rect 62 -130 96 -114
rect 62 -922 96 -906
rect 220 -130 254 -114
rect 220 -922 254 -906
rect 378 -130 412 -114
rect 378 -922 412 -906
rect -366 -999 -350 -965
rect -282 -999 -266 -965
rect -208 -999 -192 -965
rect -124 -999 -108 -965
rect -50 -999 -34 -965
rect 34 -999 50 -965
rect 108 -999 124 -965
rect 192 -999 208 -965
rect 266 -999 282 -965
rect 350 -999 366 -965
rect -526 -1067 -492 -1005
rect 492 -1067 526 -1005
rect -526 -1101 -430 -1067
rect 430 -1101 526 -1067
<< viali >>
rect -350 965 -282 999
rect -192 965 -124 999
rect -34 965 34 999
rect 124 965 192 999
rect 282 965 350 999
rect -412 130 -378 906
rect -254 130 -220 906
rect -96 130 -62 906
rect 62 130 96 906
rect 220 130 254 906
rect 378 130 412 906
rect -350 37 -282 71
rect -192 37 -124 71
rect -34 37 34 71
rect 124 37 192 71
rect 282 37 350 71
rect -350 -71 -282 -37
rect -192 -71 -124 -37
rect -34 -71 34 -37
rect 124 -71 192 -37
rect 282 -71 350 -37
rect -412 -906 -378 -130
rect -254 -906 -220 -130
rect -96 -906 -62 -130
rect 62 -906 96 -130
rect 220 -906 254 -130
rect 378 -906 412 -130
rect -350 -999 -282 -965
rect -192 -999 -124 -965
rect -34 -999 34 -965
rect 124 -999 192 -965
rect 282 -999 350 -965
<< metal1 >>
rect -362 999 -270 1005
rect -362 965 -350 999
rect -282 965 -270 999
rect -362 959 -270 965
rect -204 999 -112 1005
rect -204 965 -192 999
rect -124 965 -112 999
rect -204 959 -112 965
rect -46 999 46 1005
rect -46 965 -34 999
rect 34 965 46 999
rect -46 959 46 965
rect 112 999 204 1005
rect 112 965 124 999
rect 192 965 204 999
rect 112 959 204 965
rect 270 999 362 1005
rect 270 965 282 999
rect 350 965 362 999
rect 270 959 362 965
rect -418 906 -372 918
rect -418 130 -412 906
rect -378 130 -372 906
rect -418 118 -372 130
rect -260 906 -214 918
rect -260 130 -254 906
rect -220 130 -214 906
rect -260 118 -214 130
rect -102 906 -56 918
rect -102 130 -96 906
rect -62 130 -56 906
rect -102 118 -56 130
rect 56 906 102 918
rect 56 130 62 906
rect 96 130 102 906
rect 56 118 102 130
rect 214 906 260 918
rect 214 130 220 906
rect 254 130 260 906
rect 214 118 260 130
rect 372 906 418 918
rect 372 130 378 906
rect 412 130 418 906
rect 372 118 418 130
rect -362 71 -270 77
rect -362 37 -350 71
rect -282 37 -270 71
rect -362 31 -270 37
rect -204 71 -112 77
rect -204 37 -192 71
rect -124 37 -112 71
rect -204 31 -112 37
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect 112 71 204 77
rect 112 37 124 71
rect 192 37 204 71
rect 112 31 204 37
rect 270 71 362 77
rect 270 37 282 71
rect 350 37 362 71
rect 270 31 362 37
rect -362 -37 -270 -31
rect -362 -71 -350 -37
rect -282 -71 -270 -37
rect -362 -77 -270 -71
rect -204 -37 -112 -31
rect -204 -71 -192 -37
rect -124 -71 -112 -37
rect -204 -77 -112 -71
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect 112 -37 204 -31
rect 112 -71 124 -37
rect 192 -71 204 -37
rect 112 -77 204 -71
rect 270 -37 362 -31
rect 270 -71 282 -37
rect 350 -71 362 -37
rect 270 -77 362 -71
rect -418 -130 -372 -118
rect -418 -906 -412 -130
rect -378 -906 -372 -130
rect -418 -918 -372 -906
rect -260 -130 -214 -118
rect -260 -906 -254 -130
rect -220 -906 -214 -130
rect -260 -918 -214 -906
rect -102 -130 -56 -118
rect -102 -906 -96 -130
rect -62 -906 -56 -130
rect -102 -918 -56 -906
rect 56 -130 102 -118
rect 56 -906 62 -130
rect 96 -906 102 -130
rect 56 -918 102 -906
rect 214 -130 260 -118
rect 214 -906 220 -130
rect 254 -906 260 -130
rect 214 -918 260 -906
rect 372 -130 418 -118
rect 372 -906 378 -130
rect 412 -906 418 -130
rect 372 -918 418 -906
rect -362 -965 -270 -959
rect -362 -999 -350 -965
rect -282 -999 -270 -965
rect -362 -1005 -270 -999
rect -204 -965 -112 -959
rect -204 -999 -192 -965
rect -124 -999 -112 -965
rect -204 -1005 -112 -999
rect -46 -965 46 -959
rect -46 -999 -34 -965
rect 34 -999 46 -965
rect -46 -1005 46 -999
rect 112 -965 204 -959
rect 112 -999 124 -965
rect 192 -999 204 -965
rect 112 -1005 204 -999
rect 270 -965 362 -959
rect 270 -999 282 -965
rect 350 -999 362 -965
rect 270 -1005 362 -999
<< properties >>
string FIXED_BBOX -509 -1084 509 1084
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.0 l 0.5 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
