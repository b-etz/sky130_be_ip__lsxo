magic
tech sky130A
magscale 1 2
timestamp 1712073863
<< metal3 >>
rect -4092 3772 -120 3800
rect -4092 148 -204 3772
rect -140 148 -120 3772
rect -4092 120 -120 148
rect 120 3772 4092 3800
rect 120 148 4008 3772
rect 4072 148 4092 3772
rect 120 120 4092 148
rect -4092 -148 -120 -120
rect -4092 -3772 -204 -148
rect -140 -3772 -120 -148
rect -4092 -3800 -120 -3772
rect 120 -148 4092 -120
rect 120 -3772 4008 -148
rect 4072 -3772 4092 -148
rect 120 -3800 4092 -3772
<< via3 >>
rect -204 148 -140 3772
rect 4008 148 4072 3772
rect -204 -3772 -140 -148
rect 4008 -3772 4072 -148
<< mimcap >>
rect -4052 3720 -452 3760
rect -4052 200 -4012 3720
rect -492 200 -452 3720
rect -4052 160 -452 200
rect 160 3720 3760 3760
rect 160 200 200 3720
rect 3720 200 3760 3720
rect 160 160 3760 200
rect -4052 -200 -452 -160
rect -4052 -3720 -4012 -200
rect -492 -3720 -452 -200
rect -4052 -3760 -452 -3720
rect 160 -200 3760 -160
rect 160 -3720 200 -200
rect 3720 -3720 3760 -200
rect 160 -3760 3760 -3720
<< mimcapcontact >>
rect -4012 200 -492 3720
rect 200 200 3720 3720
rect -4012 -3720 -492 -200
rect 200 -3720 3720 -200
<< metal4 >>
rect -2304 3721 -2200 3920
rect -224 3772 -120 3920
rect -4013 3720 -491 3721
rect -4013 200 -4012 3720
rect -492 200 -491 3720
rect -4013 199 -491 200
rect -2304 -199 -2200 199
rect -224 148 -204 3772
rect -140 148 -120 3772
rect 1908 3721 2012 3920
rect 3988 3772 4092 3920
rect 199 3720 3721 3721
rect 199 200 200 3720
rect 3720 200 3721 3720
rect 199 199 3721 200
rect -224 -148 -120 148
rect -4013 -200 -491 -199
rect -4013 -3720 -4012 -200
rect -492 -3720 -491 -200
rect -4013 -3721 -491 -3720
rect -2304 -3920 -2200 -3721
rect -224 -3772 -204 -148
rect -140 -3772 -120 -148
rect 1908 -199 2012 199
rect 3988 148 4008 3772
rect 4072 148 4092 3772
rect 3988 -148 4092 148
rect 199 -200 3721 -199
rect 199 -3720 200 -200
rect 3720 -3720 3721 -200
rect 199 -3721 3721 -3720
rect -224 -3920 -120 -3772
rect 1908 -3920 2012 -3721
rect 3988 -3772 4008 -148
rect 4072 -3772 4092 -148
rect 3988 -3920 4092 -3772
<< properties >>
string FIXED_BBOX 120 120 3800 3800
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 18 l 18 val 661.68 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
