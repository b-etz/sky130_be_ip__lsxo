magic
tech sky130A
magscale 1 2
timestamp 1712848480
<< metal3 >>
rect -3798 9132 -1426 9160
rect -3798 7108 -1510 9132
rect -1446 7108 -1426 9132
rect -3798 7080 -1426 7108
rect -1186 9132 1186 9160
rect -1186 7108 1102 9132
rect 1166 7108 1186 9132
rect -1186 7080 1186 7108
rect 1426 9132 3798 9160
rect 1426 7108 3714 9132
rect 3778 7108 3798 9132
rect 1426 7080 3798 7108
rect -3798 6812 -1426 6840
rect -3798 4788 -1510 6812
rect -1446 4788 -1426 6812
rect -3798 4760 -1426 4788
rect -1186 6812 1186 6840
rect -1186 4788 1102 6812
rect 1166 4788 1186 6812
rect -1186 4760 1186 4788
rect 1426 6812 3798 6840
rect 1426 4788 3714 6812
rect 3778 4788 3798 6812
rect 1426 4760 3798 4788
rect -3798 4492 -1426 4520
rect -3798 2468 -1510 4492
rect -1446 2468 -1426 4492
rect -3798 2440 -1426 2468
rect -1186 4492 1186 4520
rect -1186 2468 1102 4492
rect 1166 2468 1186 4492
rect -1186 2440 1186 2468
rect 1426 4492 3798 4520
rect 1426 2468 3714 4492
rect 3778 2468 3798 4492
rect 1426 2440 3798 2468
rect -3798 2172 -1426 2200
rect -3798 148 -1510 2172
rect -1446 148 -1426 2172
rect -3798 120 -1426 148
rect -1186 2172 1186 2200
rect -1186 148 1102 2172
rect 1166 148 1186 2172
rect -1186 120 1186 148
rect 1426 2172 3798 2200
rect 1426 148 3714 2172
rect 3778 148 3798 2172
rect 1426 120 3798 148
rect -3798 -148 -1426 -120
rect -3798 -2172 -1510 -148
rect -1446 -2172 -1426 -148
rect -3798 -2200 -1426 -2172
rect -1186 -148 1186 -120
rect -1186 -2172 1102 -148
rect 1166 -2172 1186 -148
rect -1186 -2200 1186 -2172
rect 1426 -148 3798 -120
rect 1426 -2172 3714 -148
rect 3778 -2172 3798 -148
rect 1426 -2200 3798 -2172
rect -3798 -2468 -1426 -2440
rect -3798 -4492 -1510 -2468
rect -1446 -4492 -1426 -2468
rect -3798 -4520 -1426 -4492
rect -1186 -2468 1186 -2440
rect -1186 -4492 1102 -2468
rect 1166 -4492 1186 -2468
rect -1186 -4520 1186 -4492
rect 1426 -2468 3798 -2440
rect 1426 -4492 3714 -2468
rect 3778 -4492 3798 -2468
rect 1426 -4520 3798 -4492
rect -3798 -4788 -1426 -4760
rect -3798 -6812 -1510 -4788
rect -1446 -6812 -1426 -4788
rect -3798 -6840 -1426 -6812
rect -1186 -4788 1186 -4760
rect -1186 -6812 1102 -4788
rect 1166 -6812 1186 -4788
rect -1186 -6840 1186 -6812
rect 1426 -4788 3798 -4760
rect 1426 -6812 3714 -4788
rect 3778 -6812 3798 -4788
rect 1426 -6840 3798 -6812
rect -3798 -7108 -1426 -7080
rect -3798 -9132 -1510 -7108
rect -1446 -9132 -1426 -7108
rect -3798 -9160 -1426 -9132
rect -1186 -7108 1186 -7080
rect -1186 -9132 1102 -7108
rect 1166 -9132 1186 -7108
rect -1186 -9160 1186 -9132
rect 1426 -7108 3798 -7080
rect 1426 -9132 3714 -7108
rect 3778 -9132 3798 -7108
rect 1426 -9160 3798 -9132
<< via3 >>
rect -1510 7108 -1446 9132
rect 1102 7108 1166 9132
rect 3714 7108 3778 9132
rect -1510 4788 -1446 6812
rect 1102 4788 1166 6812
rect 3714 4788 3778 6812
rect -1510 2468 -1446 4492
rect 1102 2468 1166 4492
rect 3714 2468 3778 4492
rect -1510 148 -1446 2172
rect 1102 148 1166 2172
rect 3714 148 3778 2172
rect -1510 -2172 -1446 -148
rect 1102 -2172 1166 -148
rect 3714 -2172 3778 -148
rect -1510 -4492 -1446 -2468
rect 1102 -4492 1166 -2468
rect 3714 -4492 3778 -2468
rect -1510 -6812 -1446 -4788
rect 1102 -6812 1166 -4788
rect 3714 -6812 3778 -4788
rect -1510 -9132 -1446 -7108
rect 1102 -9132 1166 -7108
rect 3714 -9132 3778 -7108
<< mimcap >>
rect -3758 9080 -1758 9120
rect -3758 7160 -3718 9080
rect -1798 7160 -1758 9080
rect -3758 7120 -1758 7160
rect -1146 9080 854 9120
rect -1146 7160 -1106 9080
rect 814 7160 854 9080
rect -1146 7120 854 7160
rect 1466 9080 3466 9120
rect 1466 7160 1506 9080
rect 3426 7160 3466 9080
rect 1466 7120 3466 7160
rect -3758 6760 -1758 6800
rect -3758 4840 -3718 6760
rect -1798 4840 -1758 6760
rect -3758 4800 -1758 4840
rect -1146 6760 854 6800
rect -1146 4840 -1106 6760
rect 814 4840 854 6760
rect -1146 4800 854 4840
rect 1466 6760 3466 6800
rect 1466 4840 1506 6760
rect 3426 4840 3466 6760
rect 1466 4800 3466 4840
rect -3758 4440 -1758 4480
rect -3758 2520 -3718 4440
rect -1798 2520 -1758 4440
rect -3758 2480 -1758 2520
rect -1146 4440 854 4480
rect -1146 2520 -1106 4440
rect 814 2520 854 4440
rect -1146 2480 854 2520
rect 1466 4440 3466 4480
rect 1466 2520 1506 4440
rect 3426 2520 3466 4440
rect 1466 2480 3466 2520
rect -3758 2120 -1758 2160
rect -3758 200 -3718 2120
rect -1798 200 -1758 2120
rect -3758 160 -1758 200
rect -1146 2120 854 2160
rect -1146 200 -1106 2120
rect 814 200 854 2120
rect -1146 160 854 200
rect 1466 2120 3466 2160
rect 1466 200 1506 2120
rect 3426 200 3466 2120
rect 1466 160 3466 200
rect -3758 -200 -1758 -160
rect -3758 -2120 -3718 -200
rect -1798 -2120 -1758 -200
rect -3758 -2160 -1758 -2120
rect -1146 -200 854 -160
rect -1146 -2120 -1106 -200
rect 814 -2120 854 -200
rect -1146 -2160 854 -2120
rect 1466 -200 3466 -160
rect 1466 -2120 1506 -200
rect 3426 -2120 3466 -200
rect 1466 -2160 3466 -2120
rect -3758 -2520 -1758 -2480
rect -3758 -4440 -3718 -2520
rect -1798 -4440 -1758 -2520
rect -3758 -4480 -1758 -4440
rect -1146 -2520 854 -2480
rect -1146 -4440 -1106 -2520
rect 814 -4440 854 -2520
rect -1146 -4480 854 -4440
rect 1466 -2520 3466 -2480
rect 1466 -4440 1506 -2520
rect 3426 -4440 3466 -2520
rect 1466 -4480 3466 -4440
rect -3758 -4840 -1758 -4800
rect -3758 -6760 -3718 -4840
rect -1798 -6760 -1758 -4840
rect -3758 -6800 -1758 -6760
rect -1146 -4840 854 -4800
rect -1146 -6760 -1106 -4840
rect 814 -6760 854 -4840
rect -1146 -6800 854 -6760
rect 1466 -4840 3466 -4800
rect 1466 -6760 1506 -4840
rect 3426 -6760 3466 -4840
rect 1466 -6800 3466 -6760
rect -3758 -7160 -1758 -7120
rect -3758 -9080 -3718 -7160
rect -1798 -9080 -1758 -7160
rect -3758 -9120 -1758 -9080
rect -1146 -7160 854 -7120
rect -1146 -9080 -1106 -7160
rect 814 -9080 854 -7160
rect -1146 -9120 854 -9080
rect 1466 -7160 3466 -7120
rect 1466 -9080 1506 -7160
rect 3426 -9080 3466 -7160
rect 1466 -9120 3466 -9080
<< mimcapcontact >>
rect -3718 7160 -1798 9080
rect -1106 7160 814 9080
rect 1506 7160 3426 9080
rect -3718 4840 -1798 6760
rect -1106 4840 814 6760
rect 1506 4840 3426 6760
rect -3718 2520 -1798 4440
rect -1106 2520 814 4440
rect 1506 2520 3426 4440
rect -3718 200 -1798 2120
rect -1106 200 814 2120
rect 1506 200 3426 2120
rect -3718 -2120 -1798 -200
rect -1106 -2120 814 -200
rect 1506 -2120 3426 -200
rect -3718 -4440 -1798 -2520
rect -1106 -4440 814 -2520
rect 1506 -4440 3426 -2520
rect -3718 -6760 -1798 -4840
rect -1106 -6760 814 -4840
rect 1506 -6760 3426 -4840
rect -3718 -9080 -1798 -7160
rect -1106 -9080 814 -7160
rect 1506 -9080 3426 -7160
<< metal4 >>
rect -2810 9081 -2706 9280
rect -1530 9132 -1426 9280
rect -3719 9080 -1797 9081
rect -3719 7160 -3718 9080
rect -1798 7160 -1797 9080
rect -3719 7159 -1797 7160
rect -2810 6761 -2706 7159
rect -1530 7108 -1510 9132
rect -1446 7108 -1426 9132
rect -198 9081 -94 9280
rect 1082 9132 1186 9280
rect -1107 9080 815 9081
rect -1107 7160 -1106 9080
rect 814 7160 815 9080
rect -1107 7159 815 7160
rect -1530 6812 -1426 7108
rect -3719 6760 -1797 6761
rect -3719 4840 -3718 6760
rect -1798 4840 -1797 6760
rect -3719 4839 -1797 4840
rect -2810 4441 -2706 4839
rect -1530 4788 -1510 6812
rect -1446 4788 -1426 6812
rect -198 6761 -94 7159
rect 1082 7108 1102 9132
rect 1166 7108 1186 9132
rect 2414 9081 2518 9280
rect 3694 9132 3798 9280
rect 1505 9080 3427 9081
rect 1505 7160 1506 9080
rect 3426 7160 3427 9080
rect 1505 7159 3427 7160
rect 1082 6812 1186 7108
rect -1107 6760 815 6761
rect -1107 4840 -1106 6760
rect 814 4840 815 6760
rect -1107 4839 815 4840
rect -1530 4492 -1426 4788
rect -3719 4440 -1797 4441
rect -3719 2520 -3718 4440
rect -1798 2520 -1797 4440
rect -3719 2519 -1797 2520
rect -2810 2121 -2706 2519
rect -1530 2468 -1510 4492
rect -1446 2468 -1426 4492
rect -198 4441 -94 4839
rect 1082 4788 1102 6812
rect 1166 4788 1186 6812
rect 2414 6761 2518 7159
rect 3694 7108 3714 9132
rect 3778 7108 3798 9132
rect 3694 6812 3798 7108
rect 1505 6760 3427 6761
rect 1505 4840 1506 6760
rect 3426 4840 3427 6760
rect 1505 4839 3427 4840
rect 1082 4492 1186 4788
rect -1107 4440 815 4441
rect -1107 2520 -1106 4440
rect 814 2520 815 4440
rect -1107 2519 815 2520
rect -1530 2172 -1426 2468
rect -3719 2120 -1797 2121
rect -3719 200 -3718 2120
rect -1798 200 -1797 2120
rect -3719 199 -1797 200
rect -2810 -199 -2706 199
rect -1530 148 -1510 2172
rect -1446 148 -1426 2172
rect -198 2121 -94 2519
rect 1082 2468 1102 4492
rect 1166 2468 1186 4492
rect 2414 4441 2518 4839
rect 3694 4788 3714 6812
rect 3778 4788 3798 6812
rect 3694 4492 3798 4788
rect 1505 4440 3427 4441
rect 1505 2520 1506 4440
rect 3426 2520 3427 4440
rect 1505 2519 3427 2520
rect 1082 2172 1186 2468
rect -1107 2120 815 2121
rect -1107 200 -1106 2120
rect 814 200 815 2120
rect -1107 199 815 200
rect -1530 -148 -1426 148
rect -3719 -200 -1797 -199
rect -3719 -2120 -3718 -200
rect -1798 -2120 -1797 -200
rect -3719 -2121 -1797 -2120
rect -2810 -2519 -2706 -2121
rect -1530 -2172 -1510 -148
rect -1446 -2172 -1426 -148
rect -198 -199 -94 199
rect 1082 148 1102 2172
rect 1166 148 1186 2172
rect 2414 2121 2518 2519
rect 3694 2468 3714 4492
rect 3778 2468 3798 4492
rect 3694 2172 3798 2468
rect 1505 2120 3427 2121
rect 1505 200 1506 2120
rect 3426 200 3427 2120
rect 1505 199 3427 200
rect 1082 -148 1186 148
rect -1107 -200 815 -199
rect -1107 -2120 -1106 -200
rect 814 -2120 815 -200
rect -1107 -2121 815 -2120
rect -1530 -2468 -1426 -2172
rect -3719 -2520 -1797 -2519
rect -3719 -4440 -3718 -2520
rect -1798 -4440 -1797 -2520
rect -3719 -4441 -1797 -4440
rect -2810 -4839 -2706 -4441
rect -1530 -4492 -1510 -2468
rect -1446 -4492 -1426 -2468
rect -198 -2519 -94 -2121
rect 1082 -2172 1102 -148
rect 1166 -2172 1186 -148
rect 2414 -199 2518 199
rect 3694 148 3714 2172
rect 3778 148 3798 2172
rect 3694 -148 3798 148
rect 1505 -200 3427 -199
rect 1505 -2120 1506 -200
rect 3426 -2120 3427 -200
rect 1505 -2121 3427 -2120
rect 1082 -2468 1186 -2172
rect -1107 -2520 815 -2519
rect -1107 -4440 -1106 -2520
rect 814 -4440 815 -2520
rect -1107 -4441 815 -4440
rect -1530 -4788 -1426 -4492
rect -3719 -4840 -1797 -4839
rect -3719 -6760 -3718 -4840
rect -1798 -6760 -1797 -4840
rect -3719 -6761 -1797 -6760
rect -2810 -7159 -2706 -6761
rect -1530 -6812 -1510 -4788
rect -1446 -6812 -1426 -4788
rect -198 -4839 -94 -4441
rect 1082 -4492 1102 -2468
rect 1166 -4492 1186 -2468
rect 2414 -2519 2518 -2121
rect 3694 -2172 3714 -148
rect 3778 -2172 3798 -148
rect 3694 -2468 3798 -2172
rect 1505 -2520 3427 -2519
rect 1505 -4440 1506 -2520
rect 3426 -4440 3427 -2520
rect 1505 -4441 3427 -4440
rect 1082 -4788 1186 -4492
rect -1107 -4840 815 -4839
rect -1107 -6760 -1106 -4840
rect 814 -6760 815 -4840
rect -1107 -6761 815 -6760
rect -1530 -7108 -1426 -6812
rect -3719 -7160 -1797 -7159
rect -3719 -9080 -3718 -7160
rect -1798 -9080 -1797 -7160
rect -3719 -9081 -1797 -9080
rect -2810 -9280 -2706 -9081
rect -1530 -9132 -1510 -7108
rect -1446 -9132 -1426 -7108
rect -198 -7159 -94 -6761
rect 1082 -6812 1102 -4788
rect 1166 -6812 1186 -4788
rect 2414 -4839 2518 -4441
rect 3694 -4492 3714 -2468
rect 3778 -4492 3798 -2468
rect 3694 -4788 3798 -4492
rect 1505 -4840 3427 -4839
rect 1505 -6760 1506 -4840
rect 3426 -6760 3427 -4840
rect 1505 -6761 3427 -6760
rect 1082 -7108 1186 -6812
rect -1107 -7160 815 -7159
rect -1107 -9080 -1106 -7160
rect 814 -9080 815 -7160
rect -1107 -9081 815 -9080
rect -1530 -9280 -1426 -9132
rect -198 -9280 -94 -9081
rect 1082 -9132 1102 -7108
rect 1166 -9132 1186 -7108
rect 2414 -7159 2518 -6761
rect 3694 -6812 3714 -4788
rect 3778 -6812 3798 -4788
rect 3694 -7108 3798 -6812
rect 1505 -7160 3427 -7159
rect 1505 -9080 1506 -7160
rect 3426 -9080 3427 -7160
rect 1505 -9081 3427 -9080
rect 1082 -9280 1186 -9132
rect 2414 -9280 2518 -9081
rect 3694 -9132 3714 -7108
rect 3778 -9132 3798 -7108
rect 3694 -9280 3798 -9132
<< properties >>
string FIXED_BBOX 1426 7080 3506 9160
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 3 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
