magic
tech sky130A
magscale 1 2
timestamp 1712087189
<< pwell >>
rect -594 -1167 594 1167
<< mvnmos >>
rect -366 109 -266 909
rect -208 109 -108 909
rect -50 109 50 909
rect 108 109 208 909
rect 266 109 366 909
rect -366 -909 -266 -109
rect -208 -909 -108 -109
rect -50 -909 50 -109
rect 108 -909 208 -109
rect 266 -909 366 -109
<< mvndiff >>
rect -424 897 -366 909
rect -424 121 -412 897
rect -378 121 -366 897
rect -424 109 -366 121
rect -266 897 -208 909
rect -266 121 -254 897
rect -220 121 -208 897
rect -266 109 -208 121
rect -108 897 -50 909
rect -108 121 -96 897
rect -62 121 -50 897
rect -108 109 -50 121
rect 50 897 108 909
rect 50 121 62 897
rect 96 121 108 897
rect 50 109 108 121
rect 208 897 266 909
rect 208 121 220 897
rect 254 121 266 897
rect 208 109 266 121
rect 366 897 424 909
rect 366 121 378 897
rect 412 121 424 897
rect 366 109 424 121
rect -424 -121 -366 -109
rect -424 -897 -412 -121
rect -378 -897 -366 -121
rect -424 -909 -366 -897
rect -266 -121 -208 -109
rect -266 -897 -254 -121
rect -220 -897 -208 -121
rect -266 -909 -208 -897
rect -108 -121 -50 -109
rect -108 -897 -96 -121
rect -62 -897 -50 -121
rect -108 -909 -50 -897
rect 50 -121 108 -109
rect 50 -897 62 -121
rect 96 -897 108 -121
rect 50 -909 108 -897
rect 208 -121 266 -109
rect 208 -897 220 -121
rect 254 -897 266 -121
rect 208 -909 266 -897
rect 366 -121 424 -109
rect 366 -897 378 -121
rect 412 -897 424 -121
rect 366 -909 424 -897
<< mvndiffc >>
rect -412 121 -378 897
rect -254 121 -220 897
rect -96 121 -62 897
rect 62 121 96 897
rect 220 121 254 897
rect 378 121 412 897
rect -412 -897 -378 -121
rect -254 -897 -220 -121
rect -96 -897 -62 -121
rect 62 -897 96 -121
rect 220 -897 254 -121
rect 378 -897 412 -121
<< mvpsubdiff >>
rect -558 1119 558 1131
rect -558 1085 -450 1119
rect 450 1085 558 1119
rect -558 1073 558 1085
rect -558 1023 -500 1073
rect -558 -1023 -546 1023
rect -512 -1023 -500 1023
rect 500 1023 558 1073
rect -558 -1073 -500 -1023
rect 500 -1023 512 1023
rect 546 -1023 558 1023
rect 500 -1073 558 -1023
rect -558 -1085 558 -1073
rect -558 -1119 -450 -1085
rect 450 -1119 558 -1085
rect -558 -1131 558 -1119
<< mvpsubdiffcont >>
rect -450 1085 450 1119
rect -546 -1023 -512 1023
rect 512 -1023 546 1023
rect -450 -1119 450 -1085
<< poly >>
rect -366 981 -266 997
rect -366 947 -350 981
rect -282 947 -266 981
rect -366 909 -266 947
rect -208 981 -108 997
rect -208 947 -192 981
rect -124 947 -108 981
rect -208 909 -108 947
rect -50 981 50 997
rect -50 947 -34 981
rect 34 947 50 981
rect -50 909 50 947
rect 108 981 208 997
rect 108 947 124 981
rect 192 947 208 981
rect 108 909 208 947
rect 266 981 366 997
rect 266 947 282 981
rect 350 947 366 981
rect 266 909 366 947
rect -366 71 -266 109
rect -366 37 -350 71
rect -282 37 -266 71
rect -366 21 -266 37
rect -208 71 -108 109
rect -208 37 -192 71
rect -124 37 -108 71
rect -208 21 -108 37
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect 108 71 208 109
rect 108 37 124 71
rect 192 37 208 71
rect 108 21 208 37
rect 266 71 366 109
rect 266 37 282 71
rect 350 37 366 71
rect 266 21 366 37
rect -366 -37 -266 -21
rect -366 -71 -350 -37
rect -282 -71 -266 -37
rect -366 -109 -266 -71
rect -208 -37 -108 -21
rect -208 -71 -192 -37
rect -124 -71 -108 -37
rect -208 -109 -108 -71
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect 108 -37 208 -21
rect 108 -71 124 -37
rect 192 -71 208 -37
rect 108 -109 208 -71
rect 266 -37 366 -21
rect 266 -71 282 -37
rect 350 -71 366 -37
rect 266 -109 366 -71
rect -366 -947 -266 -909
rect -366 -981 -350 -947
rect -282 -981 -266 -947
rect -366 -997 -266 -981
rect -208 -947 -108 -909
rect -208 -981 -192 -947
rect -124 -981 -108 -947
rect -208 -997 -108 -981
rect -50 -947 50 -909
rect -50 -981 -34 -947
rect 34 -981 50 -947
rect -50 -997 50 -981
rect 108 -947 208 -909
rect 108 -981 124 -947
rect 192 -981 208 -947
rect 108 -997 208 -981
rect 266 -947 366 -909
rect 266 -981 282 -947
rect 350 -981 366 -947
rect 266 -997 366 -981
<< polycont >>
rect -350 947 -282 981
rect -192 947 -124 981
rect -34 947 34 981
rect 124 947 192 981
rect 282 947 350 981
rect -350 37 -282 71
rect -192 37 -124 71
rect -34 37 34 71
rect 124 37 192 71
rect 282 37 350 71
rect -350 -71 -282 -37
rect -192 -71 -124 -37
rect -34 -71 34 -37
rect 124 -71 192 -37
rect 282 -71 350 -37
rect -350 -981 -282 -947
rect -192 -981 -124 -947
rect -34 -981 34 -947
rect 124 -981 192 -947
rect 282 -981 350 -947
<< locali >>
rect -546 1085 -450 1119
rect 450 1085 546 1119
rect -546 1023 -512 1085
rect 512 1023 546 1085
rect -366 947 -350 981
rect -282 947 -266 981
rect -208 947 -192 981
rect -124 947 -108 981
rect -50 947 -34 981
rect 34 947 50 981
rect 108 947 124 981
rect 192 947 208 981
rect 266 947 282 981
rect 350 947 366 981
rect -412 897 -378 913
rect -412 105 -378 121
rect -254 897 -220 913
rect -254 105 -220 121
rect -96 897 -62 913
rect -96 105 -62 121
rect 62 897 96 913
rect 62 105 96 121
rect 220 897 254 913
rect 220 105 254 121
rect 378 897 412 913
rect 378 105 412 121
rect -366 37 -350 71
rect -282 37 -266 71
rect -208 37 -192 71
rect -124 37 -108 71
rect -50 37 -34 71
rect 34 37 50 71
rect 108 37 124 71
rect 192 37 208 71
rect 266 37 282 71
rect 350 37 366 71
rect -366 -71 -350 -37
rect -282 -71 -266 -37
rect -208 -71 -192 -37
rect -124 -71 -108 -37
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect 108 -71 124 -37
rect 192 -71 208 -37
rect 266 -71 282 -37
rect 350 -71 366 -37
rect -412 -121 -378 -105
rect -412 -913 -378 -897
rect -254 -121 -220 -105
rect -254 -913 -220 -897
rect -96 -121 -62 -105
rect -96 -913 -62 -897
rect 62 -121 96 -105
rect 62 -913 96 -897
rect 220 -121 254 -105
rect 220 -913 254 -897
rect 378 -121 412 -105
rect 378 -913 412 -897
rect -366 -981 -350 -947
rect -282 -981 -266 -947
rect -208 -981 -192 -947
rect -124 -981 -108 -947
rect -50 -981 -34 -947
rect 34 -981 50 -947
rect 108 -981 124 -947
rect 192 -981 208 -947
rect 266 -981 282 -947
rect 350 -981 366 -947
rect -546 -1085 -512 -1023
rect 512 -1085 546 -1023
rect -546 -1119 -450 -1085
rect 450 -1119 546 -1085
<< viali >>
rect -350 947 -282 981
rect -192 947 -124 981
rect -34 947 34 981
rect 124 947 192 981
rect 282 947 350 981
rect -412 121 -378 897
rect -254 121 -220 897
rect -96 121 -62 897
rect 62 121 96 897
rect 220 121 254 897
rect 378 121 412 897
rect -350 37 -282 71
rect -192 37 -124 71
rect -34 37 34 71
rect 124 37 192 71
rect 282 37 350 71
rect -350 -71 -282 -37
rect -192 -71 -124 -37
rect -34 -71 34 -37
rect 124 -71 192 -37
rect 282 -71 350 -37
rect -412 -897 -378 -121
rect -254 -897 -220 -121
rect -96 -897 -62 -121
rect 62 -897 96 -121
rect 220 -897 254 -121
rect 378 -897 412 -121
rect -350 -981 -282 -947
rect -192 -981 -124 -947
rect -34 -981 34 -947
rect 124 -981 192 -947
rect 282 -981 350 -947
<< metal1 >>
rect -362 981 -270 987
rect -362 947 -350 981
rect -282 947 -270 981
rect -362 941 -270 947
rect -204 981 -112 987
rect -204 947 -192 981
rect -124 947 -112 981
rect -204 941 -112 947
rect -46 981 46 987
rect -46 947 -34 981
rect 34 947 46 981
rect -46 941 46 947
rect 112 981 204 987
rect 112 947 124 981
rect 192 947 204 981
rect 112 941 204 947
rect 270 981 362 987
rect 270 947 282 981
rect 350 947 362 981
rect 270 941 362 947
rect -418 897 -372 909
rect -418 121 -412 897
rect -378 121 -372 897
rect -418 109 -372 121
rect -260 897 -214 909
rect -260 121 -254 897
rect -220 121 -214 897
rect -260 109 -214 121
rect -102 897 -56 909
rect -102 121 -96 897
rect -62 121 -56 897
rect -102 109 -56 121
rect 56 897 102 909
rect 56 121 62 897
rect 96 121 102 897
rect 56 109 102 121
rect 214 897 260 909
rect 214 121 220 897
rect 254 121 260 897
rect 214 109 260 121
rect 372 897 418 909
rect 372 121 378 897
rect 412 121 418 897
rect 372 109 418 121
rect -362 71 -270 77
rect -362 37 -350 71
rect -282 37 -270 71
rect -362 31 -270 37
rect -204 71 -112 77
rect -204 37 -192 71
rect -124 37 -112 71
rect -204 31 -112 37
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect 112 71 204 77
rect 112 37 124 71
rect 192 37 204 71
rect 112 31 204 37
rect 270 71 362 77
rect 270 37 282 71
rect 350 37 362 71
rect 270 31 362 37
rect -362 -37 -270 -31
rect -362 -71 -350 -37
rect -282 -71 -270 -37
rect -362 -77 -270 -71
rect -204 -37 -112 -31
rect -204 -71 -192 -37
rect -124 -71 -112 -37
rect -204 -77 -112 -71
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect 112 -37 204 -31
rect 112 -71 124 -37
rect 192 -71 204 -37
rect 112 -77 204 -71
rect 270 -37 362 -31
rect 270 -71 282 -37
rect 350 -71 362 -37
rect 270 -77 362 -71
rect -418 -121 -372 -109
rect -418 -897 -412 -121
rect -378 -897 -372 -121
rect -418 -909 -372 -897
rect -260 -121 -214 -109
rect -260 -897 -254 -121
rect -220 -897 -214 -121
rect -260 -909 -214 -897
rect -102 -121 -56 -109
rect -102 -897 -96 -121
rect -62 -897 -56 -121
rect -102 -909 -56 -897
rect 56 -121 102 -109
rect 56 -897 62 -121
rect 96 -897 102 -121
rect 56 -909 102 -897
rect 214 -121 260 -109
rect 214 -897 220 -121
rect 254 -897 260 -121
rect 214 -909 260 -897
rect 372 -121 418 -109
rect 372 -897 378 -121
rect 412 -897 418 -121
rect 372 -909 418 -897
rect -362 -947 -270 -941
rect -362 -981 -350 -947
rect -282 -981 -270 -947
rect -362 -987 -270 -981
rect -204 -947 -112 -941
rect -204 -981 -192 -947
rect -124 -981 -112 -947
rect -204 -987 -112 -981
rect -46 -947 46 -941
rect -46 -981 -34 -947
rect 34 -981 46 -947
rect -46 -987 46 -981
rect 112 -947 204 -941
rect 112 -981 124 -947
rect 192 -981 204 -947
rect 112 -987 204 -981
rect 270 -947 362 -941
rect 270 -981 282 -947
rect 350 -981 362 -947
rect 270 -987 362 -981
<< properties >>
string FIXED_BBOX -529 -1102 529 1102
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 0.5 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
