magic
tech sky130A
timestamp 1712848480
<< pwell >>
rect -514 -301 514 301
<< mvnmos >>
rect -400 130 400 172
rect -400 -21 400 21
rect -400 -172 400 -130
<< mvndiff >>
rect -429 166 -400 172
rect -429 136 -423 166
rect -406 136 -400 166
rect -429 130 -400 136
rect 400 166 429 172
rect 400 136 406 166
rect 423 136 429 166
rect 400 130 429 136
rect -429 15 -400 21
rect -429 -15 -423 15
rect -406 -15 -400 15
rect -429 -21 -400 -15
rect 400 15 429 21
rect 400 -15 406 15
rect 423 -15 429 15
rect 400 -21 429 -15
rect -429 -136 -400 -130
rect -429 -166 -423 -136
rect -406 -166 -400 -136
rect -429 -172 -400 -166
rect 400 -136 429 -130
rect 400 -166 406 -136
rect 423 -166 429 -136
rect 400 -172 429 -166
<< mvndiffc >>
rect -423 136 -406 166
rect 406 136 423 166
rect -423 -15 -406 15
rect 406 -15 423 15
rect -423 -166 -406 -136
rect 406 -166 423 -136
<< mvpsubdiff >>
rect -496 277 496 283
rect -496 260 -442 277
rect 442 260 496 277
rect -496 254 496 260
rect -496 229 -467 254
rect -496 -229 -490 229
rect -473 -229 -467 229
rect 467 229 496 254
rect -496 -254 -467 -229
rect 467 -229 473 229
rect 490 -229 496 229
rect 467 -254 496 -229
rect -496 -260 496 -254
rect -496 -277 -442 -260
rect 442 -277 496 -260
rect -496 -283 496 -277
<< mvpsubdiffcont >>
rect -442 260 442 277
rect -490 -229 -473 229
rect 473 -229 490 229
rect -442 -277 442 -260
<< poly >>
rect -400 208 400 216
rect -400 191 -392 208
rect 392 191 400 208
rect -400 172 400 191
rect -400 111 400 130
rect -400 94 -392 111
rect 392 94 400 111
rect -400 86 400 94
rect -400 57 400 65
rect -400 40 -392 57
rect 392 40 400 57
rect -400 21 400 40
rect -400 -40 400 -21
rect -400 -57 -392 -40
rect 392 -57 400 -40
rect -400 -65 400 -57
rect -400 -94 400 -86
rect -400 -111 -392 -94
rect 392 -111 400 -94
rect -400 -130 400 -111
rect -400 -191 400 -172
rect -400 -208 -392 -191
rect 392 -208 400 -191
rect -400 -216 400 -208
<< polycont >>
rect -392 191 392 208
rect -392 94 392 111
rect -392 40 392 57
rect -392 -57 392 -40
rect -392 -111 392 -94
rect -392 -208 392 -191
<< locali >>
rect -490 260 -442 277
rect 442 260 490 277
rect -490 229 -473 260
rect 473 229 490 260
rect -400 191 -392 208
rect 392 191 400 208
rect -423 166 -406 174
rect -423 128 -406 136
rect 406 166 423 174
rect 406 128 423 136
rect -400 94 -392 111
rect 392 94 400 111
rect -400 40 -392 57
rect 392 40 400 57
rect -423 15 -406 23
rect -423 -23 -406 -15
rect 406 15 423 23
rect 406 -23 423 -15
rect -400 -57 -392 -40
rect 392 -57 400 -40
rect -400 -111 -392 -94
rect 392 -111 400 -94
rect -423 -136 -406 -128
rect -423 -174 -406 -166
rect 406 -136 423 -128
rect 406 -174 423 -166
rect -400 -208 -392 -191
rect 392 -208 400 -191
rect -490 -260 -473 -229
rect 473 -260 490 -229
rect -490 -277 -442 -260
rect 442 -277 490 -260
<< viali >>
rect -392 191 392 208
rect -423 136 -406 166
rect 406 136 423 166
rect -392 94 392 111
rect -392 40 392 57
rect -423 -15 -406 15
rect 406 -15 423 15
rect -392 -57 392 -40
rect -392 -111 392 -94
rect -423 -166 -406 -136
rect 406 -166 423 -136
rect -392 -208 392 -191
<< metal1 >>
rect -398 208 398 211
rect -398 191 -392 208
rect 392 191 398 208
rect -398 188 398 191
rect -426 166 -403 172
rect -426 136 -423 166
rect -406 136 -403 166
rect -426 130 -403 136
rect 403 166 426 172
rect 403 136 406 166
rect 423 136 426 166
rect 403 130 426 136
rect -398 111 398 114
rect -398 94 -392 111
rect 392 94 398 111
rect -398 91 398 94
rect -398 57 398 60
rect -398 40 -392 57
rect 392 40 398 57
rect -398 37 398 40
rect -426 15 -403 21
rect -426 -15 -423 15
rect -406 -15 -403 15
rect -426 -21 -403 -15
rect 403 15 426 21
rect 403 -15 406 15
rect 423 -15 426 15
rect 403 -21 426 -15
rect -398 -40 398 -37
rect -398 -57 -392 -40
rect 392 -57 398 -40
rect -398 -60 398 -57
rect -398 -94 398 -91
rect -398 -111 -392 -94
rect 392 -111 398 -94
rect -398 -114 398 -111
rect -426 -136 -403 -130
rect -426 -166 -423 -136
rect -406 -166 -403 -136
rect -426 -172 -403 -166
rect 403 -136 426 -130
rect 403 -166 406 -136
rect 423 -166 426 -136
rect 403 -172 426 -166
rect -398 -191 398 -188
rect -398 -208 -392 -191
rect 392 -208 398 -191
rect -398 -211 398 -208
<< properties >>
string FIXED_BBOX -481 -268 481 268
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.420 l 8 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
