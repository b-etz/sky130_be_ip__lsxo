magic
tech sky130A
magscale 1 2
timestamp 1712782684
<< nwell >>
rect -458 -4873 458 4873
<< mvpmos >>
rect -200 3776 200 4576
rect -200 2848 200 3648
rect -200 1920 200 2720
rect -200 992 200 1792
rect -200 64 200 864
rect -200 -864 200 -64
rect -200 -1792 200 -992
rect -200 -2720 200 -1920
rect -200 -3648 200 -2848
rect -200 -4576 200 -3776
<< mvpdiff >>
rect -258 4564 -200 4576
rect -258 3788 -246 4564
rect -212 3788 -200 4564
rect -258 3776 -200 3788
rect 200 4564 258 4576
rect 200 3788 212 4564
rect 246 3788 258 4564
rect 200 3776 258 3788
rect -258 3636 -200 3648
rect -258 2860 -246 3636
rect -212 2860 -200 3636
rect -258 2848 -200 2860
rect 200 3636 258 3648
rect 200 2860 212 3636
rect 246 2860 258 3636
rect 200 2848 258 2860
rect -258 2708 -200 2720
rect -258 1932 -246 2708
rect -212 1932 -200 2708
rect -258 1920 -200 1932
rect 200 2708 258 2720
rect 200 1932 212 2708
rect 246 1932 258 2708
rect 200 1920 258 1932
rect -258 1780 -200 1792
rect -258 1004 -246 1780
rect -212 1004 -200 1780
rect -258 992 -200 1004
rect 200 1780 258 1792
rect 200 1004 212 1780
rect 246 1004 258 1780
rect 200 992 258 1004
rect -258 852 -200 864
rect -258 76 -246 852
rect -212 76 -200 852
rect -258 64 -200 76
rect 200 852 258 864
rect 200 76 212 852
rect 246 76 258 852
rect 200 64 258 76
rect -258 -76 -200 -64
rect -258 -852 -246 -76
rect -212 -852 -200 -76
rect -258 -864 -200 -852
rect 200 -76 258 -64
rect 200 -852 212 -76
rect 246 -852 258 -76
rect 200 -864 258 -852
rect -258 -1004 -200 -992
rect -258 -1780 -246 -1004
rect -212 -1780 -200 -1004
rect -258 -1792 -200 -1780
rect 200 -1004 258 -992
rect 200 -1780 212 -1004
rect 246 -1780 258 -1004
rect 200 -1792 258 -1780
rect -258 -1932 -200 -1920
rect -258 -2708 -246 -1932
rect -212 -2708 -200 -1932
rect -258 -2720 -200 -2708
rect 200 -1932 258 -1920
rect 200 -2708 212 -1932
rect 246 -2708 258 -1932
rect 200 -2720 258 -2708
rect -258 -2860 -200 -2848
rect -258 -3636 -246 -2860
rect -212 -3636 -200 -2860
rect -258 -3648 -200 -3636
rect 200 -2860 258 -2848
rect 200 -3636 212 -2860
rect 246 -3636 258 -2860
rect 200 -3648 258 -3636
rect -258 -3788 -200 -3776
rect -258 -4564 -246 -3788
rect -212 -4564 -200 -3788
rect -258 -4576 -200 -4564
rect 200 -3788 258 -3776
rect 200 -4564 212 -3788
rect 246 -4564 258 -3788
rect 200 -4576 258 -4564
<< mvpdiffc >>
rect -246 3788 -212 4564
rect 212 3788 246 4564
rect -246 2860 -212 3636
rect 212 2860 246 3636
rect -246 1932 -212 2708
rect 212 1932 246 2708
rect -246 1004 -212 1780
rect 212 1004 246 1780
rect -246 76 -212 852
rect 212 76 246 852
rect -246 -852 -212 -76
rect 212 -852 246 -76
rect -246 -1780 -212 -1004
rect 212 -1780 246 -1004
rect -246 -2708 -212 -1932
rect 212 -2708 246 -1932
rect -246 -3636 -212 -2860
rect 212 -3636 246 -2860
rect -246 -4564 -212 -3788
rect 212 -4564 246 -3788
<< mvnsubdiff >>
rect -392 4795 392 4807
rect -392 4761 -284 4795
rect 284 4761 392 4795
rect -392 4749 392 4761
rect -392 4699 -334 4749
rect -392 -4699 -380 4699
rect -346 -4699 -334 4699
rect 334 4699 392 4749
rect -392 -4749 -334 -4699
rect 334 -4699 346 4699
rect 380 -4699 392 4699
rect 334 -4749 392 -4699
rect -392 -4761 392 -4749
rect -392 -4795 -284 -4761
rect 284 -4795 392 -4761
rect -392 -4807 392 -4795
<< mvnsubdiffcont >>
rect -284 4761 284 4795
rect -380 -4699 -346 4699
rect 346 -4699 380 4699
rect -284 -4795 284 -4761
<< poly >>
rect -200 4657 200 4673
rect -200 4623 -184 4657
rect 184 4623 200 4657
rect -200 4576 200 4623
rect -200 3729 200 3776
rect -200 3695 -184 3729
rect 184 3695 200 3729
rect -200 3648 200 3695
rect -200 2801 200 2848
rect -200 2767 -184 2801
rect 184 2767 200 2801
rect -200 2720 200 2767
rect -200 1873 200 1920
rect -200 1839 -184 1873
rect 184 1839 200 1873
rect -200 1792 200 1839
rect -200 945 200 992
rect -200 911 -184 945
rect 184 911 200 945
rect -200 864 200 911
rect -200 17 200 64
rect -200 -17 -184 17
rect 184 -17 200 17
rect -200 -64 200 -17
rect -200 -911 200 -864
rect -200 -945 -184 -911
rect 184 -945 200 -911
rect -200 -992 200 -945
rect -200 -1839 200 -1792
rect -200 -1873 -184 -1839
rect 184 -1873 200 -1839
rect -200 -1920 200 -1873
rect -200 -2767 200 -2720
rect -200 -2801 -184 -2767
rect 184 -2801 200 -2767
rect -200 -2848 200 -2801
rect -200 -3695 200 -3648
rect -200 -3729 -184 -3695
rect 184 -3729 200 -3695
rect -200 -3776 200 -3729
rect -200 -4623 200 -4576
rect -200 -4657 -184 -4623
rect 184 -4657 200 -4623
rect -200 -4673 200 -4657
<< polycont >>
rect -184 4623 184 4657
rect -184 3695 184 3729
rect -184 2767 184 2801
rect -184 1839 184 1873
rect -184 911 184 945
rect -184 -17 184 17
rect -184 -945 184 -911
rect -184 -1873 184 -1839
rect -184 -2801 184 -2767
rect -184 -3729 184 -3695
rect -184 -4657 184 -4623
<< locali >>
rect -380 4761 -284 4795
rect 284 4761 380 4795
rect -380 4699 -346 4761
rect 346 4699 380 4761
rect -200 4623 -184 4657
rect 184 4623 200 4657
rect -246 4564 -212 4580
rect -246 3772 -212 3788
rect 212 4564 246 4580
rect 212 3772 246 3788
rect -200 3695 -184 3729
rect 184 3695 200 3729
rect -246 3636 -212 3652
rect -246 2844 -212 2860
rect 212 3636 246 3652
rect 212 2844 246 2860
rect -200 2767 -184 2801
rect 184 2767 200 2801
rect -246 2708 -212 2724
rect -246 1916 -212 1932
rect 212 2708 246 2724
rect 212 1916 246 1932
rect -200 1839 -184 1873
rect 184 1839 200 1873
rect -246 1780 -212 1796
rect -246 988 -212 1004
rect 212 1780 246 1796
rect 212 988 246 1004
rect -200 911 -184 945
rect 184 911 200 945
rect -246 852 -212 868
rect -246 60 -212 76
rect 212 852 246 868
rect 212 60 246 76
rect -200 -17 -184 17
rect 184 -17 200 17
rect -246 -76 -212 -60
rect -246 -868 -212 -852
rect 212 -76 246 -60
rect 212 -868 246 -852
rect -200 -945 -184 -911
rect 184 -945 200 -911
rect -246 -1004 -212 -988
rect -246 -1796 -212 -1780
rect 212 -1004 246 -988
rect 212 -1796 246 -1780
rect -200 -1873 -184 -1839
rect 184 -1873 200 -1839
rect -246 -1932 -212 -1916
rect -246 -2724 -212 -2708
rect 212 -1932 246 -1916
rect 212 -2724 246 -2708
rect -200 -2801 -184 -2767
rect 184 -2801 200 -2767
rect -246 -2860 -212 -2844
rect -246 -3652 -212 -3636
rect 212 -2860 246 -2844
rect 212 -3652 246 -3636
rect -200 -3729 -184 -3695
rect 184 -3729 200 -3695
rect -246 -3788 -212 -3772
rect -246 -4580 -212 -4564
rect 212 -3788 246 -3772
rect 212 -4580 246 -4564
rect -200 -4657 -184 -4623
rect 184 -4657 200 -4623
rect -380 -4761 -346 -4699
rect 346 -4761 380 -4699
rect -380 -4795 -284 -4761
rect 284 -4795 380 -4761
<< viali >>
rect -184 4623 184 4657
rect -246 3788 -212 4564
rect 212 3788 246 4564
rect -184 3695 184 3729
rect -246 2860 -212 3636
rect 212 2860 246 3636
rect -184 2767 184 2801
rect -246 1932 -212 2708
rect 212 1932 246 2708
rect -184 1839 184 1873
rect -246 1004 -212 1780
rect 212 1004 246 1780
rect -184 911 184 945
rect -246 76 -212 852
rect 212 76 246 852
rect -184 -17 184 17
rect -246 -852 -212 -76
rect 212 -852 246 -76
rect -184 -945 184 -911
rect -246 -1780 -212 -1004
rect 212 -1780 246 -1004
rect -184 -1873 184 -1839
rect -246 -2708 -212 -1932
rect 212 -2708 246 -1932
rect -184 -2801 184 -2767
rect -246 -3636 -212 -2860
rect 212 -3636 246 -2860
rect -184 -3729 184 -3695
rect -246 -4564 -212 -3788
rect 212 -4564 246 -3788
rect -184 -4657 184 -4623
<< metal1 >>
rect -196 4657 196 4663
rect -196 4623 -184 4657
rect 184 4623 196 4657
rect -196 4617 196 4623
rect -252 4564 -206 4576
rect -252 3788 -246 4564
rect -212 3788 -206 4564
rect -252 3776 -206 3788
rect 206 4564 252 4576
rect 206 3788 212 4564
rect 246 3788 252 4564
rect 206 3776 252 3788
rect -196 3729 196 3735
rect -196 3695 -184 3729
rect 184 3695 196 3729
rect -196 3689 196 3695
rect -252 3636 -206 3648
rect -252 2860 -246 3636
rect -212 2860 -206 3636
rect -252 2848 -206 2860
rect 206 3636 252 3648
rect 206 2860 212 3636
rect 246 2860 252 3636
rect 206 2848 252 2860
rect -196 2801 196 2807
rect -196 2767 -184 2801
rect 184 2767 196 2801
rect -196 2761 196 2767
rect -252 2708 -206 2720
rect -252 1932 -246 2708
rect -212 1932 -206 2708
rect -252 1920 -206 1932
rect 206 2708 252 2720
rect 206 1932 212 2708
rect 246 1932 252 2708
rect 206 1920 252 1932
rect -196 1873 196 1879
rect -196 1839 -184 1873
rect 184 1839 196 1873
rect -196 1833 196 1839
rect -252 1780 -206 1792
rect -252 1004 -246 1780
rect -212 1004 -206 1780
rect -252 992 -206 1004
rect 206 1780 252 1792
rect 206 1004 212 1780
rect 246 1004 252 1780
rect 206 992 252 1004
rect -196 945 196 951
rect -196 911 -184 945
rect 184 911 196 945
rect -196 905 196 911
rect -252 852 -206 864
rect -252 76 -246 852
rect -212 76 -206 852
rect -252 64 -206 76
rect 206 852 252 864
rect 206 76 212 852
rect 246 76 252 852
rect 206 64 252 76
rect -196 17 196 23
rect -196 -17 -184 17
rect 184 -17 196 17
rect -196 -23 196 -17
rect -252 -76 -206 -64
rect -252 -852 -246 -76
rect -212 -852 -206 -76
rect -252 -864 -206 -852
rect 206 -76 252 -64
rect 206 -852 212 -76
rect 246 -852 252 -76
rect 206 -864 252 -852
rect -196 -911 196 -905
rect -196 -945 -184 -911
rect 184 -945 196 -911
rect -196 -951 196 -945
rect -252 -1004 -206 -992
rect -252 -1780 -246 -1004
rect -212 -1780 -206 -1004
rect -252 -1792 -206 -1780
rect 206 -1004 252 -992
rect 206 -1780 212 -1004
rect 246 -1780 252 -1004
rect 206 -1792 252 -1780
rect -196 -1839 196 -1833
rect -196 -1873 -184 -1839
rect 184 -1873 196 -1839
rect -196 -1879 196 -1873
rect -252 -1932 -206 -1920
rect -252 -2708 -246 -1932
rect -212 -2708 -206 -1932
rect -252 -2720 -206 -2708
rect 206 -1932 252 -1920
rect 206 -2708 212 -1932
rect 246 -2708 252 -1932
rect 206 -2720 252 -2708
rect -196 -2767 196 -2761
rect -196 -2801 -184 -2767
rect 184 -2801 196 -2767
rect -196 -2807 196 -2801
rect -252 -2860 -206 -2848
rect -252 -3636 -246 -2860
rect -212 -3636 -206 -2860
rect -252 -3648 -206 -3636
rect 206 -2860 252 -2848
rect 206 -3636 212 -2860
rect 246 -3636 252 -2860
rect 206 -3648 252 -3636
rect -196 -3695 196 -3689
rect -196 -3729 -184 -3695
rect 184 -3729 196 -3695
rect -196 -3735 196 -3729
rect -252 -3788 -206 -3776
rect -252 -4564 -246 -3788
rect -212 -4564 -206 -3788
rect -252 -4576 -206 -4564
rect 206 -3788 252 -3776
rect 206 -4564 212 -3788
rect 246 -4564 252 -3788
rect 206 -4576 252 -4564
rect -196 -4623 196 -4617
rect -196 -4657 -184 -4623
rect 184 -4657 196 -4623
rect -196 -4663 196 -4657
<< properties >>
string FIXED_BBOX -363 -4778 363 4778
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 2.0 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
