magic
tech sky130A
magscale 1 2
timestamp 1712946411
<< pwell >>
rect -2193 -9082 2193 9082
<< psubdiff >>
rect -2157 9012 -2061 9046
rect 2061 9012 2157 9046
rect -2157 8950 -2123 9012
rect 2123 8950 2157 9012
rect -2157 -9012 -2123 -8950
rect 2123 -9012 2157 -8950
rect -2157 -9046 -2061 -9012
rect 2061 -9046 2157 -9012
<< psubdiffcont >>
rect -2061 9012 2061 9046
rect -2157 -8950 -2123 8950
rect 2123 -8950 2157 8950
rect -2061 -9046 2061 -9012
<< xpolycontact >>
rect -2027 8484 -1957 8916
rect -2027 -8916 -1957 -8484
rect -1861 8484 -1791 8916
rect -1861 -8916 -1791 -8484
rect -1695 8484 -1625 8916
rect -1695 -8916 -1625 -8484
rect -1529 8484 -1459 8916
rect -1529 -8916 -1459 -8484
rect -1363 8484 -1293 8916
rect -1363 -8916 -1293 -8484
rect -1197 8484 -1127 8916
rect -1197 -8916 -1127 -8484
rect -1031 8484 -961 8916
rect -1031 -8916 -961 -8484
rect -865 8484 -795 8916
rect -865 -8916 -795 -8484
rect -699 8484 -629 8916
rect -699 -8916 -629 -8484
rect -533 8484 -463 8916
rect -533 -8916 -463 -8484
rect -367 8484 -297 8916
rect -367 -8916 -297 -8484
rect -201 8484 -131 8916
rect -201 -8916 -131 -8484
rect -35 8484 35 8916
rect -35 -8916 35 -8484
rect 131 8484 201 8916
rect 131 -8916 201 -8484
rect 297 8484 367 8916
rect 297 -8916 367 -8484
rect 463 8484 533 8916
rect 463 -8916 533 -8484
rect 629 8484 699 8916
rect 629 -8916 699 -8484
rect 795 8484 865 8916
rect 795 -8916 865 -8484
rect 961 8484 1031 8916
rect 961 -8916 1031 -8484
rect 1127 8484 1197 8916
rect 1127 -8916 1197 -8484
rect 1293 8484 1363 8916
rect 1293 -8916 1363 -8484
rect 1459 8484 1529 8916
rect 1459 -8916 1529 -8484
rect 1625 8484 1695 8916
rect 1625 -8916 1695 -8484
rect 1791 8484 1861 8916
rect 1791 -8916 1861 -8484
rect 1957 8484 2027 8916
rect 1957 -8916 2027 -8484
<< xpolyres >>
rect -2027 -8484 -1957 8484
rect -1861 -8484 -1791 8484
rect -1695 -8484 -1625 8484
rect -1529 -8484 -1459 8484
rect -1363 -8484 -1293 8484
rect -1197 -8484 -1127 8484
rect -1031 -8484 -961 8484
rect -865 -8484 -795 8484
rect -699 -8484 -629 8484
rect -533 -8484 -463 8484
rect -367 -8484 -297 8484
rect -201 -8484 -131 8484
rect -35 -8484 35 8484
rect 131 -8484 201 8484
rect 297 -8484 367 8484
rect 463 -8484 533 8484
rect 629 -8484 699 8484
rect 795 -8484 865 8484
rect 961 -8484 1031 8484
rect 1127 -8484 1197 8484
rect 1293 -8484 1363 8484
rect 1459 -8484 1529 8484
rect 1625 -8484 1695 8484
rect 1791 -8484 1861 8484
rect 1957 -8484 2027 8484
<< locali >>
rect -2157 9012 -2061 9046
rect 2061 9012 2157 9046
rect -2157 8950 -2123 9012
rect 2123 8950 2157 9012
rect -2157 -9012 -2123 -8950
rect 2123 -9012 2157 -8950
rect -2157 -9046 -2061 -9012
rect 2061 -9046 2157 -9012
<< viali >>
rect -2011 8501 -1973 8898
rect -1845 8501 -1807 8898
rect -1679 8501 -1641 8898
rect -1513 8501 -1475 8898
rect -1347 8501 -1309 8898
rect -1181 8501 -1143 8898
rect -1015 8501 -977 8898
rect -849 8501 -811 8898
rect -683 8501 -645 8898
rect -517 8501 -479 8898
rect -351 8501 -313 8898
rect -185 8501 -147 8898
rect -19 8501 19 8898
rect 147 8501 185 8898
rect 313 8501 351 8898
rect 479 8501 517 8898
rect 645 8501 683 8898
rect 811 8501 849 8898
rect 977 8501 1015 8898
rect 1143 8501 1181 8898
rect 1309 8501 1347 8898
rect 1475 8501 1513 8898
rect 1641 8501 1679 8898
rect 1807 8501 1845 8898
rect 1973 8501 2011 8898
rect -2011 -8898 -1973 -8501
rect -1845 -8898 -1807 -8501
rect -1679 -8898 -1641 -8501
rect -1513 -8898 -1475 -8501
rect -1347 -8898 -1309 -8501
rect -1181 -8898 -1143 -8501
rect -1015 -8898 -977 -8501
rect -849 -8898 -811 -8501
rect -683 -8898 -645 -8501
rect -517 -8898 -479 -8501
rect -351 -8898 -313 -8501
rect -185 -8898 -147 -8501
rect -19 -8898 19 -8501
rect 147 -8898 185 -8501
rect 313 -8898 351 -8501
rect 479 -8898 517 -8501
rect 645 -8898 683 -8501
rect 811 -8898 849 -8501
rect 977 -8898 1015 -8501
rect 1143 -8898 1181 -8501
rect 1309 -8898 1347 -8501
rect 1475 -8898 1513 -8501
rect 1641 -8898 1679 -8501
rect 1807 -8898 1845 -8501
rect 1973 -8898 2011 -8501
<< metal1 >>
rect -2017 8898 -1967 8910
rect -2017 8501 -2011 8898
rect -1973 8501 -1967 8898
rect -2017 8489 -1967 8501
rect -1851 8898 -1801 8910
rect -1851 8501 -1845 8898
rect -1807 8501 -1801 8898
rect -1851 8489 -1801 8501
rect -1685 8898 -1635 8910
rect -1685 8501 -1679 8898
rect -1641 8501 -1635 8898
rect -1685 8489 -1635 8501
rect -1519 8898 -1469 8910
rect -1519 8501 -1513 8898
rect -1475 8501 -1469 8898
rect -1519 8489 -1469 8501
rect -1353 8898 -1303 8910
rect -1353 8501 -1347 8898
rect -1309 8501 -1303 8898
rect -1353 8489 -1303 8501
rect -1187 8898 -1137 8910
rect -1187 8501 -1181 8898
rect -1143 8501 -1137 8898
rect -1187 8489 -1137 8501
rect -1021 8898 -971 8910
rect -1021 8501 -1015 8898
rect -977 8501 -971 8898
rect -1021 8489 -971 8501
rect -855 8898 -805 8910
rect -855 8501 -849 8898
rect -811 8501 -805 8898
rect -855 8489 -805 8501
rect -689 8898 -639 8910
rect -689 8501 -683 8898
rect -645 8501 -639 8898
rect -689 8489 -639 8501
rect -523 8898 -473 8910
rect -523 8501 -517 8898
rect -479 8501 -473 8898
rect -523 8489 -473 8501
rect -357 8898 -307 8910
rect -357 8501 -351 8898
rect -313 8501 -307 8898
rect -357 8489 -307 8501
rect -191 8898 -141 8910
rect -191 8501 -185 8898
rect -147 8501 -141 8898
rect -191 8489 -141 8501
rect -25 8898 25 8910
rect -25 8501 -19 8898
rect 19 8501 25 8898
rect -25 8489 25 8501
rect 141 8898 191 8910
rect 141 8501 147 8898
rect 185 8501 191 8898
rect 141 8489 191 8501
rect 307 8898 357 8910
rect 307 8501 313 8898
rect 351 8501 357 8898
rect 307 8489 357 8501
rect 473 8898 523 8910
rect 473 8501 479 8898
rect 517 8501 523 8898
rect 473 8489 523 8501
rect 639 8898 689 8910
rect 639 8501 645 8898
rect 683 8501 689 8898
rect 639 8489 689 8501
rect 805 8898 855 8910
rect 805 8501 811 8898
rect 849 8501 855 8898
rect 805 8489 855 8501
rect 971 8898 1021 8910
rect 971 8501 977 8898
rect 1015 8501 1021 8898
rect 971 8489 1021 8501
rect 1137 8898 1187 8910
rect 1137 8501 1143 8898
rect 1181 8501 1187 8898
rect 1137 8489 1187 8501
rect 1303 8898 1353 8910
rect 1303 8501 1309 8898
rect 1347 8501 1353 8898
rect 1303 8489 1353 8501
rect 1469 8898 1519 8910
rect 1469 8501 1475 8898
rect 1513 8501 1519 8898
rect 1469 8489 1519 8501
rect 1635 8898 1685 8910
rect 1635 8501 1641 8898
rect 1679 8501 1685 8898
rect 1635 8489 1685 8501
rect 1801 8898 1851 8910
rect 1801 8501 1807 8898
rect 1845 8501 1851 8898
rect 1801 8489 1851 8501
rect 1967 8898 2017 8910
rect 1967 8501 1973 8898
rect 2011 8501 2017 8898
rect 1967 8489 2017 8501
rect -2017 -8501 -1967 -8489
rect -2017 -8898 -2011 -8501
rect -1973 -8898 -1967 -8501
rect -2017 -8910 -1967 -8898
rect -1851 -8501 -1801 -8489
rect -1851 -8898 -1845 -8501
rect -1807 -8898 -1801 -8501
rect -1851 -8910 -1801 -8898
rect -1685 -8501 -1635 -8489
rect -1685 -8898 -1679 -8501
rect -1641 -8898 -1635 -8501
rect -1685 -8910 -1635 -8898
rect -1519 -8501 -1469 -8489
rect -1519 -8898 -1513 -8501
rect -1475 -8898 -1469 -8501
rect -1519 -8910 -1469 -8898
rect -1353 -8501 -1303 -8489
rect -1353 -8898 -1347 -8501
rect -1309 -8898 -1303 -8501
rect -1353 -8910 -1303 -8898
rect -1187 -8501 -1137 -8489
rect -1187 -8898 -1181 -8501
rect -1143 -8898 -1137 -8501
rect -1187 -8910 -1137 -8898
rect -1021 -8501 -971 -8489
rect -1021 -8898 -1015 -8501
rect -977 -8898 -971 -8501
rect -1021 -8910 -971 -8898
rect -855 -8501 -805 -8489
rect -855 -8898 -849 -8501
rect -811 -8898 -805 -8501
rect -855 -8910 -805 -8898
rect -689 -8501 -639 -8489
rect -689 -8898 -683 -8501
rect -645 -8898 -639 -8501
rect -689 -8910 -639 -8898
rect -523 -8501 -473 -8489
rect -523 -8898 -517 -8501
rect -479 -8898 -473 -8501
rect -523 -8910 -473 -8898
rect -357 -8501 -307 -8489
rect -357 -8898 -351 -8501
rect -313 -8898 -307 -8501
rect -357 -8910 -307 -8898
rect -191 -8501 -141 -8489
rect -191 -8898 -185 -8501
rect -147 -8898 -141 -8501
rect -191 -8910 -141 -8898
rect -25 -8501 25 -8489
rect -25 -8898 -19 -8501
rect 19 -8898 25 -8501
rect -25 -8910 25 -8898
rect 141 -8501 191 -8489
rect 141 -8898 147 -8501
rect 185 -8898 191 -8501
rect 141 -8910 191 -8898
rect 307 -8501 357 -8489
rect 307 -8898 313 -8501
rect 351 -8898 357 -8501
rect 307 -8910 357 -8898
rect 473 -8501 523 -8489
rect 473 -8898 479 -8501
rect 517 -8898 523 -8501
rect 473 -8910 523 -8898
rect 639 -8501 689 -8489
rect 639 -8898 645 -8501
rect 683 -8898 689 -8501
rect 639 -8910 689 -8898
rect 805 -8501 855 -8489
rect 805 -8898 811 -8501
rect 849 -8898 855 -8501
rect 805 -8910 855 -8898
rect 971 -8501 1021 -8489
rect 971 -8898 977 -8501
rect 1015 -8898 1021 -8501
rect 971 -8910 1021 -8898
rect 1137 -8501 1187 -8489
rect 1137 -8898 1143 -8501
rect 1181 -8898 1187 -8501
rect 1137 -8910 1187 -8898
rect 1303 -8501 1353 -8489
rect 1303 -8898 1309 -8501
rect 1347 -8898 1353 -8501
rect 1303 -8910 1353 -8898
rect 1469 -8501 1519 -8489
rect 1469 -8898 1475 -8501
rect 1513 -8898 1519 -8501
rect 1469 -8910 1519 -8898
rect 1635 -8501 1685 -8489
rect 1635 -8898 1641 -8501
rect 1679 -8898 1685 -8501
rect 1635 -8910 1685 -8898
rect 1801 -8501 1851 -8489
rect 1801 -8898 1807 -8501
rect 1845 -8898 1851 -8501
rect 1801 -8910 1851 -8898
rect 1967 -8501 2017 -8489
rect 1967 -8898 1973 -8501
rect 2011 -8898 2017 -8501
rect 1967 -8910 2017 -8898
<< properties >>
string FIXED_BBOX -2140 -9029 2140 9029
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 85 m 1 nx 25 wmin 0.350 lmin 0.50 rho 2000 val 486.789k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
