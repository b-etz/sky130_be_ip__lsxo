magic
tech sky130A
magscale 1 2
timestamp 1712073300
<< metal3 >>
rect -6410 36972 -4038 37000
rect -6410 34948 -4122 36972
rect -4058 34948 -4038 36972
rect -6410 34920 -4038 34948
rect -3798 36972 -1426 37000
rect -3798 34948 -1510 36972
rect -1446 34948 -1426 36972
rect -3798 34920 -1426 34948
rect -1186 36972 1186 37000
rect -1186 34948 1102 36972
rect 1166 34948 1186 36972
rect -1186 34920 1186 34948
rect 1426 36972 3798 37000
rect 1426 34948 3714 36972
rect 3778 34948 3798 36972
rect 1426 34920 3798 34948
rect 4038 36972 6410 37000
rect 4038 34948 6326 36972
rect 6390 34948 6410 36972
rect 4038 34920 6410 34948
rect -6410 34652 -4038 34680
rect -6410 32628 -4122 34652
rect -4058 32628 -4038 34652
rect -6410 32600 -4038 32628
rect -3798 34652 -1426 34680
rect -3798 32628 -1510 34652
rect -1446 32628 -1426 34652
rect -3798 32600 -1426 32628
rect -1186 34652 1186 34680
rect -1186 32628 1102 34652
rect 1166 32628 1186 34652
rect -1186 32600 1186 32628
rect 1426 34652 3798 34680
rect 1426 32628 3714 34652
rect 3778 32628 3798 34652
rect 1426 32600 3798 32628
rect 4038 34652 6410 34680
rect 4038 32628 6326 34652
rect 6390 32628 6410 34652
rect 4038 32600 6410 32628
rect -6410 32332 -4038 32360
rect -6410 30308 -4122 32332
rect -4058 30308 -4038 32332
rect -6410 30280 -4038 30308
rect -3798 32332 -1426 32360
rect -3798 30308 -1510 32332
rect -1446 30308 -1426 32332
rect -3798 30280 -1426 30308
rect -1186 32332 1186 32360
rect -1186 30308 1102 32332
rect 1166 30308 1186 32332
rect -1186 30280 1186 30308
rect 1426 32332 3798 32360
rect 1426 30308 3714 32332
rect 3778 30308 3798 32332
rect 1426 30280 3798 30308
rect 4038 32332 6410 32360
rect 4038 30308 6326 32332
rect 6390 30308 6410 32332
rect 4038 30280 6410 30308
rect -6410 30012 -4038 30040
rect -6410 27988 -4122 30012
rect -4058 27988 -4038 30012
rect -6410 27960 -4038 27988
rect -3798 30012 -1426 30040
rect -3798 27988 -1510 30012
rect -1446 27988 -1426 30012
rect -3798 27960 -1426 27988
rect -1186 30012 1186 30040
rect -1186 27988 1102 30012
rect 1166 27988 1186 30012
rect -1186 27960 1186 27988
rect 1426 30012 3798 30040
rect 1426 27988 3714 30012
rect 3778 27988 3798 30012
rect 1426 27960 3798 27988
rect 4038 30012 6410 30040
rect 4038 27988 6326 30012
rect 6390 27988 6410 30012
rect 4038 27960 6410 27988
rect -6410 27692 -4038 27720
rect -6410 25668 -4122 27692
rect -4058 25668 -4038 27692
rect -6410 25640 -4038 25668
rect -3798 27692 -1426 27720
rect -3798 25668 -1510 27692
rect -1446 25668 -1426 27692
rect -3798 25640 -1426 25668
rect -1186 27692 1186 27720
rect -1186 25668 1102 27692
rect 1166 25668 1186 27692
rect -1186 25640 1186 25668
rect 1426 27692 3798 27720
rect 1426 25668 3714 27692
rect 3778 25668 3798 27692
rect 1426 25640 3798 25668
rect 4038 27692 6410 27720
rect 4038 25668 6326 27692
rect 6390 25668 6410 27692
rect 4038 25640 6410 25668
rect -6410 25372 -4038 25400
rect -6410 23348 -4122 25372
rect -4058 23348 -4038 25372
rect -6410 23320 -4038 23348
rect -3798 25372 -1426 25400
rect -3798 23348 -1510 25372
rect -1446 23348 -1426 25372
rect -3798 23320 -1426 23348
rect -1186 25372 1186 25400
rect -1186 23348 1102 25372
rect 1166 23348 1186 25372
rect -1186 23320 1186 23348
rect 1426 25372 3798 25400
rect 1426 23348 3714 25372
rect 3778 23348 3798 25372
rect 1426 23320 3798 23348
rect 4038 25372 6410 25400
rect 4038 23348 6326 25372
rect 6390 23348 6410 25372
rect 4038 23320 6410 23348
rect -6410 23052 -4038 23080
rect -6410 21028 -4122 23052
rect -4058 21028 -4038 23052
rect -6410 21000 -4038 21028
rect -3798 23052 -1426 23080
rect -3798 21028 -1510 23052
rect -1446 21028 -1426 23052
rect -3798 21000 -1426 21028
rect -1186 23052 1186 23080
rect -1186 21028 1102 23052
rect 1166 21028 1186 23052
rect -1186 21000 1186 21028
rect 1426 23052 3798 23080
rect 1426 21028 3714 23052
rect 3778 21028 3798 23052
rect 1426 21000 3798 21028
rect 4038 23052 6410 23080
rect 4038 21028 6326 23052
rect 6390 21028 6410 23052
rect 4038 21000 6410 21028
rect -6410 20732 -4038 20760
rect -6410 18708 -4122 20732
rect -4058 18708 -4038 20732
rect -6410 18680 -4038 18708
rect -3798 20732 -1426 20760
rect -3798 18708 -1510 20732
rect -1446 18708 -1426 20732
rect -3798 18680 -1426 18708
rect -1186 20732 1186 20760
rect -1186 18708 1102 20732
rect 1166 18708 1186 20732
rect -1186 18680 1186 18708
rect 1426 20732 3798 20760
rect 1426 18708 3714 20732
rect 3778 18708 3798 20732
rect 1426 18680 3798 18708
rect 4038 20732 6410 20760
rect 4038 18708 6326 20732
rect 6390 18708 6410 20732
rect 4038 18680 6410 18708
rect -6410 18412 -4038 18440
rect -6410 16388 -4122 18412
rect -4058 16388 -4038 18412
rect -6410 16360 -4038 16388
rect -3798 18412 -1426 18440
rect -3798 16388 -1510 18412
rect -1446 16388 -1426 18412
rect -3798 16360 -1426 16388
rect -1186 18412 1186 18440
rect -1186 16388 1102 18412
rect 1166 16388 1186 18412
rect -1186 16360 1186 16388
rect 1426 18412 3798 18440
rect 1426 16388 3714 18412
rect 3778 16388 3798 18412
rect 1426 16360 3798 16388
rect 4038 18412 6410 18440
rect 4038 16388 6326 18412
rect 6390 16388 6410 18412
rect 4038 16360 6410 16388
rect -6410 16092 -4038 16120
rect -6410 14068 -4122 16092
rect -4058 14068 -4038 16092
rect -6410 14040 -4038 14068
rect -3798 16092 -1426 16120
rect -3798 14068 -1510 16092
rect -1446 14068 -1426 16092
rect -3798 14040 -1426 14068
rect -1186 16092 1186 16120
rect -1186 14068 1102 16092
rect 1166 14068 1186 16092
rect -1186 14040 1186 14068
rect 1426 16092 3798 16120
rect 1426 14068 3714 16092
rect 3778 14068 3798 16092
rect 1426 14040 3798 14068
rect 4038 16092 6410 16120
rect 4038 14068 6326 16092
rect 6390 14068 6410 16092
rect 4038 14040 6410 14068
rect -6410 13772 -4038 13800
rect -6410 11748 -4122 13772
rect -4058 11748 -4038 13772
rect -6410 11720 -4038 11748
rect -3798 13772 -1426 13800
rect -3798 11748 -1510 13772
rect -1446 11748 -1426 13772
rect -3798 11720 -1426 11748
rect -1186 13772 1186 13800
rect -1186 11748 1102 13772
rect 1166 11748 1186 13772
rect -1186 11720 1186 11748
rect 1426 13772 3798 13800
rect 1426 11748 3714 13772
rect 3778 11748 3798 13772
rect 1426 11720 3798 11748
rect 4038 13772 6410 13800
rect 4038 11748 6326 13772
rect 6390 11748 6410 13772
rect 4038 11720 6410 11748
rect -6410 11452 -4038 11480
rect -6410 9428 -4122 11452
rect -4058 9428 -4038 11452
rect -6410 9400 -4038 9428
rect -3798 11452 -1426 11480
rect -3798 9428 -1510 11452
rect -1446 9428 -1426 11452
rect -3798 9400 -1426 9428
rect -1186 11452 1186 11480
rect -1186 9428 1102 11452
rect 1166 9428 1186 11452
rect -1186 9400 1186 9428
rect 1426 11452 3798 11480
rect 1426 9428 3714 11452
rect 3778 9428 3798 11452
rect 1426 9400 3798 9428
rect 4038 11452 6410 11480
rect 4038 9428 6326 11452
rect 6390 9428 6410 11452
rect 4038 9400 6410 9428
rect -6410 9132 -4038 9160
rect -6410 7108 -4122 9132
rect -4058 7108 -4038 9132
rect -6410 7080 -4038 7108
rect -3798 9132 -1426 9160
rect -3798 7108 -1510 9132
rect -1446 7108 -1426 9132
rect -3798 7080 -1426 7108
rect -1186 9132 1186 9160
rect -1186 7108 1102 9132
rect 1166 7108 1186 9132
rect -1186 7080 1186 7108
rect 1426 9132 3798 9160
rect 1426 7108 3714 9132
rect 3778 7108 3798 9132
rect 1426 7080 3798 7108
rect 4038 9132 6410 9160
rect 4038 7108 6326 9132
rect 6390 7108 6410 9132
rect 4038 7080 6410 7108
rect -6410 6812 -4038 6840
rect -6410 4788 -4122 6812
rect -4058 4788 -4038 6812
rect -6410 4760 -4038 4788
rect -3798 6812 -1426 6840
rect -3798 4788 -1510 6812
rect -1446 4788 -1426 6812
rect -3798 4760 -1426 4788
rect -1186 6812 1186 6840
rect -1186 4788 1102 6812
rect 1166 4788 1186 6812
rect -1186 4760 1186 4788
rect 1426 6812 3798 6840
rect 1426 4788 3714 6812
rect 3778 4788 3798 6812
rect 1426 4760 3798 4788
rect 4038 6812 6410 6840
rect 4038 4788 6326 6812
rect 6390 4788 6410 6812
rect 4038 4760 6410 4788
rect -6410 4492 -4038 4520
rect -6410 2468 -4122 4492
rect -4058 2468 -4038 4492
rect -6410 2440 -4038 2468
rect -3798 4492 -1426 4520
rect -3798 2468 -1510 4492
rect -1446 2468 -1426 4492
rect -3798 2440 -1426 2468
rect -1186 4492 1186 4520
rect -1186 2468 1102 4492
rect 1166 2468 1186 4492
rect -1186 2440 1186 2468
rect 1426 4492 3798 4520
rect 1426 2468 3714 4492
rect 3778 2468 3798 4492
rect 1426 2440 3798 2468
rect 4038 4492 6410 4520
rect 4038 2468 6326 4492
rect 6390 2468 6410 4492
rect 4038 2440 6410 2468
rect -6410 2172 -4038 2200
rect -6410 148 -4122 2172
rect -4058 148 -4038 2172
rect -6410 120 -4038 148
rect -3798 2172 -1426 2200
rect -3798 148 -1510 2172
rect -1446 148 -1426 2172
rect -3798 120 -1426 148
rect -1186 2172 1186 2200
rect -1186 148 1102 2172
rect 1166 148 1186 2172
rect -1186 120 1186 148
rect 1426 2172 3798 2200
rect 1426 148 3714 2172
rect 3778 148 3798 2172
rect 1426 120 3798 148
rect 4038 2172 6410 2200
rect 4038 148 6326 2172
rect 6390 148 6410 2172
rect 4038 120 6410 148
rect -6410 -148 -4038 -120
rect -6410 -2172 -4122 -148
rect -4058 -2172 -4038 -148
rect -6410 -2200 -4038 -2172
rect -3798 -148 -1426 -120
rect -3798 -2172 -1510 -148
rect -1446 -2172 -1426 -148
rect -3798 -2200 -1426 -2172
rect -1186 -148 1186 -120
rect -1186 -2172 1102 -148
rect 1166 -2172 1186 -148
rect -1186 -2200 1186 -2172
rect 1426 -148 3798 -120
rect 1426 -2172 3714 -148
rect 3778 -2172 3798 -148
rect 1426 -2200 3798 -2172
rect 4038 -148 6410 -120
rect 4038 -2172 6326 -148
rect 6390 -2172 6410 -148
rect 4038 -2200 6410 -2172
rect -6410 -2468 -4038 -2440
rect -6410 -4492 -4122 -2468
rect -4058 -4492 -4038 -2468
rect -6410 -4520 -4038 -4492
rect -3798 -2468 -1426 -2440
rect -3798 -4492 -1510 -2468
rect -1446 -4492 -1426 -2468
rect -3798 -4520 -1426 -4492
rect -1186 -2468 1186 -2440
rect -1186 -4492 1102 -2468
rect 1166 -4492 1186 -2468
rect -1186 -4520 1186 -4492
rect 1426 -2468 3798 -2440
rect 1426 -4492 3714 -2468
rect 3778 -4492 3798 -2468
rect 1426 -4520 3798 -4492
rect 4038 -2468 6410 -2440
rect 4038 -4492 6326 -2468
rect 6390 -4492 6410 -2468
rect 4038 -4520 6410 -4492
rect -6410 -4788 -4038 -4760
rect -6410 -6812 -4122 -4788
rect -4058 -6812 -4038 -4788
rect -6410 -6840 -4038 -6812
rect -3798 -4788 -1426 -4760
rect -3798 -6812 -1510 -4788
rect -1446 -6812 -1426 -4788
rect -3798 -6840 -1426 -6812
rect -1186 -4788 1186 -4760
rect -1186 -6812 1102 -4788
rect 1166 -6812 1186 -4788
rect -1186 -6840 1186 -6812
rect 1426 -4788 3798 -4760
rect 1426 -6812 3714 -4788
rect 3778 -6812 3798 -4788
rect 1426 -6840 3798 -6812
rect 4038 -4788 6410 -4760
rect 4038 -6812 6326 -4788
rect 6390 -6812 6410 -4788
rect 4038 -6840 6410 -6812
rect -6410 -7108 -4038 -7080
rect -6410 -9132 -4122 -7108
rect -4058 -9132 -4038 -7108
rect -6410 -9160 -4038 -9132
rect -3798 -7108 -1426 -7080
rect -3798 -9132 -1510 -7108
rect -1446 -9132 -1426 -7108
rect -3798 -9160 -1426 -9132
rect -1186 -7108 1186 -7080
rect -1186 -9132 1102 -7108
rect 1166 -9132 1186 -7108
rect -1186 -9160 1186 -9132
rect 1426 -7108 3798 -7080
rect 1426 -9132 3714 -7108
rect 3778 -9132 3798 -7108
rect 1426 -9160 3798 -9132
rect 4038 -7108 6410 -7080
rect 4038 -9132 6326 -7108
rect 6390 -9132 6410 -7108
rect 4038 -9160 6410 -9132
rect -6410 -9428 -4038 -9400
rect -6410 -11452 -4122 -9428
rect -4058 -11452 -4038 -9428
rect -6410 -11480 -4038 -11452
rect -3798 -9428 -1426 -9400
rect -3798 -11452 -1510 -9428
rect -1446 -11452 -1426 -9428
rect -3798 -11480 -1426 -11452
rect -1186 -9428 1186 -9400
rect -1186 -11452 1102 -9428
rect 1166 -11452 1186 -9428
rect -1186 -11480 1186 -11452
rect 1426 -9428 3798 -9400
rect 1426 -11452 3714 -9428
rect 3778 -11452 3798 -9428
rect 1426 -11480 3798 -11452
rect 4038 -9428 6410 -9400
rect 4038 -11452 6326 -9428
rect 6390 -11452 6410 -9428
rect 4038 -11480 6410 -11452
rect -6410 -11748 -4038 -11720
rect -6410 -13772 -4122 -11748
rect -4058 -13772 -4038 -11748
rect -6410 -13800 -4038 -13772
rect -3798 -11748 -1426 -11720
rect -3798 -13772 -1510 -11748
rect -1446 -13772 -1426 -11748
rect -3798 -13800 -1426 -13772
rect -1186 -11748 1186 -11720
rect -1186 -13772 1102 -11748
rect 1166 -13772 1186 -11748
rect -1186 -13800 1186 -13772
rect 1426 -11748 3798 -11720
rect 1426 -13772 3714 -11748
rect 3778 -13772 3798 -11748
rect 1426 -13800 3798 -13772
rect 4038 -11748 6410 -11720
rect 4038 -13772 6326 -11748
rect 6390 -13772 6410 -11748
rect 4038 -13800 6410 -13772
rect -6410 -14068 -4038 -14040
rect -6410 -16092 -4122 -14068
rect -4058 -16092 -4038 -14068
rect -6410 -16120 -4038 -16092
rect -3798 -14068 -1426 -14040
rect -3798 -16092 -1510 -14068
rect -1446 -16092 -1426 -14068
rect -3798 -16120 -1426 -16092
rect -1186 -14068 1186 -14040
rect -1186 -16092 1102 -14068
rect 1166 -16092 1186 -14068
rect -1186 -16120 1186 -16092
rect 1426 -14068 3798 -14040
rect 1426 -16092 3714 -14068
rect 3778 -16092 3798 -14068
rect 1426 -16120 3798 -16092
rect 4038 -14068 6410 -14040
rect 4038 -16092 6326 -14068
rect 6390 -16092 6410 -14068
rect 4038 -16120 6410 -16092
rect -6410 -16388 -4038 -16360
rect -6410 -18412 -4122 -16388
rect -4058 -18412 -4038 -16388
rect -6410 -18440 -4038 -18412
rect -3798 -16388 -1426 -16360
rect -3798 -18412 -1510 -16388
rect -1446 -18412 -1426 -16388
rect -3798 -18440 -1426 -18412
rect -1186 -16388 1186 -16360
rect -1186 -18412 1102 -16388
rect 1166 -18412 1186 -16388
rect -1186 -18440 1186 -18412
rect 1426 -16388 3798 -16360
rect 1426 -18412 3714 -16388
rect 3778 -18412 3798 -16388
rect 1426 -18440 3798 -18412
rect 4038 -16388 6410 -16360
rect 4038 -18412 6326 -16388
rect 6390 -18412 6410 -16388
rect 4038 -18440 6410 -18412
rect -6410 -18708 -4038 -18680
rect -6410 -20732 -4122 -18708
rect -4058 -20732 -4038 -18708
rect -6410 -20760 -4038 -20732
rect -3798 -18708 -1426 -18680
rect -3798 -20732 -1510 -18708
rect -1446 -20732 -1426 -18708
rect -3798 -20760 -1426 -20732
rect -1186 -18708 1186 -18680
rect -1186 -20732 1102 -18708
rect 1166 -20732 1186 -18708
rect -1186 -20760 1186 -20732
rect 1426 -18708 3798 -18680
rect 1426 -20732 3714 -18708
rect 3778 -20732 3798 -18708
rect 1426 -20760 3798 -20732
rect 4038 -18708 6410 -18680
rect 4038 -20732 6326 -18708
rect 6390 -20732 6410 -18708
rect 4038 -20760 6410 -20732
rect -6410 -21028 -4038 -21000
rect -6410 -23052 -4122 -21028
rect -4058 -23052 -4038 -21028
rect -6410 -23080 -4038 -23052
rect -3798 -21028 -1426 -21000
rect -3798 -23052 -1510 -21028
rect -1446 -23052 -1426 -21028
rect -3798 -23080 -1426 -23052
rect -1186 -21028 1186 -21000
rect -1186 -23052 1102 -21028
rect 1166 -23052 1186 -21028
rect -1186 -23080 1186 -23052
rect 1426 -21028 3798 -21000
rect 1426 -23052 3714 -21028
rect 3778 -23052 3798 -21028
rect 1426 -23080 3798 -23052
rect 4038 -21028 6410 -21000
rect 4038 -23052 6326 -21028
rect 6390 -23052 6410 -21028
rect 4038 -23080 6410 -23052
rect -6410 -23348 -4038 -23320
rect -6410 -25372 -4122 -23348
rect -4058 -25372 -4038 -23348
rect -6410 -25400 -4038 -25372
rect -3798 -23348 -1426 -23320
rect -3798 -25372 -1510 -23348
rect -1446 -25372 -1426 -23348
rect -3798 -25400 -1426 -25372
rect -1186 -23348 1186 -23320
rect -1186 -25372 1102 -23348
rect 1166 -25372 1186 -23348
rect -1186 -25400 1186 -25372
rect 1426 -23348 3798 -23320
rect 1426 -25372 3714 -23348
rect 3778 -25372 3798 -23348
rect 1426 -25400 3798 -25372
rect 4038 -23348 6410 -23320
rect 4038 -25372 6326 -23348
rect 6390 -25372 6410 -23348
rect 4038 -25400 6410 -25372
rect -6410 -25668 -4038 -25640
rect -6410 -27692 -4122 -25668
rect -4058 -27692 -4038 -25668
rect -6410 -27720 -4038 -27692
rect -3798 -25668 -1426 -25640
rect -3798 -27692 -1510 -25668
rect -1446 -27692 -1426 -25668
rect -3798 -27720 -1426 -27692
rect -1186 -25668 1186 -25640
rect -1186 -27692 1102 -25668
rect 1166 -27692 1186 -25668
rect -1186 -27720 1186 -27692
rect 1426 -25668 3798 -25640
rect 1426 -27692 3714 -25668
rect 3778 -27692 3798 -25668
rect 1426 -27720 3798 -27692
rect 4038 -25668 6410 -25640
rect 4038 -27692 6326 -25668
rect 6390 -27692 6410 -25668
rect 4038 -27720 6410 -27692
rect -6410 -27988 -4038 -27960
rect -6410 -30012 -4122 -27988
rect -4058 -30012 -4038 -27988
rect -6410 -30040 -4038 -30012
rect -3798 -27988 -1426 -27960
rect -3798 -30012 -1510 -27988
rect -1446 -30012 -1426 -27988
rect -3798 -30040 -1426 -30012
rect -1186 -27988 1186 -27960
rect -1186 -30012 1102 -27988
rect 1166 -30012 1186 -27988
rect -1186 -30040 1186 -30012
rect 1426 -27988 3798 -27960
rect 1426 -30012 3714 -27988
rect 3778 -30012 3798 -27988
rect 1426 -30040 3798 -30012
rect 4038 -27988 6410 -27960
rect 4038 -30012 6326 -27988
rect 6390 -30012 6410 -27988
rect 4038 -30040 6410 -30012
rect -6410 -30308 -4038 -30280
rect -6410 -32332 -4122 -30308
rect -4058 -32332 -4038 -30308
rect -6410 -32360 -4038 -32332
rect -3798 -30308 -1426 -30280
rect -3798 -32332 -1510 -30308
rect -1446 -32332 -1426 -30308
rect -3798 -32360 -1426 -32332
rect -1186 -30308 1186 -30280
rect -1186 -32332 1102 -30308
rect 1166 -32332 1186 -30308
rect -1186 -32360 1186 -32332
rect 1426 -30308 3798 -30280
rect 1426 -32332 3714 -30308
rect 3778 -32332 3798 -30308
rect 1426 -32360 3798 -32332
rect 4038 -30308 6410 -30280
rect 4038 -32332 6326 -30308
rect 6390 -32332 6410 -30308
rect 4038 -32360 6410 -32332
rect -6410 -32628 -4038 -32600
rect -6410 -34652 -4122 -32628
rect -4058 -34652 -4038 -32628
rect -6410 -34680 -4038 -34652
rect -3798 -32628 -1426 -32600
rect -3798 -34652 -1510 -32628
rect -1446 -34652 -1426 -32628
rect -3798 -34680 -1426 -34652
rect -1186 -32628 1186 -32600
rect -1186 -34652 1102 -32628
rect 1166 -34652 1186 -32628
rect -1186 -34680 1186 -34652
rect 1426 -32628 3798 -32600
rect 1426 -34652 3714 -32628
rect 3778 -34652 3798 -32628
rect 1426 -34680 3798 -34652
rect 4038 -32628 6410 -32600
rect 4038 -34652 6326 -32628
rect 6390 -34652 6410 -32628
rect 4038 -34680 6410 -34652
rect -6410 -34948 -4038 -34920
rect -6410 -36972 -4122 -34948
rect -4058 -36972 -4038 -34948
rect -6410 -37000 -4038 -36972
rect -3798 -34948 -1426 -34920
rect -3798 -36972 -1510 -34948
rect -1446 -36972 -1426 -34948
rect -3798 -37000 -1426 -36972
rect -1186 -34948 1186 -34920
rect -1186 -36972 1102 -34948
rect 1166 -36972 1186 -34948
rect -1186 -37000 1186 -36972
rect 1426 -34948 3798 -34920
rect 1426 -36972 3714 -34948
rect 3778 -36972 3798 -34948
rect 1426 -37000 3798 -36972
rect 4038 -34948 6410 -34920
rect 4038 -36972 6326 -34948
rect 6390 -36972 6410 -34948
rect 4038 -37000 6410 -36972
<< via3 >>
rect -4122 34948 -4058 36972
rect -1510 34948 -1446 36972
rect 1102 34948 1166 36972
rect 3714 34948 3778 36972
rect 6326 34948 6390 36972
rect -4122 32628 -4058 34652
rect -1510 32628 -1446 34652
rect 1102 32628 1166 34652
rect 3714 32628 3778 34652
rect 6326 32628 6390 34652
rect -4122 30308 -4058 32332
rect -1510 30308 -1446 32332
rect 1102 30308 1166 32332
rect 3714 30308 3778 32332
rect 6326 30308 6390 32332
rect -4122 27988 -4058 30012
rect -1510 27988 -1446 30012
rect 1102 27988 1166 30012
rect 3714 27988 3778 30012
rect 6326 27988 6390 30012
rect -4122 25668 -4058 27692
rect -1510 25668 -1446 27692
rect 1102 25668 1166 27692
rect 3714 25668 3778 27692
rect 6326 25668 6390 27692
rect -4122 23348 -4058 25372
rect -1510 23348 -1446 25372
rect 1102 23348 1166 25372
rect 3714 23348 3778 25372
rect 6326 23348 6390 25372
rect -4122 21028 -4058 23052
rect -1510 21028 -1446 23052
rect 1102 21028 1166 23052
rect 3714 21028 3778 23052
rect 6326 21028 6390 23052
rect -4122 18708 -4058 20732
rect -1510 18708 -1446 20732
rect 1102 18708 1166 20732
rect 3714 18708 3778 20732
rect 6326 18708 6390 20732
rect -4122 16388 -4058 18412
rect -1510 16388 -1446 18412
rect 1102 16388 1166 18412
rect 3714 16388 3778 18412
rect 6326 16388 6390 18412
rect -4122 14068 -4058 16092
rect -1510 14068 -1446 16092
rect 1102 14068 1166 16092
rect 3714 14068 3778 16092
rect 6326 14068 6390 16092
rect -4122 11748 -4058 13772
rect -1510 11748 -1446 13772
rect 1102 11748 1166 13772
rect 3714 11748 3778 13772
rect 6326 11748 6390 13772
rect -4122 9428 -4058 11452
rect -1510 9428 -1446 11452
rect 1102 9428 1166 11452
rect 3714 9428 3778 11452
rect 6326 9428 6390 11452
rect -4122 7108 -4058 9132
rect -1510 7108 -1446 9132
rect 1102 7108 1166 9132
rect 3714 7108 3778 9132
rect 6326 7108 6390 9132
rect -4122 4788 -4058 6812
rect -1510 4788 -1446 6812
rect 1102 4788 1166 6812
rect 3714 4788 3778 6812
rect 6326 4788 6390 6812
rect -4122 2468 -4058 4492
rect -1510 2468 -1446 4492
rect 1102 2468 1166 4492
rect 3714 2468 3778 4492
rect 6326 2468 6390 4492
rect -4122 148 -4058 2172
rect -1510 148 -1446 2172
rect 1102 148 1166 2172
rect 3714 148 3778 2172
rect 6326 148 6390 2172
rect -4122 -2172 -4058 -148
rect -1510 -2172 -1446 -148
rect 1102 -2172 1166 -148
rect 3714 -2172 3778 -148
rect 6326 -2172 6390 -148
rect -4122 -4492 -4058 -2468
rect -1510 -4492 -1446 -2468
rect 1102 -4492 1166 -2468
rect 3714 -4492 3778 -2468
rect 6326 -4492 6390 -2468
rect -4122 -6812 -4058 -4788
rect -1510 -6812 -1446 -4788
rect 1102 -6812 1166 -4788
rect 3714 -6812 3778 -4788
rect 6326 -6812 6390 -4788
rect -4122 -9132 -4058 -7108
rect -1510 -9132 -1446 -7108
rect 1102 -9132 1166 -7108
rect 3714 -9132 3778 -7108
rect 6326 -9132 6390 -7108
rect -4122 -11452 -4058 -9428
rect -1510 -11452 -1446 -9428
rect 1102 -11452 1166 -9428
rect 3714 -11452 3778 -9428
rect 6326 -11452 6390 -9428
rect -4122 -13772 -4058 -11748
rect -1510 -13772 -1446 -11748
rect 1102 -13772 1166 -11748
rect 3714 -13772 3778 -11748
rect 6326 -13772 6390 -11748
rect -4122 -16092 -4058 -14068
rect -1510 -16092 -1446 -14068
rect 1102 -16092 1166 -14068
rect 3714 -16092 3778 -14068
rect 6326 -16092 6390 -14068
rect -4122 -18412 -4058 -16388
rect -1510 -18412 -1446 -16388
rect 1102 -18412 1166 -16388
rect 3714 -18412 3778 -16388
rect 6326 -18412 6390 -16388
rect -4122 -20732 -4058 -18708
rect -1510 -20732 -1446 -18708
rect 1102 -20732 1166 -18708
rect 3714 -20732 3778 -18708
rect 6326 -20732 6390 -18708
rect -4122 -23052 -4058 -21028
rect -1510 -23052 -1446 -21028
rect 1102 -23052 1166 -21028
rect 3714 -23052 3778 -21028
rect 6326 -23052 6390 -21028
rect -4122 -25372 -4058 -23348
rect -1510 -25372 -1446 -23348
rect 1102 -25372 1166 -23348
rect 3714 -25372 3778 -23348
rect 6326 -25372 6390 -23348
rect -4122 -27692 -4058 -25668
rect -1510 -27692 -1446 -25668
rect 1102 -27692 1166 -25668
rect 3714 -27692 3778 -25668
rect 6326 -27692 6390 -25668
rect -4122 -30012 -4058 -27988
rect -1510 -30012 -1446 -27988
rect 1102 -30012 1166 -27988
rect 3714 -30012 3778 -27988
rect 6326 -30012 6390 -27988
rect -4122 -32332 -4058 -30308
rect -1510 -32332 -1446 -30308
rect 1102 -32332 1166 -30308
rect 3714 -32332 3778 -30308
rect 6326 -32332 6390 -30308
rect -4122 -34652 -4058 -32628
rect -1510 -34652 -1446 -32628
rect 1102 -34652 1166 -32628
rect 3714 -34652 3778 -32628
rect 6326 -34652 6390 -32628
rect -4122 -36972 -4058 -34948
rect -1510 -36972 -1446 -34948
rect 1102 -36972 1166 -34948
rect 3714 -36972 3778 -34948
rect 6326 -36972 6390 -34948
<< mimcap >>
rect -6370 36920 -4370 36960
rect -6370 35000 -6330 36920
rect -4410 35000 -4370 36920
rect -6370 34960 -4370 35000
rect -3758 36920 -1758 36960
rect -3758 35000 -3718 36920
rect -1798 35000 -1758 36920
rect -3758 34960 -1758 35000
rect -1146 36920 854 36960
rect -1146 35000 -1106 36920
rect 814 35000 854 36920
rect -1146 34960 854 35000
rect 1466 36920 3466 36960
rect 1466 35000 1506 36920
rect 3426 35000 3466 36920
rect 1466 34960 3466 35000
rect 4078 36920 6078 36960
rect 4078 35000 4118 36920
rect 6038 35000 6078 36920
rect 4078 34960 6078 35000
rect -6370 34600 -4370 34640
rect -6370 32680 -6330 34600
rect -4410 32680 -4370 34600
rect -6370 32640 -4370 32680
rect -3758 34600 -1758 34640
rect -3758 32680 -3718 34600
rect -1798 32680 -1758 34600
rect -3758 32640 -1758 32680
rect -1146 34600 854 34640
rect -1146 32680 -1106 34600
rect 814 32680 854 34600
rect -1146 32640 854 32680
rect 1466 34600 3466 34640
rect 1466 32680 1506 34600
rect 3426 32680 3466 34600
rect 1466 32640 3466 32680
rect 4078 34600 6078 34640
rect 4078 32680 4118 34600
rect 6038 32680 6078 34600
rect 4078 32640 6078 32680
rect -6370 32280 -4370 32320
rect -6370 30360 -6330 32280
rect -4410 30360 -4370 32280
rect -6370 30320 -4370 30360
rect -3758 32280 -1758 32320
rect -3758 30360 -3718 32280
rect -1798 30360 -1758 32280
rect -3758 30320 -1758 30360
rect -1146 32280 854 32320
rect -1146 30360 -1106 32280
rect 814 30360 854 32280
rect -1146 30320 854 30360
rect 1466 32280 3466 32320
rect 1466 30360 1506 32280
rect 3426 30360 3466 32280
rect 1466 30320 3466 30360
rect 4078 32280 6078 32320
rect 4078 30360 4118 32280
rect 6038 30360 6078 32280
rect 4078 30320 6078 30360
rect -6370 29960 -4370 30000
rect -6370 28040 -6330 29960
rect -4410 28040 -4370 29960
rect -6370 28000 -4370 28040
rect -3758 29960 -1758 30000
rect -3758 28040 -3718 29960
rect -1798 28040 -1758 29960
rect -3758 28000 -1758 28040
rect -1146 29960 854 30000
rect -1146 28040 -1106 29960
rect 814 28040 854 29960
rect -1146 28000 854 28040
rect 1466 29960 3466 30000
rect 1466 28040 1506 29960
rect 3426 28040 3466 29960
rect 1466 28000 3466 28040
rect 4078 29960 6078 30000
rect 4078 28040 4118 29960
rect 6038 28040 6078 29960
rect 4078 28000 6078 28040
rect -6370 27640 -4370 27680
rect -6370 25720 -6330 27640
rect -4410 25720 -4370 27640
rect -6370 25680 -4370 25720
rect -3758 27640 -1758 27680
rect -3758 25720 -3718 27640
rect -1798 25720 -1758 27640
rect -3758 25680 -1758 25720
rect -1146 27640 854 27680
rect -1146 25720 -1106 27640
rect 814 25720 854 27640
rect -1146 25680 854 25720
rect 1466 27640 3466 27680
rect 1466 25720 1506 27640
rect 3426 25720 3466 27640
rect 1466 25680 3466 25720
rect 4078 27640 6078 27680
rect 4078 25720 4118 27640
rect 6038 25720 6078 27640
rect 4078 25680 6078 25720
rect -6370 25320 -4370 25360
rect -6370 23400 -6330 25320
rect -4410 23400 -4370 25320
rect -6370 23360 -4370 23400
rect -3758 25320 -1758 25360
rect -3758 23400 -3718 25320
rect -1798 23400 -1758 25320
rect -3758 23360 -1758 23400
rect -1146 25320 854 25360
rect -1146 23400 -1106 25320
rect 814 23400 854 25320
rect -1146 23360 854 23400
rect 1466 25320 3466 25360
rect 1466 23400 1506 25320
rect 3426 23400 3466 25320
rect 1466 23360 3466 23400
rect 4078 25320 6078 25360
rect 4078 23400 4118 25320
rect 6038 23400 6078 25320
rect 4078 23360 6078 23400
rect -6370 23000 -4370 23040
rect -6370 21080 -6330 23000
rect -4410 21080 -4370 23000
rect -6370 21040 -4370 21080
rect -3758 23000 -1758 23040
rect -3758 21080 -3718 23000
rect -1798 21080 -1758 23000
rect -3758 21040 -1758 21080
rect -1146 23000 854 23040
rect -1146 21080 -1106 23000
rect 814 21080 854 23000
rect -1146 21040 854 21080
rect 1466 23000 3466 23040
rect 1466 21080 1506 23000
rect 3426 21080 3466 23000
rect 1466 21040 3466 21080
rect 4078 23000 6078 23040
rect 4078 21080 4118 23000
rect 6038 21080 6078 23000
rect 4078 21040 6078 21080
rect -6370 20680 -4370 20720
rect -6370 18760 -6330 20680
rect -4410 18760 -4370 20680
rect -6370 18720 -4370 18760
rect -3758 20680 -1758 20720
rect -3758 18760 -3718 20680
rect -1798 18760 -1758 20680
rect -3758 18720 -1758 18760
rect -1146 20680 854 20720
rect -1146 18760 -1106 20680
rect 814 18760 854 20680
rect -1146 18720 854 18760
rect 1466 20680 3466 20720
rect 1466 18760 1506 20680
rect 3426 18760 3466 20680
rect 1466 18720 3466 18760
rect 4078 20680 6078 20720
rect 4078 18760 4118 20680
rect 6038 18760 6078 20680
rect 4078 18720 6078 18760
rect -6370 18360 -4370 18400
rect -6370 16440 -6330 18360
rect -4410 16440 -4370 18360
rect -6370 16400 -4370 16440
rect -3758 18360 -1758 18400
rect -3758 16440 -3718 18360
rect -1798 16440 -1758 18360
rect -3758 16400 -1758 16440
rect -1146 18360 854 18400
rect -1146 16440 -1106 18360
rect 814 16440 854 18360
rect -1146 16400 854 16440
rect 1466 18360 3466 18400
rect 1466 16440 1506 18360
rect 3426 16440 3466 18360
rect 1466 16400 3466 16440
rect 4078 18360 6078 18400
rect 4078 16440 4118 18360
rect 6038 16440 6078 18360
rect 4078 16400 6078 16440
rect -6370 16040 -4370 16080
rect -6370 14120 -6330 16040
rect -4410 14120 -4370 16040
rect -6370 14080 -4370 14120
rect -3758 16040 -1758 16080
rect -3758 14120 -3718 16040
rect -1798 14120 -1758 16040
rect -3758 14080 -1758 14120
rect -1146 16040 854 16080
rect -1146 14120 -1106 16040
rect 814 14120 854 16040
rect -1146 14080 854 14120
rect 1466 16040 3466 16080
rect 1466 14120 1506 16040
rect 3426 14120 3466 16040
rect 1466 14080 3466 14120
rect 4078 16040 6078 16080
rect 4078 14120 4118 16040
rect 6038 14120 6078 16040
rect 4078 14080 6078 14120
rect -6370 13720 -4370 13760
rect -6370 11800 -6330 13720
rect -4410 11800 -4370 13720
rect -6370 11760 -4370 11800
rect -3758 13720 -1758 13760
rect -3758 11800 -3718 13720
rect -1798 11800 -1758 13720
rect -3758 11760 -1758 11800
rect -1146 13720 854 13760
rect -1146 11800 -1106 13720
rect 814 11800 854 13720
rect -1146 11760 854 11800
rect 1466 13720 3466 13760
rect 1466 11800 1506 13720
rect 3426 11800 3466 13720
rect 1466 11760 3466 11800
rect 4078 13720 6078 13760
rect 4078 11800 4118 13720
rect 6038 11800 6078 13720
rect 4078 11760 6078 11800
rect -6370 11400 -4370 11440
rect -6370 9480 -6330 11400
rect -4410 9480 -4370 11400
rect -6370 9440 -4370 9480
rect -3758 11400 -1758 11440
rect -3758 9480 -3718 11400
rect -1798 9480 -1758 11400
rect -3758 9440 -1758 9480
rect -1146 11400 854 11440
rect -1146 9480 -1106 11400
rect 814 9480 854 11400
rect -1146 9440 854 9480
rect 1466 11400 3466 11440
rect 1466 9480 1506 11400
rect 3426 9480 3466 11400
rect 1466 9440 3466 9480
rect 4078 11400 6078 11440
rect 4078 9480 4118 11400
rect 6038 9480 6078 11400
rect 4078 9440 6078 9480
rect -6370 9080 -4370 9120
rect -6370 7160 -6330 9080
rect -4410 7160 -4370 9080
rect -6370 7120 -4370 7160
rect -3758 9080 -1758 9120
rect -3758 7160 -3718 9080
rect -1798 7160 -1758 9080
rect -3758 7120 -1758 7160
rect -1146 9080 854 9120
rect -1146 7160 -1106 9080
rect 814 7160 854 9080
rect -1146 7120 854 7160
rect 1466 9080 3466 9120
rect 1466 7160 1506 9080
rect 3426 7160 3466 9080
rect 1466 7120 3466 7160
rect 4078 9080 6078 9120
rect 4078 7160 4118 9080
rect 6038 7160 6078 9080
rect 4078 7120 6078 7160
rect -6370 6760 -4370 6800
rect -6370 4840 -6330 6760
rect -4410 4840 -4370 6760
rect -6370 4800 -4370 4840
rect -3758 6760 -1758 6800
rect -3758 4840 -3718 6760
rect -1798 4840 -1758 6760
rect -3758 4800 -1758 4840
rect -1146 6760 854 6800
rect -1146 4840 -1106 6760
rect 814 4840 854 6760
rect -1146 4800 854 4840
rect 1466 6760 3466 6800
rect 1466 4840 1506 6760
rect 3426 4840 3466 6760
rect 1466 4800 3466 4840
rect 4078 6760 6078 6800
rect 4078 4840 4118 6760
rect 6038 4840 6078 6760
rect 4078 4800 6078 4840
rect -6370 4440 -4370 4480
rect -6370 2520 -6330 4440
rect -4410 2520 -4370 4440
rect -6370 2480 -4370 2520
rect -3758 4440 -1758 4480
rect -3758 2520 -3718 4440
rect -1798 2520 -1758 4440
rect -3758 2480 -1758 2520
rect -1146 4440 854 4480
rect -1146 2520 -1106 4440
rect 814 2520 854 4440
rect -1146 2480 854 2520
rect 1466 4440 3466 4480
rect 1466 2520 1506 4440
rect 3426 2520 3466 4440
rect 1466 2480 3466 2520
rect 4078 4440 6078 4480
rect 4078 2520 4118 4440
rect 6038 2520 6078 4440
rect 4078 2480 6078 2520
rect -6370 2120 -4370 2160
rect -6370 200 -6330 2120
rect -4410 200 -4370 2120
rect -6370 160 -4370 200
rect -3758 2120 -1758 2160
rect -3758 200 -3718 2120
rect -1798 200 -1758 2120
rect -3758 160 -1758 200
rect -1146 2120 854 2160
rect -1146 200 -1106 2120
rect 814 200 854 2120
rect -1146 160 854 200
rect 1466 2120 3466 2160
rect 1466 200 1506 2120
rect 3426 200 3466 2120
rect 1466 160 3466 200
rect 4078 2120 6078 2160
rect 4078 200 4118 2120
rect 6038 200 6078 2120
rect 4078 160 6078 200
rect -6370 -200 -4370 -160
rect -6370 -2120 -6330 -200
rect -4410 -2120 -4370 -200
rect -6370 -2160 -4370 -2120
rect -3758 -200 -1758 -160
rect -3758 -2120 -3718 -200
rect -1798 -2120 -1758 -200
rect -3758 -2160 -1758 -2120
rect -1146 -200 854 -160
rect -1146 -2120 -1106 -200
rect 814 -2120 854 -200
rect -1146 -2160 854 -2120
rect 1466 -200 3466 -160
rect 1466 -2120 1506 -200
rect 3426 -2120 3466 -200
rect 1466 -2160 3466 -2120
rect 4078 -200 6078 -160
rect 4078 -2120 4118 -200
rect 6038 -2120 6078 -200
rect 4078 -2160 6078 -2120
rect -6370 -2520 -4370 -2480
rect -6370 -4440 -6330 -2520
rect -4410 -4440 -4370 -2520
rect -6370 -4480 -4370 -4440
rect -3758 -2520 -1758 -2480
rect -3758 -4440 -3718 -2520
rect -1798 -4440 -1758 -2520
rect -3758 -4480 -1758 -4440
rect -1146 -2520 854 -2480
rect -1146 -4440 -1106 -2520
rect 814 -4440 854 -2520
rect -1146 -4480 854 -4440
rect 1466 -2520 3466 -2480
rect 1466 -4440 1506 -2520
rect 3426 -4440 3466 -2520
rect 1466 -4480 3466 -4440
rect 4078 -2520 6078 -2480
rect 4078 -4440 4118 -2520
rect 6038 -4440 6078 -2520
rect 4078 -4480 6078 -4440
rect -6370 -4840 -4370 -4800
rect -6370 -6760 -6330 -4840
rect -4410 -6760 -4370 -4840
rect -6370 -6800 -4370 -6760
rect -3758 -4840 -1758 -4800
rect -3758 -6760 -3718 -4840
rect -1798 -6760 -1758 -4840
rect -3758 -6800 -1758 -6760
rect -1146 -4840 854 -4800
rect -1146 -6760 -1106 -4840
rect 814 -6760 854 -4840
rect -1146 -6800 854 -6760
rect 1466 -4840 3466 -4800
rect 1466 -6760 1506 -4840
rect 3426 -6760 3466 -4840
rect 1466 -6800 3466 -6760
rect 4078 -4840 6078 -4800
rect 4078 -6760 4118 -4840
rect 6038 -6760 6078 -4840
rect 4078 -6800 6078 -6760
rect -6370 -7160 -4370 -7120
rect -6370 -9080 -6330 -7160
rect -4410 -9080 -4370 -7160
rect -6370 -9120 -4370 -9080
rect -3758 -7160 -1758 -7120
rect -3758 -9080 -3718 -7160
rect -1798 -9080 -1758 -7160
rect -3758 -9120 -1758 -9080
rect -1146 -7160 854 -7120
rect -1146 -9080 -1106 -7160
rect 814 -9080 854 -7160
rect -1146 -9120 854 -9080
rect 1466 -7160 3466 -7120
rect 1466 -9080 1506 -7160
rect 3426 -9080 3466 -7160
rect 1466 -9120 3466 -9080
rect 4078 -7160 6078 -7120
rect 4078 -9080 4118 -7160
rect 6038 -9080 6078 -7160
rect 4078 -9120 6078 -9080
rect -6370 -9480 -4370 -9440
rect -6370 -11400 -6330 -9480
rect -4410 -11400 -4370 -9480
rect -6370 -11440 -4370 -11400
rect -3758 -9480 -1758 -9440
rect -3758 -11400 -3718 -9480
rect -1798 -11400 -1758 -9480
rect -3758 -11440 -1758 -11400
rect -1146 -9480 854 -9440
rect -1146 -11400 -1106 -9480
rect 814 -11400 854 -9480
rect -1146 -11440 854 -11400
rect 1466 -9480 3466 -9440
rect 1466 -11400 1506 -9480
rect 3426 -11400 3466 -9480
rect 1466 -11440 3466 -11400
rect 4078 -9480 6078 -9440
rect 4078 -11400 4118 -9480
rect 6038 -11400 6078 -9480
rect 4078 -11440 6078 -11400
rect -6370 -11800 -4370 -11760
rect -6370 -13720 -6330 -11800
rect -4410 -13720 -4370 -11800
rect -6370 -13760 -4370 -13720
rect -3758 -11800 -1758 -11760
rect -3758 -13720 -3718 -11800
rect -1798 -13720 -1758 -11800
rect -3758 -13760 -1758 -13720
rect -1146 -11800 854 -11760
rect -1146 -13720 -1106 -11800
rect 814 -13720 854 -11800
rect -1146 -13760 854 -13720
rect 1466 -11800 3466 -11760
rect 1466 -13720 1506 -11800
rect 3426 -13720 3466 -11800
rect 1466 -13760 3466 -13720
rect 4078 -11800 6078 -11760
rect 4078 -13720 4118 -11800
rect 6038 -13720 6078 -11800
rect 4078 -13760 6078 -13720
rect -6370 -14120 -4370 -14080
rect -6370 -16040 -6330 -14120
rect -4410 -16040 -4370 -14120
rect -6370 -16080 -4370 -16040
rect -3758 -14120 -1758 -14080
rect -3758 -16040 -3718 -14120
rect -1798 -16040 -1758 -14120
rect -3758 -16080 -1758 -16040
rect -1146 -14120 854 -14080
rect -1146 -16040 -1106 -14120
rect 814 -16040 854 -14120
rect -1146 -16080 854 -16040
rect 1466 -14120 3466 -14080
rect 1466 -16040 1506 -14120
rect 3426 -16040 3466 -14120
rect 1466 -16080 3466 -16040
rect 4078 -14120 6078 -14080
rect 4078 -16040 4118 -14120
rect 6038 -16040 6078 -14120
rect 4078 -16080 6078 -16040
rect -6370 -16440 -4370 -16400
rect -6370 -18360 -6330 -16440
rect -4410 -18360 -4370 -16440
rect -6370 -18400 -4370 -18360
rect -3758 -16440 -1758 -16400
rect -3758 -18360 -3718 -16440
rect -1798 -18360 -1758 -16440
rect -3758 -18400 -1758 -18360
rect -1146 -16440 854 -16400
rect -1146 -18360 -1106 -16440
rect 814 -18360 854 -16440
rect -1146 -18400 854 -18360
rect 1466 -16440 3466 -16400
rect 1466 -18360 1506 -16440
rect 3426 -18360 3466 -16440
rect 1466 -18400 3466 -18360
rect 4078 -16440 6078 -16400
rect 4078 -18360 4118 -16440
rect 6038 -18360 6078 -16440
rect 4078 -18400 6078 -18360
rect -6370 -18760 -4370 -18720
rect -6370 -20680 -6330 -18760
rect -4410 -20680 -4370 -18760
rect -6370 -20720 -4370 -20680
rect -3758 -18760 -1758 -18720
rect -3758 -20680 -3718 -18760
rect -1798 -20680 -1758 -18760
rect -3758 -20720 -1758 -20680
rect -1146 -18760 854 -18720
rect -1146 -20680 -1106 -18760
rect 814 -20680 854 -18760
rect -1146 -20720 854 -20680
rect 1466 -18760 3466 -18720
rect 1466 -20680 1506 -18760
rect 3426 -20680 3466 -18760
rect 1466 -20720 3466 -20680
rect 4078 -18760 6078 -18720
rect 4078 -20680 4118 -18760
rect 6038 -20680 6078 -18760
rect 4078 -20720 6078 -20680
rect -6370 -21080 -4370 -21040
rect -6370 -23000 -6330 -21080
rect -4410 -23000 -4370 -21080
rect -6370 -23040 -4370 -23000
rect -3758 -21080 -1758 -21040
rect -3758 -23000 -3718 -21080
rect -1798 -23000 -1758 -21080
rect -3758 -23040 -1758 -23000
rect -1146 -21080 854 -21040
rect -1146 -23000 -1106 -21080
rect 814 -23000 854 -21080
rect -1146 -23040 854 -23000
rect 1466 -21080 3466 -21040
rect 1466 -23000 1506 -21080
rect 3426 -23000 3466 -21080
rect 1466 -23040 3466 -23000
rect 4078 -21080 6078 -21040
rect 4078 -23000 4118 -21080
rect 6038 -23000 6078 -21080
rect 4078 -23040 6078 -23000
rect -6370 -23400 -4370 -23360
rect -6370 -25320 -6330 -23400
rect -4410 -25320 -4370 -23400
rect -6370 -25360 -4370 -25320
rect -3758 -23400 -1758 -23360
rect -3758 -25320 -3718 -23400
rect -1798 -25320 -1758 -23400
rect -3758 -25360 -1758 -25320
rect -1146 -23400 854 -23360
rect -1146 -25320 -1106 -23400
rect 814 -25320 854 -23400
rect -1146 -25360 854 -25320
rect 1466 -23400 3466 -23360
rect 1466 -25320 1506 -23400
rect 3426 -25320 3466 -23400
rect 1466 -25360 3466 -25320
rect 4078 -23400 6078 -23360
rect 4078 -25320 4118 -23400
rect 6038 -25320 6078 -23400
rect 4078 -25360 6078 -25320
rect -6370 -25720 -4370 -25680
rect -6370 -27640 -6330 -25720
rect -4410 -27640 -4370 -25720
rect -6370 -27680 -4370 -27640
rect -3758 -25720 -1758 -25680
rect -3758 -27640 -3718 -25720
rect -1798 -27640 -1758 -25720
rect -3758 -27680 -1758 -27640
rect -1146 -25720 854 -25680
rect -1146 -27640 -1106 -25720
rect 814 -27640 854 -25720
rect -1146 -27680 854 -27640
rect 1466 -25720 3466 -25680
rect 1466 -27640 1506 -25720
rect 3426 -27640 3466 -25720
rect 1466 -27680 3466 -27640
rect 4078 -25720 6078 -25680
rect 4078 -27640 4118 -25720
rect 6038 -27640 6078 -25720
rect 4078 -27680 6078 -27640
rect -6370 -28040 -4370 -28000
rect -6370 -29960 -6330 -28040
rect -4410 -29960 -4370 -28040
rect -6370 -30000 -4370 -29960
rect -3758 -28040 -1758 -28000
rect -3758 -29960 -3718 -28040
rect -1798 -29960 -1758 -28040
rect -3758 -30000 -1758 -29960
rect -1146 -28040 854 -28000
rect -1146 -29960 -1106 -28040
rect 814 -29960 854 -28040
rect -1146 -30000 854 -29960
rect 1466 -28040 3466 -28000
rect 1466 -29960 1506 -28040
rect 3426 -29960 3466 -28040
rect 1466 -30000 3466 -29960
rect 4078 -28040 6078 -28000
rect 4078 -29960 4118 -28040
rect 6038 -29960 6078 -28040
rect 4078 -30000 6078 -29960
rect -6370 -30360 -4370 -30320
rect -6370 -32280 -6330 -30360
rect -4410 -32280 -4370 -30360
rect -6370 -32320 -4370 -32280
rect -3758 -30360 -1758 -30320
rect -3758 -32280 -3718 -30360
rect -1798 -32280 -1758 -30360
rect -3758 -32320 -1758 -32280
rect -1146 -30360 854 -30320
rect -1146 -32280 -1106 -30360
rect 814 -32280 854 -30360
rect -1146 -32320 854 -32280
rect 1466 -30360 3466 -30320
rect 1466 -32280 1506 -30360
rect 3426 -32280 3466 -30360
rect 1466 -32320 3466 -32280
rect 4078 -30360 6078 -30320
rect 4078 -32280 4118 -30360
rect 6038 -32280 6078 -30360
rect 4078 -32320 6078 -32280
rect -6370 -32680 -4370 -32640
rect -6370 -34600 -6330 -32680
rect -4410 -34600 -4370 -32680
rect -6370 -34640 -4370 -34600
rect -3758 -32680 -1758 -32640
rect -3758 -34600 -3718 -32680
rect -1798 -34600 -1758 -32680
rect -3758 -34640 -1758 -34600
rect -1146 -32680 854 -32640
rect -1146 -34600 -1106 -32680
rect 814 -34600 854 -32680
rect -1146 -34640 854 -34600
rect 1466 -32680 3466 -32640
rect 1466 -34600 1506 -32680
rect 3426 -34600 3466 -32680
rect 1466 -34640 3466 -34600
rect 4078 -32680 6078 -32640
rect 4078 -34600 4118 -32680
rect 6038 -34600 6078 -32680
rect 4078 -34640 6078 -34600
rect -6370 -35000 -4370 -34960
rect -6370 -36920 -6330 -35000
rect -4410 -36920 -4370 -35000
rect -6370 -36960 -4370 -36920
rect -3758 -35000 -1758 -34960
rect -3758 -36920 -3718 -35000
rect -1798 -36920 -1758 -35000
rect -3758 -36960 -1758 -36920
rect -1146 -35000 854 -34960
rect -1146 -36920 -1106 -35000
rect 814 -36920 854 -35000
rect -1146 -36960 854 -36920
rect 1466 -35000 3466 -34960
rect 1466 -36920 1506 -35000
rect 3426 -36920 3466 -35000
rect 1466 -36960 3466 -36920
rect 4078 -35000 6078 -34960
rect 4078 -36920 4118 -35000
rect 6038 -36920 6078 -35000
rect 4078 -36960 6078 -36920
<< mimcapcontact >>
rect -6330 35000 -4410 36920
rect -3718 35000 -1798 36920
rect -1106 35000 814 36920
rect 1506 35000 3426 36920
rect 4118 35000 6038 36920
rect -6330 32680 -4410 34600
rect -3718 32680 -1798 34600
rect -1106 32680 814 34600
rect 1506 32680 3426 34600
rect 4118 32680 6038 34600
rect -6330 30360 -4410 32280
rect -3718 30360 -1798 32280
rect -1106 30360 814 32280
rect 1506 30360 3426 32280
rect 4118 30360 6038 32280
rect -6330 28040 -4410 29960
rect -3718 28040 -1798 29960
rect -1106 28040 814 29960
rect 1506 28040 3426 29960
rect 4118 28040 6038 29960
rect -6330 25720 -4410 27640
rect -3718 25720 -1798 27640
rect -1106 25720 814 27640
rect 1506 25720 3426 27640
rect 4118 25720 6038 27640
rect -6330 23400 -4410 25320
rect -3718 23400 -1798 25320
rect -1106 23400 814 25320
rect 1506 23400 3426 25320
rect 4118 23400 6038 25320
rect -6330 21080 -4410 23000
rect -3718 21080 -1798 23000
rect -1106 21080 814 23000
rect 1506 21080 3426 23000
rect 4118 21080 6038 23000
rect -6330 18760 -4410 20680
rect -3718 18760 -1798 20680
rect -1106 18760 814 20680
rect 1506 18760 3426 20680
rect 4118 18760 6038 20680
rect -6330 16440 -4410 18360
rect -3718 16440 -1798 18360
rect -1106 16440 814 18360
rect 1506 16440 3426 18360
rect 4118 16440 6038 18360
rect -6330 14120 -4410 16040
rect -3718 14120 -1798 16040
rect -1106 14120 814 16040
rect 1506 14120 3426 16040
rect 4118 14120 6038 16040
rect -6330 11800 -4410 13720
rect -3718 11800 -1798 13720
rect -1106 11800 814 13720
rect 1506 11800 3426 13720
rect 4118 11800 6038 13720
rect -6330 9480 -4410 11400
rect -3718 9480 -1798 11400
rect -1106 9480 814 11400
rect 1506 9480 3426 11400
rect 4118 9480 6038 11400
rect -6330 7160 -4410 9080
rect -3718 7160 -1798 9080
rect -1106 7160 814 9080
rect 1506 7160 3426 9080
rect 4118 7160 6038 9080
rect -6330 4840 -4410 6760
rect -3718 4840 -1798 6760
rect -1106 4840 814 6760
rect 1506 4840 3426 6760
rect 4118 4840 6038 6760
rect -6330 2520 -4410 4440
rect -3718 2520 -1798 4440
rect -1106 2520 814 4440
rect 1506 2520 3426 4440
rect 4118 2520 6038 4440
rect -6330 200 -4410 2120
rect -3718 200 -1798 2120
rect -1106 200 814 2120
rect 1506 200 3426 2120
rect 4118 200 6038 2120
rect -6330 -2120 -4410 -200
rect -3718 -2120 -1798 -200
rect -1106 -2120 814 -200
rect 1506 -2120 3426 -200
rect 4118 -2120 6038 -200
rect -6330 -4440 -4410 -2520
rect -3718 -4440 -1798 -2520
rect -1106 -4440 814 -2520
rect 1506 -4440 3426 -2520
rect 4118 -4440 6038 -2520
rect -6330 -6760 -4410 -4840
rect -3718 -6760 -1798 -4840
rect -1106 -6760 814 -4840
rect 1506 -6760 3426 -4840
rect 4118 -6760 6038 -4840
rect -6330 -9080 -4410 -7160
rect -3718 -9080 -1798 -7160
rect -1106 -9080 814 -7160
rect 1506 -9080 3426 -7160
rect 4118 -9080 6038 -7160
rect -6330 -11400 -4410 -9480
rect -3718 -11400 -1798 -9480
rect -1106 -11400 814 -9480
rect 1506 -11400 3426 -9480
rect 4118 -11400 6038 -9480
rect -6330 -13720 -4410 -11800
rect -3718 -13720 -1798 -11800
rect -1106 -13720 814 -11800
rect 1506 -13720 3426 -11800
rect 4118 -13720 6038 -11800
rect -6330 -16040 -4410 -14120
rect -3718 -16040 -1798 -14120
rect -1106 -16040 814 -14120
rect 1506 -16040 3426 -14120
rect 4118 -16040 6038 -14120
rect -6330 -18360 -4410 -16440
rect -3718 -18360 -1798 -16440
rect -1106 -18360 814 -16440
rect 1506 -18360 3426 -16440
rect 4118 -18360 6038 -16440
rect -6330 -20680 -4410 -18760
rect -3718 -20680 -1798 -18760
rect -1106 -20680 814 -18760
rect 1506 -20680 3426 -18760
rect 4118 -20680 6038 -18760
rect -6330 -23000 -4410 -21080
rect -3718 -23000 -1798 -21080
rect -1106 -23000 814 -21080
rect 1506 -23000 3426 -21080
rect 4118 -23000 6038 -21080
rect -6330 -25320 -4410 -23400
rect -3718 -25320 -1798 -23400
rect -1106 -25320 814 -23400
rect 1506 -25320 3426 -23400
rect 4118 -25320 6038 -23400
rect -6330 -27640 -4410 -25720
rect -3718 -27640 -1798 -25720
rect -1106 -27640 814 -25720
rect 1506 -27640 3426 -25720
rect 4118 -27640 6038 -25720
rect -6330 -29960 -4410 -28040
rect -3718 -29960 -1798 -28040
rect -1106 -29960 814 -28040
rect 1506 -29960 3426 -28040
rect 4118 -29960 6038 -28040
rect -6330 -32280 -4410 -30360
rect -3718 -32280 -1798 -30360
rect -1106 -32280 814 -30360
rect 1506 -32280 3426 -30360
rect 4118 -32280 6038 -30360
rect -6330 -34600 -4410 -32680
rect -3718 -34600 -1798 -32680
rect -1106 -34600 814 -32680
rect 1506 -34600 3426 -32680
rect 4118 -34600 6038 -32680
rect -6330 -36920 -4410 -35000
rect -3718 -36920 -1798 -35000
rect -1106 -36920 814 -35000
rect 1506 -36920 3426 -35000
rect 4118 -36920 6038 -35000
<< metal4 >>
rect -5422 36921 -5318 37120
rect -4142 36972 -4038 37120
rect -6331 36920 -4409 36921
rect -6331 35000 -6330 36920
rect -4410 35000 -4409 36920
rect -6331 34999 -4409 35000
rect -5422 34601 -5318 34999
rect -4142 34948 -4122 36972
rect -4058 34948 -4038 36972
rect -2810 36921 -2706 37120
rect -1530 36972 -1426 37120
rect -3719 36920 -1797 36921
rect -3719 35000 -3718 36920
rect -1798 35000 -1797 36920
rect -3719 34999 -1797 35000
rect -4142 34652 -4038 34948
rect -6331 34600 -4409 34601
rect -6331 32680 -6330 34600
rect -4410 32680 -4409 34600
rect -6331 32679 -4409 32680
rect -5422 32281 -5318 32679
rect -4142 32628 -4122 34652
rect -4058 32628 -4038 34652
rect -2810 34601 -2706 34999
rect -1530 34948 -1510 36972
rect -1446 34948 -1426 36972
rect -198 36921 -94 37120
rect 1082 36972 1186 37120
rect -1107 36920 815 36921
rect -1107 35000 -1106 36920
rect 814 35000 815 36920
rect -1107 34999 815 35000
rect -1530 34652 -1426 34948
rect -3719 34600 -1797 34601
rect -3719 32680 -3718 34600
rect -1798 32680 -1797 34600
rect -3719 32679 -1797 32680
rect -4142 32332 -4038 32628
rect -6331 32280 -4409 32281
rect -6331 30360 -6330 32280
rect -4410 30360 -4409 32280
rect -6331 30359 -4409 30360
rect -5422 29961 -5318 30359
rect -4142 30308 -4122 32332
rect -4058 30308 -4038 32332
rect -2810 32281 -2706 32679
rect -1530 32628 -1510 34652
rect -1446 32628 -1426 34652
rect -198 34601 -94 34999
rect 1082 34948 1102 36972
rect 1166 34948 1186 36972
rect 2414 36921 2518 37120
rect 3694 36972 3798 37120
rect 1505 36920 3427 36921
rect 1505 35000 1506 36920
rect 3426 35000 3427 36920
rect 1505 34999 3427 35000
rect 1082 34652 1186 34948
rect -1107 34600 815 34601
rect -1107 32680 -1106 34600
rect 814 32680 815 34600
rect -1107 32679 815 32680
rect -1530 32332 -1426 32628
rect -3719 32280 -1797 32281
rect -3719 30360 -3718 32280
rect -1798 30360 -1797 32280
rect -3719 30359 -1797 30360
rect -4142 30012 -4038 30308
rect -6331 29960 -4409 29961
rect -6331 28040 -6330 29960
rect -4410 28040 -4409 29960
rect -6331 28039 -4409 28040
rect -5422 27641 -5318 28039
rect -4142 27988 -4122 30012
rect -4058 27988 -4038 30012
rect -2810 29961 -2706 30359
rect -1530 30308 -1510 32332
rect -1446 30308 -1426 32332
rect -198 32281 -94 32679
rect 1082 32628 1102 34652
rect 1166 32628 1186 34652
rect 2414 34601 2518 34999
rect 3694 34948 3714 36972
rect 3778 34948 3798 36972
rect 5026 36921 5130 37120
rect 6306 36972 6410 37120
rect 4117 36920 6039 36921
rect 4117 35000 4118 36920
rect 6038 35000 6039 36920
rect 4117 34999 6039 35000
rect 3694 34652 3798 34948
rect 1505 34600 3427 34601
rect 1505 32680 1506 34600
rect 3426 32680 3427 34600
rect 1505 32679 3427 32680
rect 1082 32332 1186 32628
rect -1107 32280 815 32281
rect -1107 30360 -1106 32280
rect 814 30360 815 32280
rect -1107 30359 815 30360
rect -1530 30012 -1426 30308
rect -3719 29960 -1797 29961
rect -3719 28040 -3718 29960
rect -1798 28040 -1797 29960
rect -3719 28039 -1797 28040
rect -4142 27692 -4038 27988
rect -6331 27640 -4409 27641
rect -6331 25720 -6330 27640
rect -4410 25720 -4409 27640
rect -6331 25719 -4409 25720
rect -5422 25321 -5318 25719
rect -4142 25668 -4122 27692
rect -4058 25668 -4038 27692
rect -2810 27641 -2706 28039
rect -1530 27988 -1510 30012
rect -1446 27988 -1426 30012
rect -198 29961 -94 30359
rect 1082 30308 1102 32332
rect 1166 30308 1186 32332
rect 2414 32281 2518 32679
rect 3694 32628 3714 34652
rect 3778 32628 3798 34652
rect 5026 34601 5130 34999
rect 6306 34948 6326 36972
rect 6390 34948 6410 36972
rect 6306 34652 6410 34948
rect 4117 34600 6039 34601
rect 4117 32680 4118 34600
rect 6038 32680 6039 34600
rect 4117 32679 6039 32680
rect 3694 32332 3798 32628
rect 1505 32280 3427 32281
rect 1505 30360 1506 32280
rect 3426 30360 3427 32280
rect 1505 30359 3427 30360
rect 1082 30012 1186 30308
rect -1107 29960 815 29961
rect -1107 28040 -1106 29960
rect 814 28040 815 29960
rect -1107 28039 815 28040
rect -1530 27692 -1426 27988
rect -3719 27640 -1797 27641
rect -3719 25720 -3718 27640
rect -1798 25720 -1797 27640
rect -3719 25719 -1797 25720
rect -4142 25372 -4038 25668
rect -6331 25320 -4409 25321
rect -6331 23400 -6330 25320
rect -4410 23400 -4409 25320
rect -6331 23399 -4409 23400
rect -5422 23001 -5318 23399
rect -4142 23348 -4122 25372
rect -4058 23348 -4038 25372
rect -2810 25321 -2706 25719
rect -1530 25668 -1510 27692
rect -1446 25668 -1426 27692
rect -198 27641 -94 28039
rect 1082 27988 1102 30012
rect 1166 27988 1186 30012
rect 2414 29961 2518 30359
rect 3694 30308 3714 32332
rect 3778 30308 3798 32332
rect 5026 32281 5130 32679
rect 6306 32628 6326 34652
rect 6390 32628 6410 34652
rect 6306 32332 6410 32628
rect 4117 32280 6039 32281
rect 4117 30360 4118 32280
rect 6038 30360 6039 32280
rect 4117 30359 6039 30360
rect 3694 30012 3798 30308
rect 1505 29960 3427 29961
rect 1505 28040 1506 29960
rect 3426 28040 3427 29960
rect 1505 28039 3427 28040
rect 1082 27692 1186 27988
rect -1107 27640 815 27641
rect -1107 25720 -1106 27640
rect 814 25720 815 27640
rect -1107 25719 815 25720
rect -1530 25372 -1426 25668
rect -3719 25320 -1797 25321
rect -3719 23400 -3718 25320
rect -1798 23400 -1797 25320
rect -3719 23399 -1797 23400
rect -4142 23052 -4038 23348
rect -6331 23000 -4409 23001
rect -6331 21080 -6330 23000
rect -4410 21080 -4409 23000
rect -6331 21079 -4409 21080
rect -5422 20681 -5318 21079
rect -4142 21028 -4122 23052
rect -4058 21028 -4038 23052
rect -2810 23001 -2706 23399
rect -1530 23348 -1510 25372
rect -1446 23348 -1426 25372
rect -198 25321 -94 25719
rect 1082 25668 1102 27692
rect 1166 25668 1186 27692
rect 2414 27641 2518 28039
rect 3694 27988 3714 30012
rect 3778 27988 3798 30012
rect 5026 29961 5130 30359
rect 6306 30308 6326 32332
rect 6390 30308 6410 32332
rect 6306 30012 6410 30308
rect 4117 29960 6039 29961
rect 4117 28040 4118 29960
rect 6038 28040 6039 29960
rect 4117 28039 6039 28040
rect 3694 27692 3798 27988
rect 1505 27640 3427 27641
rect 1505 25720 1506 27640
rect 3426 25720 3427 27640
rect 1505 25719 3427 25720
rect 1082 25372 1186 25668
rect -1107 25320 815 25321
rect -1107 23400 -1106 25320
rect 814 23400 815 25320
rect -1107 23399 815 23400
rect -1530 23052 -1426 23348
rect -3719 23000 -1797 23001
rect -3719 21080 -3718 23000
rect -1798 21080 -1797 23000
rect -3719 21079 -1797 21080
rect -4142 20732 -4038 21028
rect -6331 20680 -4409 20681
rect -6331 18760 -6330 20680
rect -4410 18760 -4409 20680
rect -6331 18759 -4409 18760
rect -5422 18361 -5318 18759
rect -4142 18708 -4122 20732
rect -4058 18708 -4038 20732
rect -2810 20681 -2706 21079
rect -1530 21028 -1510 23052
rect -1446 21028 -1426 23052
rect -198 23001 -94 23399
rect 1082 23348 1102 25372
rect 1166 23348 1186 25372
rect 2414 25321 2518 25719
rect 3694 25668 3714 27692
rect 3778 25668 3798 27692
rect 5026 27641 5130 28039
rect 6306 27988 6326 30012
rect 6390 27988 6410 30012
rect 6306 27692 6410 27988
rect 4117 27640 6039 27641
rect 4117 25720 4118 27640
rect 6038 25720 6039 27640
rect 4117 25719 6039 25720
rect 3694 25372 3798 25668
rect 1505 25320 3427 25321
rect 1505 23400 1506 25320
rect 3426 23400 3427 25320
rect 1505 23399 3427 23400
rect 1082 23052 1186 23348
rect -1107 23000 815 23001
rect -1107 21080 -1106 23000
rect 814 21080 815 23000
rect -1107 21079 815 21080
rect -1530 20732 -1426 21028
rect -3719 20680 -1797 20681
rect -3719 18760 -3718 20680
rect -1798 18760 -1797 20680
rect -3719 18759 -1797 18760
rect -4142 18412 -4038 18708
rect -6331 18360 -4409 18361
rect -6331 16440 -6330 18360
rect -4410 16440 -4409 18360
rect -6331 16439 -4409 16440
rect -5422 16041 -5318 16439
rect -4142 16388 -4122 18412
rect -4058 16388 -4038 18412
rect -2810 18361 -2706 18759
rect -1530 18708 -1510 20732
rect -1446 18708 -1426 20732
rect -198 20681 -94 21079
rect 1082 21028 1102 23052
rect 1166 21028 1186 23052
rect 2414 23001 2518 23399
rect 3694 23348 3714 25372
rect 3778 23348 3798 25372
rect 5026 25321 5130 25719
rect 6306 25668 6326 27692
rect 6390 25668 6410 27692
rect 6306 25372 6410 25668
rect 4117 25320 6039 25321
rect 4117 23400 4118 25320
rect 6038 23400 6039 25320
rect 4117 23399 6039 23400
rect 3694 23052 3798 23348
rect 1505 23000 3427 23001
rect 1505 21080 1506 23000
rect 3426 21080 3427 23000
rect 1505 21079 3427 21080
rect 1082 20732 1186 21028
rect -1107 20680 815 20681
rect -1107 18760 -1106 20680
rect 814 18760 815 20680
rect -1107 18759 815 18760
rect -1530 18412 -1426 18708
rect -3719 18360 -1797 18361
rect -3719 16440 -3718 18360
rect -1798 16440 -1797 18360
rect -3719 16439 -1797 16440
rect -4142 16092 -4038 16388
rect -6331 16040 -4409 16041
rect -6331 14120 -6330 16040
rect -4410 14120 -4409 16040
rect -6331 14119 -4409 14120
rect -5422 13721 -5318 14119
rect -4142 14068 -4122 16092
rect -4058 14068 -4038 16092
rect -2810 16041 -2706 16439
rect -1530 16388 -1510 18412
rect -1446 16388 -1426 18412
rect -198 18361 -94 18759
rect 1082 18708 1102 20732
rect 1166 18708 1186 20732
rect 2414 20681 2518 21079
rect 3694 21028 3714 23052
rect 3778 21028 3798 23052
rect 5026 23001 5130 23399
rect 6306 23348 6326 25372
rect 6390 23348 6410 25372
rect 6306 23052 6410 23348
rect 4117 23000 6039 23001
rect 4117 21080 4118 23000
rect 6038 21080 6039 23000
rect 4117 21079 6039 21080
rect 3694 20732 3798 21028
rect 1505 20680 3427 20681
rect 1505 18760 1506 20680
rect 3426 18760 3427 20680
rect 1505 18759 3427 18760
rect 1082 18412 1186 18708
rect -1107 18360 815 18361
rect -1107 16440 -1106 18360
rect 814 16440 815 18360
rect -1107 16439 815 16440
rect -1530 16092 -1426 16388
rect -3719 16040 -1797 16041
rect -3719 14120 -3718 16040
rect -1798 14120 -1797 16040
rect -3719 14119 -1797 14120
rect -4142 13772 -4038 14068
rect -6331 13720 -4409 13721
rect -6331 11800 -6330 13720
rect -4410 11800 -4409 13720
rect -6331 11799 -4409 11800
rect -5422 11401 -5318 11799
rect -4142 11748 -4122 13772
rect -4058 11748 -4038 13772
rect -2810 13721 -2706 14119
rect -1530 14068 -1510 16092
rect -1446 14068 -1426 16092
rect -198 16041 -94 16439
rect 1082 16388 1102 18412
rect 1166 16388 1186 18412
rect 2414 18361 2518 18759
rect 3694 18708 3714 20732
rect 3778 18708 3798 20732
rect 5026 20681 5130 21079
rect 6306 21028 6326 23052
rect 6390 21028 6410 23052
rect 6306 20732 6410 21028
rect 4117 20680 6039 20681
rect 4117 18760 4118 20680
rect 6038 18760 6039 20680
rect 4117 18759 6039 18760
rect 3694 18412 3798 18708
rect 1505 18360 3427 18361
rect 1505 16440 1506 18360
rect 3426 16440 3427 18360
rect 1505 16439 3427 16440
rect 1082 16092 1186 16388
rect -1107 16040 815 16041
rect -1107 14120 -1106 16040
rect 814 14120 815 16040
rect -1107 14119 815 14120
rect -1530 13772 -1426 14068
rect -3719 13720 -1797 13721
rect -3719 11800 -3718 13720
rect -1798 11800 -1797 13720
rect -3719 11799 -1797 11800
rect -4142 11452 -4038 11748
rect -6331 11400 -4409 11401
rect -6331 9480 -6330 11400
rect -4410 9480 -4409 11400
rect -6331 9479 -4409 9480
rect -5422 9081 -5318 9479
rect -4142 9428 -4122 11452
rect -4058 9428 -4038 11452
rect -2810 11401 -2706 11799
rect -1530 11748 -1510 13772
rect -1446 11748 -1426 13772
rect -198 13721 -94 14119
rect 1082 14068 1102 16092
rect 1166 14068 1186 16092
rect 2414 16041 2518 16439
rect 3694 16388 3714 18412
rect 3778 16388 3798 18412
rect 5026 18361 5130 18759
rect 6306 18708 6326 20732
rect 6390 18708 6410 20732
rect 6306 18412 6410 18708
rect 4117 18360 6039 18361
rect 4117 16440 4118 18360
rect 6038 16440 6039 18360
rect 4117 16439 6039 16440
rect 3694 16092 3798 16388
rect 1505 16040 3427 16041
rect 1505 14120 1506 16040
rect 3426 14120 3427 16040
rect 1505 14119 3427 14120
rect 1082 13772 1186 14068
rect -1107 13720 815 13721
rect -1107 11800 -1106 13720
rect 814 11800 815 13720
rect -1107 11799 815 11800
rect -1530 11452 -1426 11748
rect -3719 11400 -1797 11401
rect -3719 9480 -3718 11400
rect -1798 9480 -1797 11400
rect -3719 9479 -1797 9480
rect -4142 9132 -4038 9428
rect -6331 9080 -4409 9081
rect -6331 7160 -6330 9080
rect -4410 7160 -4409 9080
rect -6331 7159 -4409 7160
rect -5422 6761 -5318 7159
rect -4142 7108 -4122 9132
rect -4058 7108 -4038 9132
rect -2810 9081 -2706 9479
rect -1530 9428 -1510 11452
rect -1446 9428 -1426 11452
rect -198 11401 -94 11799
rect 1082 11748 1102 13772
rect 1166 11748 1186 13772
rect 2414 13721 2518 14119
rect 3694 14068 3714 16092
rect 3778 14068 3798 16092
rect 5026 16041 5130 16439
rect 6306 16388 6326 18412
rect 6390 16388 6410 18412
rect 6306 16092 6410 16388
rect 4117 16040 6039 16041
rect 4117 14120 4118 16040
rect 6038 14120 6039 16040
rect 4117 14119 6039 14120
rect 3694 13772 3798 14068
rect 1505 13720 3427 13721
rect 1505 11800 1506 13720
rect 3426 11800 3427 13720
rect 1505 11799 3427 11800
rect 1082 11452 1186 11748
rect -1107 11400 815 11401
rect -1107 9480 -1106 11400
rect 814 9480 815 11400
rect -1107 9479 815 9480
rect -1530 9132 -1426 9428
rect -3719 9080 -1797 9081
rect -3719 7160 -3718 9080
rect -1798 7160 -1797 9080
rect -3719 7159 -1797 7160
rect -4142 6812 -4038 7108
rect -6331 6760 -4409 6761
rect -6331 4840 -6330 6760
rect -4410 4840 -4409 6760
rect -6331 4839 -4409 4840
rect -5422 4441 -5318 4839
rect -4142 4788 -4122 6812
rect -4058 4788 -4038 6812
rect -2810 6761 -2706 7159
rect -1530 7108 -1510 9132
rect -1446 7108 -1426 9132
rect -198 9081 -94 9479
rect 1082 9428 1102 11452
rect 1166 9428 1186 11452
rect 2414 11401 2518 11799
rect 3694 11748 3714 13772
rect 3778 11748 3798 13772
rect 5026 13721 5130 14119
rect 6306 14068 6326 16092
rect 6390 14068 6410 16092
rect 6306 13772 6410 14068
rect 4117 13720 6039 13721
rect 4117 11800 4118 13720
rect 6038 11800 6039 13720
rect 4117 11799 6039 11800
rect 3694 11452 3798 11748
rect 1505 11400 3427 11401
rect 1505 9480 1506 11400
rect 3426 9480 3427 11400
rect 1505 9479 3427 9480
rect 1082 9132 1186 9428
rect -1107 9080 815 9081
rect -1107 7160 -1106 9080
rect 814 7160 815 9080
rect -1107 7159 815 7160
rect -1530 6812 -1426 7108
rect -3719 6760 -1797 6761
rect -3719 4840 -3718 6760
rect -1798 4840 -1797 6760
rect -3719 4839 -1797 4840
rect -4142 4492 -4038 4788
rect -6331 4440 -4409 4441
rect -6331 2520 -6330 4440
rect -4410 2520 -4409 4440
rect -6331 2519 -4409 2520
rect -5422 2121 -5318 2519
rect -4142 2468 -4122 4492
rect -4058 2468 -4038 4492
rect -2810 4441 -2706 4839
rect -1530 4788 -1510 6812
rect -1446 4788 -1426 6812
rect -198 6761 -94 7159
rect 1082 7108 1102 9132
rect 1166 7108 1186 9132
rect 2414 9081 2518 9479
rect 3694 9428 3714 11452
rect 3778 9428 3798 11452
rect 5026 11401 5130 11799
rect 6306 11748 6326 13772
rect 6390 11748 6410 13772
rect 6306 11452 6410 11748
rect 4117 11400 6039 11401
rect 4117 9480 4118 11400
rect 6038 9480 6039 11400
rect 4117 9479 6039 9480
rect 3694 9132 3798 9428
rect 1505 9080 3427 9081
rect 1505 7160 1506 9080
rect 3426 7160 3427 9080
rect 1505 7159 3427 7160
rect 1082 6812 1186 7108
rect -1107 6760 815 6761
rect -1107 4840 -1106 6760
rect 814 4840 815 6760
rect -1107 4839 815 4840
rect -1530 4492 -1426 4788
rect -3719 4440 -1797 4441
rect -3719 2520 -3718 4440
rect -1798 2520 -1797 4440
rect -3719 2519 -1797 2520
rect -4142 2172 -4038 2468
rect -6331 2120 -4409 2121
rect -6331 200 -6330 2120
rect -4410 200 -4409 2120
rect -6331 199 -4409 200
rect -5422 -199 -5318 199
rect -4142 148 -4122 2172
rect -4058 148 -4038 2172
rect -2810 2121 -2706 2519
rect -1530 2468 -1510 4492
rect -1446 2468 -1426 4492
rect -198 4441 -94 4839
rect 1082 4788 1102 6812
rect 1166 4788 1186 6812
rect 2414 6761 2518 7159
rect 3694 7108 3714 9132
rect 3778 7108 3798 9132
rect 5026 9081 5130 9479
rect 6306 9428 6326 11452
rect 6390 9428 6410 11452
rect 6306 9132 6410 9428
rect 4117 9080 6039 9081
rect 4117 7160 4118 9080
rect 6038 7160 6039 9080
rect 4117 7159 6039 7160
rect 3694 6812 3798 7108
rect 1505 6760 3427 6761
rect 1505 4840 1506 6760
rect 3426 4840 3427 6760
rect 1505 4839 3427 4840
rect 1082 4492 1186 4788
rect -1107 4440 815 4441
rect -1107 2520 -1106 4440
rect 814 2520 815 4440
rect -1107 2519 815 2520
rect -1530 2172 -1426 2468
rect -3719 2120 -1797 2121
rect -3719 200 -3718 2120
rect -1798 200 -1797 2120
rect -3719 199 -1797 200
rect -4142 -148 -4038 148
rect -6331 -200 -4409 -199
rect -6331 -2120 -6330 -200
rect -4410 -2120 -4409 -200
rect -6331 -2121 -4409 -2120
rect -5422 -2519 -5318 -2121
rect -4142 -2172 -4122 -148
rect -4058 -2172 -4038 -148
rect -2810 -199 -2706 199
rect -1530 148 -1510 2172
rect -1446 148 -1426 2172
rect -198 2121 -94 2519
rect 1082 2468 1102 4492
rect 1166 2468 1186 4492
rect 2414 4441 2518 4839
rect 3694 4788 3714 6812
rect 3778 4788 3798 6812
rect 5026 6761 5130 7159
rect 6306 7108 6326 9132
rect 6390 7108 6410 9132
rect 6306 6812 6410 7108
rect 4117 6760 6039 6761
rect 4117 4840 4118 6760
rect 6038 4840 6039 6760
rect 4117 4839 6039 4840
rect 3694 4492 3798 4788
rect 1505 4440 3427 4441
rect 1505 2520 1506 4440
rect 3426 2520 3427 4440
rect 1505 2519 3427 2520
rect 1082 2172 1186 2468
rect -1107 2120 815 2121
rect -1107 200 -1106 2120
rect 814 200 815 2120
rect -1107 199 815 200
rect -1530 -148 -1426 148
rect -3719 -200 -1797 -199
rect -3719 -2120 -3718 -200
rect -1798 -2120 -1797 -200
rect -3719 -2121 -1797 -2120
rect -4142 -2468 -4038 -2172
rect -6331 -2520 -4409 -2519
rect -6331 -4440 -6330 -2520
rect -4410 -4440 -4409 -2520
rect -6331 -4441 -4409 -4440
rect -5422 -4839 -5318 -4441
rect -4142 -4492 -4122 -2468
rect -4058 -4492 -4038 -2468
rect -2810 -2519 -2706 -2121
rect -1530 -2172 -1510 -148
rect -1446 -2172 -1426 -148
rect -198 -199 -94 199
rect 1082 148 1102 2172
rect 1166 148 1186 2172
rect 2414 2121 2518 2519
rect 3694 2468 3714 4492
rect 3778 2468 3798 4492
rect 5026 4441 5130 4839
rect 6306 4788 6326 6812
rect 6390 4788 6410 6812
rect 6306 4492 6410 4788
rect 4117 4440 6039 4441
rect 4117 2520 4118 4440
rect 6038 2520 6039 4440
rect 4117 2519 6039 2520
rect 3694 2172 3798 2468
rect 1505 2120 3427 2121
rect 1505 200 1506 2120
rect 3426 200 3427 2120
rect 1505 199 3427 200
rect 1082 -148 1186 148
rect -1107 -200 815 -199
rect -1107 -2120 -1106 -200
rect 814 -2120 815 -200
rect -1107 -2121 815 -2120
rect -1530 -2468 -1426 -2172
rect -3719 -2520 -1797 -2519
rect -3719 -4440 -3718 -2520
rect -1798 -4440 -1797 -2520
rect -3719 -4441 -1797 -4440
rect -4142 -4788 -4038 -4492
rect -6331 -4840 -4409 -4839
rect -6331 -6760 -6330 -4840
rect -4410 -6760 -4409 -4840
rect -6331 -6761 -4409 -6760
rect -5422 -7159 -5318 -6761
rect -4142 -6812 -4122 -4788
rect -4058 -6812 -4038 -4788
rect -2810 -4839 -2706 -4441
rect -1530 -4492 -1510 -2468
rect -1446 -4492 -1426 -2468
rect -198 -2519 -94 -2121
rect 1082 -2172 1102 -148
rect 1166 -2172 1186 -148
rect 2414 -199 2518 199
rect 3694 148 3714 2172
rect 3778 148 3798 2172
rect 5026 2121 5130 2519
rect 6306 2468 6326 4492
rect 6390 2468 6410 4492
rect 6306 2172 6410 2468
rect 4117 2120 6039 2121
rect 4117 200 4118 2120
rect 6038 200 6039 2120
rect 4117 199 6039 200
rect 3694 -148 3798 148
rect 1505 -200 3427 -199
rect 1505 -2120 1506 -200
rect 3426 -2120 3427 -200
rect 1505 -2121 3427 -2120
rect 1082 -2468 1186 -2172
rect -1107 -2520 815 -2519
rect -1107 -4440 -1106 -2520
rect 814 -4440 815 -2520
rect -1107 -4441 815 -4440
rect -1530 -4788 -1426 -4492
rect -3719 -4840 -1797 -4839
rect -3719 -6760 -3718 -4840
rect -1798 -6760 -1797 -4840
rect -3719 -6761 -1797 -6760
rect -4142 -7108 -4038 -6812
rect -6331 -7160 -4409 -7159
rect -6331 -9080 -6330 -7160
rect -4410 -9080 -4409 -7160
rect -6331 -9081 -4409 -9080
rect -5422 -9479 -5318 -9081
rect -4142 -9132 -4122 -7108
rect -4058 -9132 -4038 -7108
rect -2810 -7159 -2706 -6761
rect -1530 -6812 -1510 -4788
rect -1446 -6812 -1426 -4788
rect -198 -4839 -94 -4441
rect 1082 -4492 1102 -2468
rect 1166 -4492 1186 -2468
rect 2414 -2519 2518 -2121
rect 3694 -2172 3714 -148
rect 3778 -2172 3798 -148
rect 5026 -199 5130 199
rect 6306 148 6326 2172
rect 6390 148 6410 2172
rect 6306 -148 6410 148
rect 4117 -200 6039 -199
rect 4117 -2120 4118 -200
rect 6038 -2120 6039 -200
rect 4117 -2121 6039 -2120
rect 3694 -2468 3798 -2172
rect 1505 -2520 3427 -2519
rect 1505 -4440 1506 -2520
rect 3426 -4440 3427 -2520
rect 1505 -4441 3427 -4440
rect 1082 -4788 1186 -4492
rect -1107 -4840 815 -4839
rect -1107 -6760 -1106 -4840
rect 814 -6760 815 -4840
rect -1107 -6761 815 -6760
rect -1530 -7108 -1426 -6812
rect -3719 -7160 -1797 -7159
rect -3719 -9080 -3718 -7160
rect -1798 -9080 -1797 -7160
rect -3719 -9081 -1797 -9080
rect -4142 -9428 -4038 -9132
rect -6331 -9480 -4409 -9479
rect -6331 -11400 -6330 -9480
rect -4410 -11400 -4409 -9480
rect -6331 -11401 -4409 -11400
rect -5422 -11799 -5318 -11401
rect -4142 -11452 -4122 -9428
rect -4058 -11452 -4038 -9428
rect -2810 -9479 -2706 -9081
rect -1530 -9132 -1510 -7108
rect -1446 -9132 -1426 -7108
rect -198 -7159 -94 -6761
rect 1082 -6812 1102 -4788
rect 1166 -6812 1186 -4788
rect 2414 -4839 2518 -4441
rect 3694 -4492 3714 -2468
rect 3778 -4492 3798 -2468
rect 5026 -2519 5130 -2121
rect 6306 -2172 6326 -148
rect 6390 -2172 6410 -148
rect 6306 -2468 6410 -2172
rect 4117 -2520 6039 -2519
rect 4117 -4440 4118 -2520
rect 6038 -4440 6039 -2520
rect 4117 -4441 6039 -4440
rect 3694 -4788 3798 -4492
rect 1505 -4840 3427 -4839
rect 1505 -6760 1506 -4840
rect 3426 -6760 3427 -4840
rect 1505 -6761 3427 -6760
rect 1082 -7108 1186 -6812
rect -1107 -7160 815 -7159
rect -1107 -9080 -1106 -7160
rect 814 -9080 815 -7160
rect -1107 -9081 815 -9080
rect -1530 -9428 -1426 -9132
rect -3719 -9480 -1797 -9479
rect -3719 -11400 -3718 -9480
rect -1798 -11400 -1797 -9480
rect -3719 -11401 -1797 -11400
rect -4142 -11748 -4038 -11452
rect -6331 -11800 -4409 -11799
rect -6331 -13720 -6330 -11800
rect -4410 -13720 -4409 -11800
rect -6331 -13721 -4409 -13720
rect -5422 -14119 -5318 -13721
rect -4142 -13772 -4122 -11748
rect -4058 -13772 -4038 -11748
rect -2810 -11799 -2706 -11401
rect -1530 -11452 -1510 -9428
rect -1446 -11452 -1426 -9428
rect -198 -9479 -94 -9081
rect 1082 -9132 1102 -7108
rect 1166 -9132 1186 -7108
rect 2414 -7159 2518 -6761
rect 3694 -6812 3714 -4788
rect 3778 -6812 3798 -4788
rect 5026 -4839 5130 -4441
rect 6306 -4492 6326 -2468
rect 6390 -4492 6410 -2468
rect 6306 -4788 6410 -4492
rect 4117 -4840 6039 -4839
rect 4117 -6760 4118 -4840
rect 6038 -6760 6039 -4840
rect 4117 -6761 6039 -6760
rect 3694 -7108 3798 -6812
rect 1505 -7160 3427 -7159
rect 1505 -9080 1506 -7160
rect 3426 -9080 3427 -7160
rect 1505 -9081 3427 -9080
rect 1082 -9428 1186 -9132
rect -1107 -9480 815 -9479
rect -1107 -11400 -1106 -9480
rect 814 -11400 815 -9480
rect -1107 -11401 815 -11400
rect -1530 -11748 -1426 -11452
rect -3719 -11800 -1797 -11799
rect -3719 -13720 -3718 -11800
rect -1798 -13720 -1797 -11800
rect -3719 -13721 -1797 -13720
rect -4142 -14068 -4038 -13772
rect -6331 -14120 -4409 -14119
rect -6331 -16040 -6330 -14120
rect -4410 -16040 -4409 -14120
rect -6331 -16041 -4409 -16040
rect -5422 -16439 -5318 -16041
rect -4142 -16092 -4122 -14068
rect -4058 -16092 -4038 -14068
rect -2810 -14119 -2706 -13721
rect -1530 -13772 -1510 -11748
rect -1446 -13772 -1426 -11748
rect -198 -11799 -94 -11401
rect 1082 -11452 1102 -9428
rect 1166 -11452 1186 -9428
rect 2414 -9479 2518 -9081
rect 3694 -9132 3714 -7108
rect 3778 -9132 3798 -7108
rect 5026 -7159 5130 -6761
rect 6306 -6812 6326 -4788
rect 6390 -6812 6410 -4788
rect 6306 -7108 6410 -6812
rect 4117 -7160 6039 -7159
rect 4117 -9080 4118 -7160
rect 6038 -9080 6039 -7160
rect 4117 -9081 6039 -9080
rect 3694 -9428 3798 -9132
rect 1505 -9480 3427 -9479
rect 1505 -11400 1506 -9480
rect 3426 -11400 3427 -9480
rect 1505 -11401 3427 -11400
rect 1082 -11748 1186 -11452
rect -1107 -11800 815 -11799
rect -1107 -13720 -1106 -11800
rect 814 -13720 815 -11800
rect -1107 -13721 815 -13720
rect -1530 -14068 -1426 -13772
rect -3719 -14120 -1797 -14119
rect -3719 -16040 -3718 -14120
rect -1798 -16040 -1797 -14120
rect -3719 -16041 -1797 -16040
rect -4142 -16388 -4038 -16092
rect -6331 -16440 -4409 -16439
rect -6331 -18360 -6330 -16440
rect -4410 -18360 -4409 -16440
rect -6331 -18361 -4409 -18360
rect -5422 -18759 -5318 -18361
rect -4142 -18412 -4122 -16388
rect -4058 -18412 -4038 -16388
rect -2810 -16439 -2706 -16041
rect -1530 -16092 -1510 -14068
rect -1446 -16092 -1426 -14068
rect -198 -14119 -94 -13721
rect 1082 -13772 1102 -11748
rect 1166 -13772 1186 -11748
rect 2414 -11799 2518 -11401
rect 3694 -11452 3714 -9428
rect 3778 -11452 3798 -9428
rect 5026 -9479 5130 -9081
rect 6306 -9132 6326 -7108
rect 6390 -9132 6410 -7108
rect 6306 -9428 6410 -9132
rect 4117 -9480 6039 -9479
rect 4117 -11400 4118 -9480
rect 6038 -11400 6039 -9480
rect 4117 -11401 6039 -11400
rect 3694 -11748 3798 -11452
rect 1505 -11800 3427 -11799
rect 1505 -13720 1506 -11800
rect 3426 -13720 3427 -11800
rect 1505 -13721 3427 -13720
rect 1082 -14068 1186 -13772
rect -1107 -14120 815 -14119
rect -1107 -16040 -1106 -14120
rect 814 -16040 815 -14120
rect -1107 -16041 815 -16040
rect -1530 -16388 -1426 -16092
rect -3719 -16440 -1797 -16439
rect -3719 -18360 -3718 -16440
rect -1798 -18360 -1797 -16440
rect -3719 -18361 -1797 -18360
rect -4142 -18708 -4038 -18412
rect -6331 -18760 -4409 -18759
rect -6331 -20680 -6330 -18760
rect -4410 -20680 -4409 -18760
rect -6331 -20681 -4409 -20680
rect -5422 -21079 -5318 -20681
rect -4142 -20732 -4122 -18708
rect -4058 -20732 -4038 -18708
rect -2810 -18759 -2706 -18361
rect -1530 -18412 -1510 -16388
rect -1446 -18412 -1426 -16388
rect -198 -16439 -94 -16041
rect 1082 -16092 1102 -14068
rect 1166 -16092 1186 -14068
rect 2414 -14119 2518 -13721
rect 3694 -13772 3714 -11748
rect 3778 -13772 3798 -11748
rect 5026 -11799 5130 -11401
rect 6306 -11452 6326 -9428
rect 6390 -11452 6410 -9428
rect 6306 -11748 6410 -11452
rect 4117 -11800 6039 -11799
rect 4117 -13720 4118 -11800
rect 6038 -13720 6039 -11800
rect 4117 -13721 6039 -13720
rect 3694 -14068 3798 -13772
rect 1505 -14120 3427 -14119
rect 1505 -16040 1506 -14120
rect 3426 -16040 3427 -14120
rect 1505 -16041 3427 -16040
rect 1082 -16388 1186 -16092
rect -1107 -16440 815 -16439
rect -1107 -18360 -1106 -16440
rect 814 -18360 815 -16440
rect -1107 -18361 815 -18360
rect -1530 -18708 -1426 -18412
rect -3719 -18760 -1797 -18759
rect -3719 -20680 -3718 -18760
rect -1798 -20680 -1797 -18760
rect -3719 -20681 -1797 -20680
rect -4142 -21028 -4038 -20732
rect -6331 -21080 -4409 -21079
rect -6331 -23000 -6330 -21080
rect -4410 -23000 -4409 -21080
rect -6331 -23001 -4409 -23000
rect -5422 -23399 -5318 -23001
rect -4142 -23052 -4122 -21028
rect -4058 -23052 -4038 -21028
rect -2810 -21079 -2706 -20681
rect -1530 -20732 -1510 -18708
rect -1446 -20732 -1426 -18708
rect -198 -18759 -94 -18361
rect 1082 -18412 1102 -16388
rect 1166 -18412 1186 -16388
rect 2414 -16439 2518 -16041
rect 3694 -16092 3714 -14068
rect 3778 -16092 3798 -14068
rect 5026 -14119 5130 -13721
rect 6306 -13772 6326 -11748
rect 6390 -13772 6410 -11748
rect 6306 -14068 6410 -13772
rect 4117 -14120 6039 -14119
rect 4117 -16040 4118 -14120
rect 6038 -16040 6039 -14120
rect 4117 -16041 6039 -16040
rect 3694 -16388 3798 -16092
rect 1505 -16440 3427 -16439
rect 1505 -18360 1506 -16440
rect 3426 -18360 3427 -16440
rect 1505 -18361 3427 -18360
rect 1082 -18708 1186 -18412
rect -1107 -18760 815 -18759
rect -1107 -20680 -1106 -18760
rect 814 -20680 815 -18760
rect -1107 -20681 815 -20680
rect -1530 -21028 -1426 -20732
rect -3719 -21080 -1797 -21079
rect -3719 -23000 -3718 -21080
rect -1798 -23000 -1797 -21080
rect -3719 -23001 -1797 -23000
rect -4142 -23348 -4038 -23052
rect -6331 -23400 -4409 -23399
rect -6331 -25320 -6330 -23400
rect -4410 -25320 -4409 -23400
rect -6331 -25321 -4409 -25320
rect -5422 -25719 -5318 -25321
rect -4142 -25372 -4122 -23348
rect -4058 -25372 -4038 -23348
rect -2810 -23399 -2706 -23001
rect -1530 -23052 -1510 -21028
rect -1446 -23052 -1426 -21028
rect -198 -21079 -94 -20681
rect 1082 -20732 1102 -18708
rect 1166 -20732 1186 -18708
rect 2414 -18759 2518 -18361
rect 3694 -18412 3714 -16388
rect 3778 -18412 3798 -16388
rect 5026 -16439 5130 -16041
rect 6306 -16092 6326 -14068
rect 6390 -16092 6410 -14068
rect 6306 -16388 6410 -16092
rect 4117 -16440 6039 -16439
rect 4117 -18360 4118 -16440
rect 6038 -18360 6039 -16440
rect 4117 -18361 6039 -18360
rect 3694 -18708 3798 -18412
rect 1505 -18760 3427 -18759
rect 1505 -20680 1506 -18760
rect 3426 -20680 3427 -18760
rect 1505 -20681 3427 -20680
rect 1082 -21028 1186 -20732
rect -1107 -21080 815 -21079
rect -1107 -23000 -1106 -21080
rect 814 -23000 815 -21080
rect -1107 -23001 815 -23000
rect -1530 -23348 -1426 -23052
rect -3719 -23400 -1797 -23399
rect -3719 -25320 -3718 -23400
rect -1798 -25320 -1797 -23400
rect -3719 -25321 -1797 -25320
rect -4142 -25668 -4038 -25372
rect -6331 -25720 -4409 -25719
rect -6331 -27640 -6330 -25720
rect -4410 -27640 -4409 -25720
rect -6331 -27641 -4409 -27640
rect -5422 -28039 -5318 -27641
rect -4142 -27692 -4122 -25668
rect -4058 -27692 -4038 -25668
rect -2810 -25719 -2706 -25321
rect -1530 -25372 -1510 -23348
rect -1446 -25372 -1426 -23348
rect -198 -23399 -94 -23001
rect 1082 -23052 1102 -21028
rect 1166 -23052 1186 -21028
rect 2414 -21079 2518 -20681
rect 3694 -20732 3714 -18708
rect 3778 -20732 3798 -18708
rect 5026 -18759 5130 -18361
rect 6306 -18412 6326 -16388
rect 6390 -18412 6410 -16388
rect 6306 -18708 6410 -18412
rect 4117 -18760 6039 -18759
rect 4117 -20680 4118 -18760
rect 6038 -20680 6039 -18760
rect 4117 -20681 6039 -20680
rect 3694 -21028 3798 -20732
rect 1505 -21080 3427 -21079
rect 1505 -23000 1506 -21080
rect 3426 -23000 3427 -21080
rect 1505 -23001 3427 -23000
rect 1082 -23348 1186 -23052
rect -1107 -23400 815 -23399
rect -1107 -25320 -1106 -23400
rect 814 -25320 815 -23400
rect -1107 -25321 815 -25320
rect -1530 -25668 -1426 -25372
rect -3719 -25720 -1797 -25719
rect -3719 -27640 -3718 -25720
rect -1798 -27640 -1797 -25720
rect -3719 -27641 -1797 -27640
rect -4142 -27988 -4038 -27692
rect -6331 -28040 -4409 -28039
rect -6331 -29960 -6330 -28040
rect -4410 -29960 -4409 -28040
rect -6331 -29961 -4409 -29960
rect -5422 -30359 -5318 -29961
rect -4142 -30012 -4122 -27988
rect -4058 -30012 -4038 -27988
rect -2810 -28039 -2706 -27641
rect -1530 -27692 -1510 -25668
rect -1446 -27692 -1426 -25668
rect -198 -25719 -94 -25321
rect 1082 -25372 1102 -23348
rect 1166 -25372 1186 -23348
rect 2414 -23399 2518 -23001
rect 3694 -23052 3714 -21028
rect 3778 -23052 3798 -21028
rect 5026 -21079 5130 -20681
rect 6306 -20732 6326 -18708
rect 6390 -20732 6410 -18708
rect 6306 -21028 6410 -20732
rect 4117 -21080 6039 -21079
rect 4117 -23000 4118 -21080
rect 6038 -23000 6039 -21080
rect 4117 -23001 6039 -23000
rect 3694 -23348 3798 -23052
rect 1505 -23400 3427 -23399
rect 1505 -25320 1506 -23400
rect 3426 -25320 3427 -23400
rect 1505 -25321 3427 -25320
rect 1082 -25668 1186 -25372
rect -1107 -25720 815 -25719
rect -1107 -27640 -1106 -25720
rect 814 -27640 815 -25720
rect -1107 -27641 815 -27640
rect -1530 -27988 -1426 -27692
rect -3719 -28040 -1797 -28039
rect -3719 -29960 -3718 -28040
rect -1798 -29960 -1797 -28040
rect -3719 -29961 -1797 -29960
rect -4142 -30308 -4038 -30012
rect -6331 -30360 -4409 -30359
rect -6331 -32280 -6330 -30360
rect -4410 -32280 -4409 -30360
rect -6331 -32281 -4409 -32280
rect -5422 -32679 -5318 -32281
rect -4142 -32332 -4122 -30308
rect -4058 -32332 -4038 -30308
rect -2810 -30359 -2706 -29961
rect -1530 -30012 -1510 -27988
rect -1446 -30012 -1426 -27988
rect -198 -28039 -94 -27641
rect 1082 -27692 1102 -25668
rect 1166 -27692 1186 -25668
rect 2414 -25719 2518 -25321
rect 3694 -25372 3714 -23348
rect 3778 -25372 3798 -23348
rect 5026 -23399 5130 -23001
rect 6306 -23052 6326 -21028
rect 6390 -23052 6410 -21028
rect 6306 -23348 6410 -23052
rect 4117 -23400 6039 -23399
rect 4117 -25320 4118 -23400
rect 6038 -25320 6039 -23400
rect 4117 -25321 6039 -25320
rect 3694 -25668 3798 -25372
rect 1505 -25720 3427 -25719
rect 1505 -27640 1506 -25720
rect 3426 -27640 3427 -25720
rect 1505 -27641 3427 -27640
rect 1082 -27988 1186 -27692
rect -1107 -28040 815 -28039
rect -1107 -29960 -1106 -28040
rect 814 -29960 815 -28040
rect -1107 -29961 815 -29960
rect -1530 -30308 -1426 -30012
rect -3719 -30360 -1797 -30359
rect -3719 -32280 -3718 -30360
rect -1798 -32280 -1797 -30360
rect -3719 -32281 -1797 -32280
rect -4142 -32628 -4038 -32332
rect -6331 -32680 -4409 -32679
rect -6331 -34600 -6330 -32680
rect -4410 -34600 -4409 -32680
rect -6331 -34601 -4409 -34600
rect -5422 -34999 -5318 -34601
rect -4142 -34652 -4122 -32628
rect -4058 -34652 -4038 -32628
rect -2810 -32679 -2706 -32281
rect -1530 -32332 -1510 -30308
rect -1446 -32332 -1426 -30308
rect -198 -30359 -94 -29961
rect 1082 -30012 1102 -27988
rect 1166 -30012 1186 -27988
rect 2414 -28039 2518 -27641
rect 3694 -27692 3714 -25668
rect 3778 -27692 3798 -25668
rect 5026 -25719 5130 -25321
rect 6306 -25372 6326 -23348
rect 6390 -25372 6410 -23348
rect 6306 -25668 6410 -25372
rect 4117 -25720 6039 -25719
rect 4117 -27640 4118 -25720
rect 6038 -27640 6039 -25720
rect 4117 -27641 6039 -27640
rect 3694 -27988 3798 -27692
rect 1505 -28040 3427 -28039
rect 1505 -29960 1506 -28040
rect 3426 -29960 3427 -28040
rect 1505 -29961 3427 -29960
rect 1082 -30308 1186 -30012
rect -1107 -30360 815 -30359
rect -1107 -32280 -1106 -30360
rect 814 -32280 815 -30360
rect -1107 -32281 815 -32280
rect -1530 -32628 -1426 -32332
rect -3719 -32680 -1797 -32679
rect -3719 -34600 -3718 -32680
rect -1798 -34600 -1797 -32680
rect -3719 -34601 -1797 -34600
rect -4142 -34948 -4038 -34652
rect -6331 -35000 -4409 -34999
rect -6331 -36920 -6330 -35000
rect -4410 -36920 -4409 -35000
rect -6331 -36921 -4409 -36920
rect -5422 -37120 -5318 -36921
rect -4142 -36972 -4122 -34948
rect -4058 -36972 -4038 -34948
rect -2810 -34999 -2706 -34601
rect -1530 -34652 -1510 -32628
rect -1446 -34652 -1426 -32628
rect -198 -32679 -94 -32281
rect 1082 -32332 1102 -30308
rect 1166 -32332 1186 -30308
rect 2414 -30359 2518 -29961
rect 3694 -30012 3714 -27988
rect 3778 -30012 3798 -27988
rect 5026 -28039 5130 -27641
rect 6306 -27692 6326 -25668
rect 6390 -27692 6410 -25668
rect 6306 -27988 6410 -27692
rect 4117 -28040 6039 -28039
rect 4117 -29960 4118 -28040
rect 6038 -29960 6039 -28040
rect 4117 -29961 6039 -29960
rect 3694 -30308 3798 -30012
rect 1505 -30360 3427 -30359
rect 1505 -32280 1506 -30360
rect 3426 -32280 3427 -30360
rect 1505 -32281 3427 -32280
rect 1082 -32628 1186 -32332
rect -1107 -32680 815 -32679
rect -1107 -34600 -1106 -32680
rect 814 -34600 815 -32680
rect -1107 -34601 815 -34600
rect -1530 -34948 -1426 -34652
rect -3719 -35000 -1797 -34999
rect -3719 -36920 -3718 -35000
rect -1798 -36920 -1797 -35000
rect -3719 -36921 -1797 -36920
rect -4142 -37120 -4038 -36972
rect -2810 -37120 -2706 -36921
rect -1530 -36972 -1510 -34948
rect -1446 -36972 -1426 -34948
rect -198 -34999 -94 -34601
rect 1082 -34652 1102 -32628
rect 1166 -34652 1186 -32628
rect 2414 -32679 2518 -32281
rect 3694 -32332 3714 -30308
rect 3778 -32332 3798 -30308
rect 5026 -30359 5130 -29961
rect 6306 -30012 6326 -27988
rect 6390 -30012 6410 -27988
rect 6306 -30308 6410 -30012
rect 4117 -30360 6039 -30359
rect 4117 -32280 4118 -30360
rect 6038 -32280 6039 -30360
rect 4117 -32281 6039 -32280
rect 3694 -32628 3798 -32332
rect 1505 -32680 3427 -32679
rect 1505 -34600 1506 -32680
rect 3426 -34600 3427 -32680
rect 1505 -34601 3427 -34600
rect 1082 -34948 1186 -34652
rect -1107 -35000 815 -34999
rect -1107 -36920 -1106 -35000
rect 814 -36920 815 -35000
rect -1107 -36921 815 -36920
rect -1530 -37120 -1426 -36972
rect -198 -37120 -94 -36921
rect 1082 -36972 1102 -34948
rect 1166 -36972 1186 -34948
rect 2414 -34999 2518 -34601
rect 3694 -34652 3714 -32628
rect 3778 -34652 3798 -32628
rect 5026 -32679 5130 -32281
rect 6306 -32332 6326 -30308
rect 6390 -32332 6410 -30308
rect 6306 -32628 6410 -32332
rect 4117 -32680 6039 -32679
rect 4117 -34600 4118 -32680
rect 6038 -34600 6039 -32680
rect 4117 -34601 6039 -34600
rect 3694 -34948 3798 -34652
rect 1505 -35000 3427 -34999
rect 1505 -36920 1506 -35000
rect 3426 -36920 3427 -35000
rect 1505 -36921 3427 -36920
rect 1082 -37120 1186 -36972
rect 2414 -37120 2518 -36921
rect 3694 -36972 3714 -34948
rect 3778 -36972 3798 -34948
rect 5026 -34999 5130 -34601
rect 6306 -34652 6326 -32628
rect 6390 -34652 6410 -32628
rect 6306 -34948 6410 -34652
rect 4117 -35000 6039 -34999
rect 4117 -36920 4118 -35000
rect 6038 -36920 6039 -35000
rect 4117 -36921 6039 -36920
rect 3694 -37120 3798 -36972
rect 5026 -37120 5130 -36921
rect 6306 -36972 6326 -34948
rect 6390 -36972 6410 -34948
rect 6306 -37120 6410 -36972
<< properties >>
string FIXED_BBOX 4038 34920 6118 37000
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 5 ny 32 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
