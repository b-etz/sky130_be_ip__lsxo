magic
tech sky130A
magscale 1 2
timestamp 1712954147
<< pwell >>
rect -1612 -6832 1612 6832
<< psubdiff >>
rect -1576 6762 -1480 6796
rect 1480 6762 1576 6796
rect -1576 6700 -1542 6762
rect 1542 6700 1576 6762
rect -1576 -6762 -1542 -6700
rect 1542 -6762 1576 -6700
rect -1576 -6796 -1480 -6762
rect 1480 -6796 1576 -6762
<< psubdiffcont >>
rect -1480 6762 1480 6796
rect -1576 -6700 -1542 6700
rect 1542 -6700 1576 6700
rect -1480 -6796 1480 -6762
<< xpolycontact >>
rect -1446 6234 -1376 6666
rect -1446 -6666 -1376 -6234
rect -1280 6234 -1210 6666
rect -1280 -6666 -1210 -6234
rect -1114 6234 -1044 6666
rect -1114 -6666 -1044 -6234
rect -948 6234 -878 6666
rect -948 -6666 -878 -6234
rect -782 6234 -712 6666
rect -782 -6666 -712 -6234
rect -616 6234 -546 6666
rect -616 -6666 -546 -6234
rect -450 6234 -380 6666
rect -450 -6666 -380 -6234
rect -284 6234 -214 6666
rect -284 -6666 -214 -6234
rect -118 6234 -48 6666
rect -118 -6666 -48 -6234
rect 48 6234 118 6666
rect 48 -6666 118 -6234
rect 214 6234 284 6666
rect 214 -6666 284 -6234
rect 380 6234 450 6666
rect 380 -6666 450 -6234
rect 546 6234 616 6666
rect 546 -6666 616 -6234
rect 712 6234 782 6666
rect 712 -6666 782 -6234
rect 878 6234 948 6666
rect 878 -6666 948 -6234
rect 1044 6234 1114 6666
rect 1044 -6666 1114 -6234
rect 1210 6234 1280 6666
rect 1210 -6666 1280 -6234
rect 1376 6234 1446 6666
rect 1376 -6666 1446 -6234
<< xpolyres >>
rect -1446 -6234 -1376 6234
rect -1280 -6234 -1210 6234
rect -1114 -6234 -1044 6234
rect -948 -6234 -878 6234
rect -782 -6234 -712 6234
rect -616 -6234 -546 6234
rect -450 -6234 -380 6234
rect -284 -6234 -214 6234
rect -118 -6234 -48 6234
rect 48 -6234 118 6234
rect 214 -6234 284 6234
rect 380 -6234 450 6234
rect 546 -6234 616 6234
rect 712 -6234 782 6234
rect 878 -6234 948 6234
rect 1044 -6234 1114 6234
rect 1210 -6234 1280 6234
rect 1376 -6234 1446 6234
<< locali >>
rect -1576 6762 -1480 6796
rect 1480 6762 1576 6796
rect -1576 6700 -1542 6762
rect 1542 6700 1576 6762
rect -1576 -6762 -1542 -6700
rect 1542 -6762 1576 -6700
rect -1576 -6796 -1480 -6762
rect 1480 -6796 1576 -6762
<< viali >>
rect -1430 6251 -1392 6648
rect -1264 6251 -1226 6648
rect -1098 6251 -1060 6648
rect -932 6251 -894 6648
rect -766 6251 -728 6648
rect -600 6251 -562 6648
rect -434 6251 -396 6648
rect -268 6251 -230 6648
rect -102 6251 -64 6648
rect 64 6251 102 6648
rect 230 6251 268 6648
rect 396 6251 434 6648
rect 562 6251 600 6648
rect 728 6251 766 6648
rect 894 6251 932 6648
rect 1060 6251 1098 6648
rect 1226 6251 1264 6648
rect 1392 6251 1430 6648
rect -1430 -6648 -1392 -6251
rect -1264 -6648 -1226 -6251
rect -1098 -6648 -1060 -6251
rect -932 -6648 -894 -6251
rect -766 -6648 -728 -6251
rect -600 -6648 -562 -6251
rect -434 -6648 -396 -6251
rect -268 -6648 -230 -6251
rect -102 -6648 -64 -6251
rect 64 -6648 102 -6251
rect 230 -6648 268 -6251
rect 396 -6648 434 -6251
rect 562 -6648 600 -6251
rect 728 -6648 766 -6251
rect 894 -6648 932 -6251
rect 1060 -6648 1098 -6251
rect 1226 -6648 1264 -6251
rect 1392 -6648 1430 -6251
<< metal1 >>
rect -1436 6648 -1386 6660
rect -1436 6251 -1430 6648
rect -1392 6251 -1386 6648
rect -1436 6239 -1386 6251
rect -1270 6648 -1220 6660
rect -1270 6251 -1264 6648
rect -1226 6251 -1220 6648
rect -1270 6239 -1220 6251
rect -1104 6648 -1054 6660
rect -1104 6251 -1098 6648
rect -1060 6251 -1054 6648
rect -1104 6239 -1054 6251
rect -938 6648 -888 6660
rect -938 6251 -932 6648
rect -894 6251 -888 6648
rect -938 6239 -888 6251
rect -772 6648 -722 6660
rect -772 6251 -766 6648
rect -728 6251 -722 6648
rect -772 6239 -722 6251
rect -606 6648 -556 6660
rect -606 6251 -600 6648
rect -562 6251 -556 6648
rect -606 6239 -556 6251
rect -440 6648 -390 6660
rect -440 6251 -434 6648
rect -396 6251 -390 6648
rect -440 6239 -390 6251
rect -274 6648 -224 6660
rect -274 6251 -268 6648
rect -230 6251 -224 6648
rect -274 6239 -224 6251
rect -108 6648 -58 6660
rect -108 6251 -102 6648
rect -64 6251 -58 6648
rect -108 6239 -58 6251
rect 58 6648 108 6660
rect 58 6251 64 6648
rect 102 6251 108 6648
rect 58 6239 108 6251
rect 224 6648 274 6660
rect 224 6251 230 6648
rect 268 6251 274 6648
rect 224 6239 274 6251
rect 390 6648 440 6660
rect 390 6251 396 6648
rect 434 6251 440 6648
rect 390 6239 440 6251
rect 556 6648 606 6660
rect 556 6251 562 6648
rect 600 6251 606 6648
rect 556 6239 606 6251
rect 722 6648 772 6660
rect 722 6251 728 6648
rect 766 6251 772 6648
rect 722 6239 772 6251
rect 888 6648 938 6660
rect 888 6251 894 6648
rect 932 6251 938 6648
rect 888 6239 938 6251
rect 1054 6648 1104 6660
rect 1054 6251 1060 6648
rect 1098 6251 1104 6648
rect 1054 6239 1104 6251
rect 1220 6648 1270 6660
rect 1220 6251 1226 6648
rect 1264 6251 1270 6648
rect 1220 6239 1270 6251
rect 1386 6648 1436 6660
rect 1386 6251 1392 6648
rect 1430 6251 1436 6648
rect 1386 6239 1436 6251
rect -1436 -6251 -1386 -6239
rect -1436 -6648 -1430 -6251
rect -1392 -6648 -1386 -6251
rect -1436 -6660 -1386 -6648
rect -1270 -6251 -1220 -6239
rect -1270 -6648 -1264 -6251
rect -1226 -6648 -1220 -6251
rect -1270 -6660 -1220 -6648
rect -1104 -6251 -1054 -6239
rect -1104 -6648 -1098 -6251
rect -1060 -6648 -1054 -6251
rect -1104 -6660 -1054 -6648
rect -938 -6251 -888 -6239
rect -938 -6648 -932 -6251
rect -894 -6648 -888 -6251
rect -938 -6660 -888 -6648
rect -772 -6251 -722 -6239
rect -772 -6648 -766 -6251
rect -728 -6648 -722 -6251
rect -772 -6660 -722 -6648
rect -606 -6251 -556 -6239
rect -606 -6648 -600 -6251
rect -562 -6648 -556 -6251
rect -606 -6660 -556 -6648
rect -440 -6251 -390 -6239
rect -440 -6648 -434 -6251
rect -396 -6648 -390 -6251
rect -440 -6660 -390 -6648
rect -274 -6251 -224 -6239
rect -274 -6648 -268 -6251
rect -230 -6648 -224 -6251
rect -274 -6660 -224 -6648
rect -108 -6251 -58 -6239
rect -108 -6648 -102 -6251
rect -64 -6648 -58 -6251
rect -108 -6660 -58 -6648
rect 58 -6251 108 -6239
rect 58 -6648 64 -6251
rect 102 -6648 108 -6251
rect 58 -6660 108 -6648
rect 224 -6251 274 -6239
rect 224 -6648 230 -6251
rect 268 -6648 274 -6251
rect 224 -6660 274 -6648
rect 390 -6251 440 -6239
rect 390 -6648 396 -6251
rect 434 -6648 440 -6251
rect 390 -6660 440 -6648
rect 556 -6251 606 -6239
rect 556 -6648 562 -6251
rect 600 -6648 606 -6251
rect 556 -6660 606 -6648
rect 722 -6251 772 -6239
rect 722 -6648 728 -6251
rect 766 -6648 772 -6251
rect 722 -6660 772 -6648
rect 888 -6251 938 -6239
rect 888 -6648 894 -6251
rect 932 -6648 938 -6251
rect 888 -6660 938 -6648
rect 1054 -6251 1104 -6239
rect 1054 -6648 1060 -6251
rect 1098 -6648 1104 -6251
rect 1054 -6660 1104 -6648
rect 1220 -6251 1270 -6239
rect 1220 -6648 1226 -6251
rect 1264 -6648 1270 -6251
rect 1220 -6660 1270 -6648
rect 1386 -6251 1436 -6239
rect 1386 -6648 1392 -6251
rect 1430 -6648 1436 -6251
rect 1386 -6660 1436 -6648
<< properties >>
string FIXED_BBOX -1559 -6779 1559 6779
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 62.5 m 1 nx 18 wmin 0.350 lmin 0.50 rho 2000 val 358.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
