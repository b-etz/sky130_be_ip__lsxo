magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< pwell >>
rect -278 -5239 278 5239
<< mvnmos >>
rect -50 4181 50 4981
rect -50 3163 50 3963
rect -50 2145 50 2945
rect -50 1127 50 1927
rect -50 109 50 909
rect -50 -909 50 -109
rect -50 -1927 50 -1127
rect -50 -2945 50 -2145
rect -50 -3963 50 -3163
rect -50 -4981 50 -4181
<< mvndiff >>
rect -108 4969 -50 4981
rect -108 4193 -96 4969
rect -62 4193 -50 4969
rect -108 4181 -50 4193
rect 50 4969 108 4981
rect 50 4193 62 4969
rect 96 4193 108 4969
rect 50 4181 108 4193
rect -108 3951 -50 3963
rect -108 3175 -96 3951
rect -62 3175 -50 3951
rect -108 3163 -50 3175
rect 50 3951 108 3963
rect 50 3175 62 3951
rect 96 3175 108 3951
rect 50 3163 108 3175
rect -108 2933 -50 2945
rect -108 2157 -96 2933
rect -62 2157 -50 2933
rect -108 2145 -50 2157
rect 50 2933 108 2945
rect 50 2157 62 2933
rect 96 2157 108 2933
rect 50 2145 108 2157
rect -108 1915 -50 1927
rect -108 1139 -96 1915
rect -62 1139 -50 1915
rect -108 1127 -50 1139
rect 50 1915 108 1927
rect 50 1139 62 1915
rect 96 1139 108 1915
rect 50 1127 108 1139
rect -108 897 -50 909
rect -108 121 -96 897
rect -62 121 -50 897
rect -108 109 -50 121
rect 50 897 108 909
rect 50 121 62 897
rect 96 121 108 897
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -897 -96 -121
rect -62 -897 -50 -121
rect -108 -909 -50 -897
rect 50 -121 108 -109
rect 50 -897 62 -121
rect 96 -897 108 -121
rect 50 -909 108 -897
rect -108 -1139 -50 -1127
rect -108 -1915 -96 -1139
rect -62 -1915 -50 -1139
rect -108 -1927 -50 -1915
rect 50 -1139 108 -1127
rect 50 -1915 62 -1139
rect 96 -1915 108 -1139
rect 50 -1927 108 -1915
rect -108 -2157 -50 -2145
rect -108 -2933 -96 -2157
rect -62 -2933 -50 -2157
rect -108 -2945 -50 -2933
rect 50 -2157 108 -2145
rect 50 -2933 62 -2157
rect 96 -2933 108 -2157
rect 50 -2945 108 -2933
rect -108 -3175 -50 -3163
rect -108 -3951 -96 -3175
rect -62 -3951 -50 -3175
rect -108 -3963 -50 -3951
rect 50 -3175 108 -3163
rect 50 -3951 62 -3175
rect 96 -3951 108 -3175
rect 50 -3963 108 -3951
rect -108 -4193 -50 -4181
rect -108 -4969 -96 -4193
rect -62 -4969 -50 -4193
rect -108 -4981 -50 -4969
rect 50 -4193 108 -4181
rect 50 -4969 62 -4193
rect 96 -4969 108 -4193
rect 50 -4981 108 -4969
<< mvndiffc >>
rect -96 4193 -62 4969
rect 62 4193 96 4969
rect -96 3175 -62 3951
rect 62 3175 96 3951
rect -96 2157 -62 2933
rect 62 2157 96 2933
rect -96 1139 -62 1915
rect 62 1139 96 1915
rect -96 121 -62 897
rect 62 121 96 897
rect -96 -897 -62 -121
rect 62 -897 96 -121
rect -96 -1915 -62 -1139
rect 62 -1915 96 -1139
rect -96 -2933 -62 -2157
rect 62 -2933 96 -2157
rect -96 -3951 -62 -3175
rect 62 -3951 96 -3175
rect -96 -4969 -62 -4193
rect 62 -4969 96 -4193
<< mvpsubdiff >>
rect -242 5191 242 5203
rect -242 5157 -134 5191
rect 134 5157 242 5191
rect -242 5145 242 5157
rect -242 5095 -184 5145
rect -242 -5095 -230 5095
rect -196 -5095 -184 5095
rect 184 5095 242 5145
rect -242 -5145 -184 -5095
rect 184 -5095 196 5095
rect 230 -5095 242 5095
rect 184 -5145 242 -5095
rect -242 -5157 242 -5145
rect -242 -5191 -134 -5157
rect 134 -5191 242 -5157
rect -242 -5203 242 -5191
<< mvpsubdiffcont >>
rect -134 5157 134 5191
rect -230 -5095 -196 5095
rect 196 -5095 230 5095
rect -134 -5191 134 -5157
<< poly >>
rect -50 5053 50 5069
rect -50 5019 -34 5053
rect 34 5019 50 5053
rect -50 4981 50 5019
rect -50 4143 50 4181
rect -50 4109 -34 4143
rect 34 4109 50 4143
rect -50 4093 50 4109
rect -50 4035 50 4051
rect -50 4001 -34 4035
rect 34 4001 50 4035
rect -50 3963 50 4001
rect -50 3125 50 3163
rect -50 3091 -34 3125
rect 34 3091 50 3125
rect -50 3075 50 3091
rect -50 3017 50 3033
rect -50 2983 -34 3017
rect 34 2983 50 3017
rect -50 2945 50 2983
rect -50 2107 50 2145
rect -50 2073 -34 2107
rect 34 2073 50 2107
rect -50 2057 50 2073
rect -50 1999 50 2015
rect -50 1965 -34 1999
rect 34 1965 50 1999
rect -50 1927 50 1965
rect -50 1089 50 1127
rect -50 1055 -34 1089
rect 34 1055 50 1089
rect -50 1039 50 1055
rect -50 981 50 997
rect -50 947 -34 981
rect 34 947 50 981
rect -50 909 50 947
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -947 50 -909
rect -50 -981 -34 -947
rect 34 -981 50 -947
rect -50 -997 50 -981
rect -50 -1055 50 -1039
rect -50 -1089 -34 -1055
rect 34 -1089 50 -1055
rect -50 -1127 50 -1089
rect -50 -1965 50 -1927
rect -50 -1999 -34 -1965
rect 34 -1999 50 -1965
rect -50 -2015 50 -1999
rect -50 -2073 50 -2057
rect -50 -2107 -34 -2073
rect 34 -2107 50 -2073
rect -50 -2145 50 -2107
rect -50 -2983 50 -2945
rect -50 -3017 -34 -2983
rect 34 -3017 50 -2983
rect -50 -3033 50 -3017
rect -50 -3091 50 -3075
rect -50 -3125 -34 -3091
rect 34 -3125 50 -3091
rect -50 -3163 50 -3125
rect -50 -4001 50 -3963
rect -50 -4035 -34 -4001
rect 34 -4035 50 -4001
rect -50 -4051 50 -4035
rect -50 -4109 50 -4093
rect -50 -4143 -34 -4109
rect 34 -4143 50 -4109
rect -50 -4181 50 -4143
rect -50 -5019 50 -4981
rect -50 -5053 -34 -5019
rect 34 -5053 50 -5019
rect -50 -5069 50 -5053
<< polycont >>
rect -34 5019 34 5053
rect -34 4109 34 4143
rect -34 4001 34 4035
rect -34 3091 34 3125
rect -34 2983 34 3017
rect -34 2073 34 2107
rect -34 1965 34 1999
rect -34 1055 34 1089
rect -34 947 34 981
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -981 34 -947
rect -34 -1089 34 -1055
rect -34 -1999 34 -1965
rect -34 -2107 34 -2073
rect -34 -3017 34 -2983
rect -34 -3125 34 -3091
rect -34 -4035 34 -4001
rect -34 -4143 34 -4109
rect -34 -5053 34 -5019
<< locali >>
rect -230 5157 -134 5191
rect 134 5157 230 5191
rect -230 5095 -196 5157
rect 196 5095 230 5157
rect -50 5019 -34 5053
rect 34 5019 50 5053
rect -96 4969 -62 4985
rect -96 4177 -62 4193
rect 62 4969 96 4985
rect 62 4177 96 4193
rect -50 4109 -34 4143
rect 34 4109 50 4143
rect -50 4001 -34 4035
rect 34 4001 50 4035
rect -96 3951 -62 3967
rect -96 3159 -62 3175
rect 62 3951 96 3967
rect 62 3159 96 3175
rect -50 3091 -34 3125
rect 34 3091 50 3125
rect -50 2983 -34 3017
rect 34 2983 50 3017
rect -96 2933 -62 2949
rect -96 2141 -62 2157
rect 62 2933 96 2949
rect 62 2141 96 2157
rect -50 2073 -34 2107
rect 34 2073 50 2107
rect -50 1965 -34 1999
rect 34 1965 50 1999
rect -96 1915 -62 1931
rect -96 1123 -62 1139
rect 62 1915 96 1931
rect 62 1123 96 1139
rect -50 1055 -34 1089
rect 34 1055 50 1089
rect -50 947 -34 981
rect 34 947 50 981
rect -96 897 -62 913
rect -96 105 -62 121
rect 62 897 96 913
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -913 -62 -897
rect 62 -121 96 -105
rect 62 -913 96 -897
rect -50 -981 -34 -947
rect 34 -981 50 -947
rect -50 -1089 -34 -1055
rect 34 -1089 50 -1055
rect -96 -1139 -62 -1123
rect -96 -1931 -62 -1915
rect 62 -1139 96 -1123
rect 62 -1931 96 -1915
rect -50 -1999 -34 -1965
rect 34 -1999 50 -1965
rect -50 -2107 -34 -2073
rect 34 -2107 50 -2073
rect -96 -2157 -62 -2141
rect -96 -2949 -62 -2933
rect 62 -2157 96 -2141
rect 62 -2949 96 -2933
rect -50 -3017 -34 -2983
rect 34 -3017 50 -2983
rect -50 -3125 -34 -3091
rect 34 -3125 50 -3091
rect -96 -3175 -62 -3159
rect -96 -3967 -62 -3951
rect 62 -3175 96 -3159
rect 62 -3967 96 -3951
rect -50 -4035 -34 -4001
rect 34 -4035 50 -4001
rect -50 -4143 -34 -4109
rect 34 -4143 50 -4109
rect -96 -4193 -62 -4177
rect -96 -4985 -62 -4969
rect 62 -4193 96 -4177
rect 62 -4985 96 -4969
rect -50 -5053 -34 -5019
rect 34 -5053 50 -5019
rect -230 -5157 -196 -5095
rect 196 -5157 230 -5095
rect -230 -5191 -134 -5157
rect 134 -5191 230 -5157
<< viali >>
rect -34 5019 34 5053
rect -96 4193 -62 4969
rect 62 4193 96 4969
rect -34 4109 34 4143
rect -34 4001 34 4035
rect -96 3175 -62 3951
rect 62 3175 96 3951
rect -34 3091 34 3125
rect -34 2983 34 3017
rect -96 2157 -62 2933
rect 62 2157 96 2933
rect -34 2073 34 2107
rect -34 1965 34 1999
rect -96 1139 -62 1915
rect 62 1139 96 1915
rect -34 1055 34 1089
rect -34 947 34 981
rect -96 121 -62 897
rect 62 121 96 897
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -897 -62 -121
rect 62 -897 96 -121
rect -34 -981 34 -947
rect -34 -1089 34 -1055
rect -96 -1915 -62 -1139
rect 62 -1915 96 -1139
rect -34 -1999 34 -1965
rect -34 -2107 34 -2073
rect -96 -2933 -62 -2157
rect 62 -2933 96 -2157
rect -34 -3017 34 -2983
rect -34 -3125 34 -3091
rect -96 -3951 -62 -3175
rect 62 -3951 96 -3175
rect -34 -4035 34 -4001
rect -34 -4143 34 -4109
rect -96 -4969 -62 -4193
rect 62 -4969 96 -4193
rect -34 -5053 34 -5019
<< metal1 >>
rect -46 5053 46 5059
rect -46 5019 -34 5053
rect 34 5019 46 5053
rect -46 5013 46 5019
rect -102 4969 -56 4981
rect -102 4193 -96 4969
rect -62 4193 -56 4969
rect -102 4181 -56 4193
rect 56 4969 102 4981
rect 56 4193 62 4969
rect 96 4193 102 4969
rect 56 4181 102 4193
rect -46 4143 46 4149
rect -46 4109 -34 4143
rect 34 4109 46 4143
rect -46 4103 46 4109
rect -46 4035 46 4041
rect -46 4001 -34 4035
rect 34 4001 46 4035
rect -46 3995 46 4001
rect -102 3951 -56 3963
rect -102 3175 -96 3951
rect -62 3175 -56 3951
rect -102 3163 -56 3175
rect 56 3951 102 3963
rect 56 3175 62 3951
rect 96 3175 102 3951
rect 56 3163 102 3175
rect -46 3125 46 3131
rect -46 3091 -34 3125
rect 34 3091 46 3125
rect -46 3085 46 3091
rect -46 3017 46 3023
rect -46 2983 -34 3017
rect 34 2983 46 3017
rect -46 2977 46 2983
rect -102 2933 -56 2945
rect -102 2157 -96 2933
rect -62 2157 -56 2933
rect -102 2145 -56 2157
rect 56 2933 102 2945
rect 56 2157 62 2933
rect 96 2157 102 2933
rect 56 2145 102 2157
rect -46 2107 46 2113
rect -46 2073 -34 2107
rect 34 2073 46 2107
rect -46 2067 46 2073
rect -46 1999 46 2005
rect -46 1965 -34 1999
rect 34 1965 46 1999
rect -46 1959 46 1965
rect -102 1915 -56 1927
rect -102 1139 -96 1915
rect -62 1139 -56 1915
rect -102 1127 -56 1139
rect 56 1915 102 1927
rect 56 1139 62 1915
rect 96 1139 102 1915
rect 56 1127 102 1139
rect -46 1089 46 1095
rect -46 1055 -34 1089
rect 34 1055 46 1089
rect -46 1049 46 1055
rect -46 981 46 987
rect -46 947 -34 981
rect 34 947 46 981
rect -46 941 46 947
rect -102 897 -56 909
rect -102 121 -96 897
rect -62 121 -56 897
rect -102 109 -56 121
rect 56 897 102 909
rect 56 121 62 897
rect 96 121 102 897
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -897 -96 -121
rect -62 -897 -56 -121
rect -102 -909 -56 -897
rect 56 -121 102 -109
rect 56 -897 62 -121
rect 96 -897 102 -121
rect 56 -909 102 -897
rect -46 -947 46 -941
rect -46 -981 -34 -947
rect 34 -981 46 -947
rect -46 -987 46 -981
rect -46 -1055 46 -1049
rect -46 -1089 -34 -1055
rect 34 -1089 46 -1055
rect -46 -1095 46 -1089
rect -102 -1139 -56 -1127
rect -102 -1915 -96 -1139
rect -62 -1915 -56 -1139
rect -102 -1927 -56 -1915
rect 56 -1139 102 -1127
rect 56 -1915 62 -1139
rect 96 -1915 102 -1139
rect 56 -1927 102 -1915
rect -46 -1965 46 -1959
rect -46 -1999 -34 -1965
rect 34 -1999 46 -1965
rect -46 -2005 46 -1999
rect -46 -2073 46 -2067
rect -46 -2107 -34 -2073
rect 34 -2107 46 -2073
rect -46 -2113 46 -2107
rect -102 -2157 -56 -2145
rect -102 -2933 -96 -2157
rect -62 -2933 -56 -2157
rect -102 -2945 -56 -2933
rect 56 -2157 102 -2145
rect 56 -2933 62 -2157
rect 96 -2933 102 -2157
rect 56 -2945 102 -2933
rect -46 -2983 46 -2977
rect -46 -3017 -34 -2983
rect 34 -3017 46 -2983
rect -46 -3023 46 -3017
rect -46 -3091 46 -3085
rect -46 -3125 -34 -3091
rect 34 -3125 46 -3091
rect -46 -3131 46 -3125
rect -102 -3175 -56 -3163
rect -102 -3951 -96 -3175
rect -62 -3951 -56 -3175
rect -102 -3963 -56 -3951
rect 56 -3175 102 -3163
rect 56 -3951 62 -3175
rect 96 -3951 102 -3175
rect 56 -3963 102 -3951
rect -46 -4001 46 -3995
rect -46 -4035 -34 -4001
rect 34 -4035 46 -4001
rect -46 -4041 46 -4035
rect -46 -4109 46 -4103
rect -46 -4143 -34 -4109
rect 34 -4143 46 -4109
rect -46 -4149 46 -4143
rect -102 -4193 -56 -4181
rect -102 -4969 -96 -4193
rect -62 -4969 -56 -4193
rect -102 -4981 -56 -4969
rect 56 -4193 102 -4181
rect 56 -4969 62 -4193
rect 96 -4969 102 -4193
rect 56 -4981 102 -4969
rect -46 -5019 46 -5013
rect -46 -5053 -34 -5019
rect 34 -5053 46 -5019
rect -46 -5059 46 -5053
<< properties >>
string FIXED_BBOX -213 -5174 213 5174
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 0.5 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
