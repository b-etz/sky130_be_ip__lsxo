magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
use sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B  sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B_0
timestamp 1712071977
transform 1 0 2529 0 1 -1234
box -357 -558 357 558
use sky130_fd_pr__nfet_01v8_69TQ3K  XM1
timestamp 1712071977
transform 1 0 897 0 1 -2007
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_3HMWVM  XM2
timestamp 1712071977
transform 1 0 937 0 1 -1052
box -296 -319 296 319
use sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B  XM3
timestamp 1712071977
transform 1 0 1822 0 1 -1234
box -357 -558 357 558
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM5
timestamp 1712071977
transform 1 0 1411 0 1 83
box -658 -397 658 397
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM6
timestamp 1712071977
transform 1 0 2537 0 1 83
box -658 -397 658 397
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 128 0 0 0 avdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 128 0 0 0 dvdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 128 0 0 0 out
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 128 0 0 0 out_b
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 128 0 0 0 in
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 128 0 0 0 dvss
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 128 0 0 0 avss
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 128 0 0 0 in_b
port 7 nsew
<< end >>
