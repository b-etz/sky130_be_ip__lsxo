magic
tech sky130A
magscale 1 2
timestamp 1713225924
<< metal3 >>
rect -2386 7200 2092 11680
rect -2386 2480 2092 6960
rect -2386 -2240 2092 2240
rect -2386 -6960 2092 -2480
rect -2386 -11678 2092 -7200
rect -2386 -11680 -286 -11678
rect 12 -11680 2092 -11678
<< mimcap >>
rect -2346 11600 2054 11640
rect -2346 7280 -2306 11600
rect 2014 7280 2054 11600
rect -2346 7240 2054 7280
rect -2346 6880 2054 6920
rect -2346 2560 -2306 6880
rect 2014 2560 2054 6880
rect -2346 2520 2054 2560
rect -2346 2160 2054 2200
rect -2346 -2160 -2306 2160
rect 2014 -2160 2054 2160
rect -2346 -2200 2054 -2160
rect -2346 -2560 2054 -2520
rect -2346 -6880 -2306 -2560
rect 2014 -6880 2054 -2560
rect -2346 -6920 2054 -6880
rect -2346 -7280 2054 -7240
rect -2346 -11600 -2306 -7280
rect 2014 -11600 2054 -7280
rect -2346 -11640 2054 -11600
<< mimcapcontact >>
rect -2306 7280 2014 11600
rect -2306 2560 2014 6880
rect -2306 -2160 2014 2160
rect -2306 -6880 2014 -2560
rect -2306 -11600 2014 -7280
<< metal4 >>
rect -198 11601 -94 11684
rect -2307 11600 2015 11601
rect -2307 7280 -2306 11600
rect 2014 7280 2015 11600
rect -2307 7279 2015 7280
rect -198 6881 -94 7279
rect -2307 6880 2015 6881
rect -2307 2560 -2306 6880
rect 2014 2560 2015 6880
rect -2307 2559 2015 2560
rect -198 2161 -94 2559
rect -2307 2160 2015 2161
rect -2307 -2160 -2306 2160
rect 2014 -2160 2015 2160
rect -2307 -2161 2015 -2160
rect -198 -2559 -94 -2161
rect -2307 -2560 2015 -2559
rect -2307 -6880 -2306 -2560
rect 2014 -6880 2015 -2560
rect -2307 -6881 2015 -6880
rect -198 -7279 -94 -6881
rect -2307 -7280 2015 -7279
rect -2307 -11600 -2306 -7280
rect 2014 -11600 2015 -7280
rect -2307 -11601 2015 -11600
rect -198 -11678 -94 -11601
<< properties >>
string FIXED_BBOX -2386 7200 2094 11680
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 22 l 22 val 984.72 carea 2.00 cperi 0.19 nx 1 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
