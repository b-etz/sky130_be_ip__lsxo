magic
tech sky130A
magscale 1 2
timestamp 1712878565
<< pwell >>
rect -2359 -10982 2359 10982
<< psubdiff >>
rect -2323 10912 -2227 10946
rect 2227 10912 2323 10946
rect -2323 10850 -2289 10912
rect 2289 10850 2323 10912
rect -2323 -10912 -2289 -10850
rect 2289 -10912 2323 -10850
rect -2323 -10946 -2227 -10912
rect 2227 -10946 2323 -10912
<< psubdiffcont >>
rect -2227 10912 2227 10946
rect -2323 -10850 -2289 10850
rect 2289 -10850 2323 10850
rect -2227 -10946 2227 -10912
<< xpolycontact >>
rect -2193 10384 -2123 10816
rect -2193 -10816 -2123 -10384
rect -2027 10384 -1957 10816
rect -2027 -10816 -1957 -10384
rect -1861 10384 -1791 10816
rect -1861 -10816 -1791 -10384
rect -1695 10384 -1625 10816
rect -1695 -10816 -1625 -10384
rect -1529 10384 -1459 10816
rect -1529 -10816 -1459 -10384
rect -1363 10384 -1293 10816
rect -1363 -10816 -1293 -10384
rect -1197 10384 -1127 10816
rect -1197 -10816 -1127 -10384
rect -1031 10384 -961 10816
rect -1031 -10816 -961 -10384
rect -865 10384 -795 10816
rect -865 -10816 -795 -10384
rect -699 10384 -629 10816
rect -699 -10816 -629 -10384
rect -533 10384 -463 10816
rect -533 -10816 -463 -10384
rect -367 10384 -297 10816
rect -367 -10816 -297 -10384
rect -201 10384 -131 10816
rect -201 -10816 -131 -10384
rect -35 10384 35 10816
rect -35 -10816 35 -10384
rect 131 10384 201 10816
rect 131 -10816 201 -10384
rect 297 10384 367 10816
rect 297 -10816 367 -10384
rect 463 10384 533 10816
rect 463 -10816 533 -10384
rect 629 10384 699 10816
rect 629 -10816 699 -10384
rect 795 10384 865 10816
rect 795 -10816 865 -10384
rect 961 10384 1031 10816
rect 961 -10816 1031 -10384
rect 1127 10384 1197 10816
rect 1127 -10816 1197 -10384
rect 1293 10384 1363 10816
rect 1293 -10816 1363 -10384
rect 1459 10384 1529 10816
rect 1459 -10816 1529 -10384
rect 1625 10384 1695 10816
rect 1625 -10816 1695 -10384
rect 1791 10384 1861 10816
rect 1791 -10816 1861 -10384
rect 1957 10384 2027 10816
rect 1957 -10816 2027 -10384
rect 2123 10384 2193 10816
rect 2123 -10816 2193 -10384
<< xpolyres >>
rect -2193 -10384 -2123 10384
rect -2027 -10384 -1957 10384
rect -1861 -10384 -1791 10384
rect -1695 -10384 -1625 10384
rect -1529 -10384 -1459 10384
rect -1363 -10384 -1293 10384
rect -1197 -10384 -1127 10384
rect -1031 -10384 -961 10384
rect -865 -10384 -795 10384
rect -699 -10384 -629 10384
rect -533 -10384 -463 10384
rect -367 -10384 -297 10384
rect -201 -10384 -131 10384
rect -35 -10384 35 10384
rect 131 -10384 201 10384
rect 297 -10384 367 10384
rect 463 -10384 533 10384
rect 629 -10384 699 10384
rect 795 -10384 865 10384
rect 961 -10384 1031 10384
rect 1127 -10384 1197 10384
rect 1293 -10384 1363 10384
rect 1459 -10384 1529 10384
rect 1625 -10384 1695 10384
rect 1791 -10384 1861 10384
rect 1957 -10384 2027 10384
rect 2123 -10384 2193 10384
<< locali >>
rect -2323 10912 -2227 10946
rect 2227 10912 2323 10946
rect -2323 10850 -2289 10912
rect 2289 10850 2323 10912
rect -2323 -10912 -2289 -10850
rect 2289 -10912 2323 -10850
rect -2323 -10946 -2227 -10912
rect 2227 -10946 2323 -10912
<< viali >>
rect -2177 10401 -2139 10798
rect -2011 10401 -1973 10798
rect -1845 10401 -1807 10798
rect -1679 10401 -1641 10798
rect -1513 10401 -1475 10798
rect -1347 10401 -1309 10798
rect -1181 10401 -1143 10798
rect -1015 10401 -977 10798
rect -849 10401 -811 10798
rect -683 10401 -645 10798
rect -517 10401 -479 10798
rect -351 10401 -313 10798
rect -185 10401 -147 10798
rect -19 10401 19 10798
rect 147 10401 185 10798
rect 313 10401 351 10798
rect 479 10401 517 10798
rect 645 10401 683 10798
rect 811 10401 849 10798
rect 977 10401 1015 10798
rect 1143 10401 1181 10798
rect 1309 10401 1347 10798
rect 1475 10401 1513 10798
rect 1641 10401 1679 10798
rect 1807 10401 1845 10798
rect 1973 10401 2011 10798
rect 2139 10401 2177 10798
rect -2177 -10798 -2139 -10401
rect -2011 -10798 -1973 -10401
rect -1845 -10798 -1807 -10401
rect -1679 -10798 -1641 -10401
rect -1513 -10798 -1475 -10401
rect -1347 -10798 -1309 -10401
rect -1181 -10798 -1143 -10401
rect -1015 -10798 -977 -10401
rect -849 -10798 -811 -10401
rect -683 -10798 -645 -10401
rect -517 -10798 -479 -10401
rect -351 -10798 -313 -10401
rect -185 -10798 -147 -10401
rect -19 -10798 19 -10401
rect 147 -10798 185 -10401
rect 313 -10798 351 -10401
rect 479 -10798 517 -10401
rect 645 -10798 683 -10401
rect 811 -10798 849 -10401
rect 977 -10798 1015 -10401
rect 1143 -10798 1181 -10401
rect 1309 -10798 1347 -10401
rect 1475 -10798 1513 -10401
rect 1641 -10798 1679 -10401
rect 1807 -10798 1845 -10401
rect 1973 -10798 2011 -10401
rect 2139 -10798 2177 -10401
<< metal1 >>
rect -2183 10798 -2133 10810
rect -2183 10401 -2177 10798
rect -2139 10401 -2133 10798
rect -2183 10389 -2133 10401
rect -2017 10798 -1967 10810
rect -2017 10401 -2011 10798
rect -1973 10401 -1967 10798
rect -2017 10389 -1967 10401
rect -1851 10798 -1801 10810
rect -1851 10401 -1845 10798
rect -1807 10401 -1801 10798
rect -1851 10389 -1801 10401
rect -1685 10798 -1635 10810
rect -1685 10401 -1679 10798
rect -1641 10401 -1635 10798
rect -1685 10389 -1635 10401
rect -1519 10798 -1469 10810
rect -1519 10401 -1513 10798
rect -1475 10401 -1469 10798
rect -1519 10389 -1469 10401
rect -1353 10798 -1303 10810
rect -1353 10401 -1347 10798
rect -1309 10401 -1303 10798
rect -1353 10389 -1303 10401
rect -1187 10798 -1137 10810
rect -1187 10401 -1181 10798
rect -1143 10401 -1137 10798
rect -1187 10389 -1137 10401
rect -1021 10798 -971 10810
rect -1021 10401 -1015 10798
rect -977 10401 -971 10798
rect -1021 10389 -971 10401
rect -855 10798 -805 10810
rect -855 10401 -849 10798
rect -811 10401 -805 10798
rect -855 10389 -805 10401
rect -689 10798 -639 10810
rect -689 10401 -683 10798
rect -645 10401 -639 10798
rect -689 10389 -639 10401
rect -523 10798 -473 10810
rect -523 10401 -517 10798
rect -479 10401 -473 10798
rect -523 10389 -473 10401
rect -357 10798 -307 10810
rect -357 10401 -351 10798
rect -313 10401 -307 10798
rect -357 10389 -307 10401
rect -191 10798 -141 10810
rect -191 10401 -185 10798
rect -147 10401 -141 10798
rect -191 10389 -141 10401
rect -25 10798 25 10810
rect -25 10401 -19 10798
rect 19 10401 25 10798
rect -25 10389 25 10401
rect 141 10798 191 10810
rect 141 10401 147 10798
rect 185 10401 191 10798
rect 141 10389 191 10401
rect 307 10798 357 10810
rect 307 10401 313 10798
rect 351 10401 357 10798
rect 307 10389 357 10401
rect 473 10798 523 10810
rect 473 10401 479 10798
rect 517 10401 523 10798
rect 473 10389 523 10401
rect 639 10798 689 10810
rect 639 10401 645 10798
rect 683 10401 689 10798
rect 639 10389 689 10401
rect 805 10798 855 10810
rect 805 10401 811 10798
rect 849 10401 855 10798
rect 805 10389 855 10401
rect 971 10798 1021 10810
rect 971 10401 977 10798
rect 1015 10401 1021 10798
rect 971 10389 1021 10401
rect 1137 10798 1187 10810
rect 1137 10401 1143 10798
rect 1181 10401 1187 10798
rect 1137 10389 1187 10401
rect 1303 10798 1353 10810
rect 1303 10401 1309 10798
rect 1347 10401 1353 10798
rect 1303 10389 1353 10401
rect 1469 10798 1519 10810
rect 1469 10401 1475 10798
rect 1513 10401 1519 10798
rect 1469 10389 1519 10401
rect 1635 10798 1685 10810
rect 1635 10401 1641 10798
rect 1679 10401 1685 10798
rect 1635 10389 1685 10401
rect 1801 10798 1851 10810
rect 1801 10401 1807 10798
rect 1845 10401 1851 10798
rect 1801 10389 1851 10401
rect 1967 10798 2017 10810
rect 1967 10401 1973 10798
rect 2011 10401 2017 10798
rect 1967 10389 2017 10401
rect 2133 10798 2183 10810
rect 2133 10401 2139 10798
rect 2177 10401 2183 10798
rect 2133 10389 2183 10401
rect -2183 -10401 -2133 -10389
rect -2183 -10798 -2177 -10401
rect -2139 -10798 -2133 -10401
rect -2183 -10810 -2133 -10798
rect -2017 -10401 -1967 -10389
rect -2017 -10798 -2011 -10401
rect -1973 -10798 -1967 -10401
rect -2017 -10810 -1967 -10798
rect -1851 -10401 -1801 -10389
rect -1851 -10798 -1845 -10401
rect -1807 -10798 -1801 -10401
rect -1851 -10810 -1801 -10798
rect -1685 -10401 -1635 -10389
rect -1685 -10798 -1679 -10401
rect -1641 -10798 -1635 -10401
rect -1685 -10810 -1635 -10798
rect -1519 -10401 -1469 -10389
rect -1519 -10798 -1513 -10401
rect -1475 -10798 -1469 -10401
rect -1519 -10810 -1469 -10798
rect -1353 -10401 -1303 -10389
rect -1353 -10798 -1347 -10401
rect -1309 -10798 -1303 -10401
rect -1353 -10810 -1303 -10798
rect -1187 -10401 -1137 -10389
rect -1187 -10798 -1181 -10401
rect -1143 -10798 -1137 -10401
rect -1187 -10810 -1137 -10798
rect -1021 -10401 -971 -10389
rect -1021 -10798 -1015 -10401
rect -977 -10798 -971 -10401
rect -1021 -10810 -971 -10798
rect -855 -10401 -805 -10389
rect -855 -10798 -849 -10401
rect -811 -10798 -805 -10401
rect -855 -10810 -805 -10798
rect -689 -10401 -639 -10389
rect -689 -10798 -683 -10401
rect -645 -10798 -639 -10401
rect -689 -10810 -639 -10798
rect -523 -10401 -473 -10389
rect -523 -10798 -517 -10401
rect -479 -10798 -473 -10401
rect -523 -10810 -473 -10798
rect -357 -10401 -307 -10389
rect -357 -10798 -351 -10401
rect -313 -10798 -307 -10401
rect -357 -10810 -307 -10798
rect -191 -10401 -141 -10389
rect -191 -10798 -185 -10401
rect -147 -10798 -141 -10401
rect -191 -10810 -141 -10798
rect -25 -10401 25 -10389
rect -25 -10798 -19 -10401
rect 19 -10798 25 -10401
rect -25 -10810 25 -10798
rect 141 -10401 191 -10389
rect 141 -10798 147 -10401
rect 185 -10798 191 -10401
rect 141 -10810 191 -10798
rect 307 -10401 357 -10389
rect 307 -10798 313 -10401
rect 351 -10798 357 -10401
rect 307 -10810 357 -10798
rect 473 -10401 523 -10389
rect 473 -10798 479 -10401
rect 517 -10798 523 -10401
rect 473 -10810 523 -10798
rect 639 -10401 689 -10389
rect 639 -10798 645 -10401
rect 683 -10798 689 -10401
rect 639 -10810 689 -10798
rect 805 -10401 855 -10389
rect 805 -10798 811 -10401
rect 849 -10798 855 -10401
rect 805 -10810 855 -10798
rect 971 -10401 1021 -10389
rect 971 -10798 977 -10401
rect 1015 -10798 1021 -10401
rect 971 -10810 1021 -10798
rect 1137 -10401 1187 -10389
rect 1137 -10798 1143 -10401
rect 1181 -10798 1187 -10401
rect 1137 -10810 1187 -10798
rect 1303 -10401 1353 -10389
rect 1303 -10798 1309 -10401
rect 1347 -10798 1353 -10401
rect 1303 -10810 1353 -10798
rect 1469 -10401 1519 -10389
rect 1469 -10798 1475 -10401
rect 1513 -10798 1519 -10401
rect 1469 -10810 1519 -10798
rect 1635 -10401 1685 -10389
rect 1635 -10798 1641 -10401
rect 1679 -10798 1685 -10401
rect 1635 -10810 1685 -10798
rect 1801 -10401 1851 -10389
rect 1801 -10798 1807 -10401
rect 1845 -10798 1851 -10401
rect 1801 -10810 1851 -10798
rect 1967 -10401 2017 -10389
rect 1967 -10798 1973 -10401
rect 2011 -10798 2017 -10401
rect 1967 -10810 2017 -10798
rect 2133 -10401 2183 -10389
rect 2133 -10798 2139 -10401
rect 2177 -10798 2183 -10401
rect 2133 -10810 2183 -10798
<< properties >>
string FIXED_BBOX -2306 -10929 2306 10929
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 104.0 m 1 nx 27 wmin 0.350 lmin 0.50 rho 2000 val 595.361k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
