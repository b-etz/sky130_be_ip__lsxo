magic
tech sky130A
magscale 1 2
timestamp 1712954292
<< dnwell >>
rect 1932 -9000 6418 -3442
rect 8780 -10312 25248 -4220
rect 1706 -23624 25490 -11618
<< nwell >>
rect 1852 -3648 6498 -3362
rect 1852 -8794 2138 -3648
rect 6212 -8794 6498 -3648
rect 1852 -9080 6498 -8794
rect 8700 -4426 25328 -4140
rect 8700 -10106 8986 -4426
rect 25042 -10106 25328 -4426
rect 8700 -10392 25328 -10106
rect 1626 -11824 25570 -11538
rect 1626 -23418 1912 -11824
rect 25284 -23418 25570 -11824
rect 1626 -23704 25570 -23418
<< nsubdiff >>
rect 1889 -3419 6461 -3399
rect 1889 -3453 1969 -3419
rect 6381 -3453 6461 -3419
rect 1889 -3473 6461 -3453
rect 1889 -3479 1963 -3473
rect 1889 -8963 1909 -3479
rect 1943 -8963 1963 -3479
rect 1889 -8969 1963 -8963
rect 6387 -3479 6461 -3473
rect 6387 -8963 6407 -3479
rect 6441 -8963 6461 -3479
rect 6387 -8969 6461 -8963
rect 1889 -8989 6461 -8969
rect 1889 -9023 1969 -8989
rect 6381 -9023 6461 -8989
rect 1889 -9043 6461 -9023
rect 8737 -4197 25291 -4177
rect 8737 -4231 8817 -4197
rect 25211 -4231 25291 -4197
rect 8737 -4251 25291 -4231
rect 8737 -4257 8811 -4251
rect 8737 -10275 8757 -4257
rect 8791 -10275 8811 -4257
rect 8737 -10281 8811 -10275
rect 25217 -4257 25291 -4251
rect 25217 -10275 25237 -4257
rect 25271 -10275 25291 -4257
rect 25217 -10281 25291 -10275
rect 8737 -10301 25291 -10281
rect 8737 -10335 8817 -10301
rect 25211 -10335 25291 -10301
rect 8737 -10355 25291 -10335
rect 1663 -11595 25533 -11575
rect 1663 -11629 1743 -11595
rect 25453 -11629 25533 -11595
rect 1663 -11649 25533 -11629
rect 1663 -11655 1737 -11649
rect 1663 -23587 1683 -11655
rect 1717 -23587 1737 -11655
rect 1663 -23593 1737 -23587
rect 25459 -11655 25533 -11649
rect 25459 -23587 25479 -11655
rect 25513 -23587 25533 -11655
rect 25459 -23593 25533 -23587
rect 1663 -23613 25533 -23593
rect 1663 -23647 1743 -23613
rect 25453 -23647 25533 -23613
rect 1663 -23667 25533 -23647
<< nsubdiffcont >>
rect 1969 -3453 6381 -3419
rect 1909 -8963 1943 -3479
rect 6407 -8963 6441 -3479
rect 1969 -9023 6381 -8989
rect 8817 -4231 25211 -4197
rect 8757 -10275 8791 -4257
rect 25237 -10275 25271 -4257
rect 8817 -10335 25211 -10301
rect 1743 -11629 25453 -11595
rect 1683 -23587 1717 -11655
rect 25479 -23587 25513 -11655
rect 1743 -23647 25453 -23613
<< locali >>
rect 1909 -3453 1969 -3419
rect 6381 -3453 6441 -3419
rect 1909 -3479 1943 -3453
rect 6407 -3479 6441 -3453
rect 3872 -7142 4600 -7134
rect 2500 -7152 3228 -7142
rect 2500 -7216 2512 -7152
rect 3872 -7208 3888 -7142
rect 4588 -7208 4600 -7142
rect 2406 -7266 2526 -7254
rect 2406 -8042 2420 -7266
rect 2512 -8042 2526 -7266
rect 2406 -8054 2526 -8042
rect 2564 -7266 2684 -7254
rect 2564 -8042 2578 -7266
rect 2670 -8042 2684 -7266
rect 2564 -8054 2684 -8042
rect 2722 -7266 2842 -7254
rect 2722 -8042 2736 -7266
rect 2828 -8042 2842 -7266
rect 2722 -8054 2842 -8042
rect 2880 -7266 3000 -7254
rect 2880 -8042 2894 -7266
rect 2986 -8042 3000 -7266
rect 2880 -8054 3000 -8042
rect 3036 -7266 3156 -7254
rect 3036 -8042 3050 -7266
rect 3142 -8042 3156 -7266
rect 3036 -8054 3156 -8042
rect 3196 -7266 3316 -7254
rect 3196 -8042 3210 -7266
rect 3302 -8042 3316 -7266
rect 3196 -8054 3316 -8042
rect 3782 -7266 3902 -7254
rect 3782 -8044 3796 -7266
rect 3888 -8044 3902 -7266
rect 3782 -8054 3902 -8044
rect 3940 -7266 4060 -7254
rect 3940 -8044 3954 -7266
rect 4046 -8044 4060 -7266
rect 3940 -8054 4060 -8044
rect 4098 -7266 4218 -7254
rect 4098 -8044 4112 -7266
rect 4204 -8044 4218 -7266
rect 4098 -8054 4218 -8044
rect 4256 -7266 4376 -7254
rect 4256 -8044 4270 -7266
rect 4362 -8044 4376 -7266
rect 4256 -8054 4376 -8044
rect 4414 -7266 4534 -7254
rect 4414 -8044 4428 -7266
rect 4520 -8044 4534 -7266
rect 4414 -8054 4534 -8044
rect 4572 -7266 4692 -7254
rect 4572 -8044 4586 -7266
rect 4678 -8044 4692 -7266
rect 4572 -8054 4692 -8044
rect 2500 -8158 2512 -8092
rect 3212 -8158 3228 -8092
rect 2500 -8166 3228 -8158
rect 3872 -8168 3888 -8102
rect 4588 -8168 4600 -8102
rect 3872 -8176 4600 -8168
rect 1909 -8989 1943 -8963
rect 6407 -8989 6441 -8963
rect 1909 -9023 1969 -8989
rect 6381 -9023 6441 -8989
rect 8757 -4231 8817 -4197
rect 25211 -4231 25271 -4197
rect 8757 -4257 8791 -4231
rect 8757 -10301 8791 -10275
rect 25237 -4257 25271 -4231
rect 25237 -10301 25271 -10275
rect 8757 -10335 8817 -10301
rect 25211 -10335 25271 -10301
rect 1683 -11629 1743 -11595
rect 25453 -11629 25513 -11595
rect 1683 -11655 1717 -11629
rect 1683 -23613 1717 -23587
rect 25479 -11655 25513 -11629
rect 25479 -23613 25513 -23587
rect 1683 -23647 1743 -23613
rect 25453 -23647 25513 -23613
<< viali >>
rect 2512 -7216 3230 -7152
rect 3888 -7208 4588 -7142
rect 2420 -8042 2512 -7266
rect 2578 -8042 2670 -7266
rect 2736 -8042 2828 -7266
rect 2894 -8042 2986 -7266
rect 3050 -8042 3142 -7266
rect 3210 -8042 3302 -7266
rect 3796 -8044 3888 -7266
rect 3954 -8044 4046 -7266
rect 4112 -8044 4204 -7266
rect 4270 -8044 4362 -7266
rect 4428 -8044 4520 -7266
rect 4586 -8044 4678 -7266
rect 2512 -8158 3212 -8092
rect 3888 -8168 4588 -8102
<< metal1 >>
rect 3264 -872 3464 -672
rect 4922 -872 5122 -672
rect 1890 -1200 2090 -1000
rect 2242 -1202 2442 -1002
rect 7066 -1128 7266 -928
rect 9806 -958 10006 -758
rect 11378 -950 11578 -750
rect 23862 -1102 24062 -902
rect 3364 -7142 3370 -6962
rect 2500 -7152 3370 -7142
rect 2500 -7216 2512 -7152
rect 3230 -7216 3370 -7152
rect 2500 -7222 3370 -7216
rect 3478 -7222 3484 -6962
rect 3614 -7214 3620 -6954
rect 3728 -7134 3734 -6954
rect 3728 -7142 4600 -7134
rect 3728 -7208 3888 -7142
rect 4588 -7208 4600 -7142
rect 3728 -7214 4600 -7208
rect 2406 -8054 2412 -7254
rect 2520 -8054 2526 -7254
rect 2564 -8054 2570 -7254
rect 2678 -8054 2684 -7254
rect 2722 -8054 2728 -7254
rect 2836 -8054 2842 -7254
rect 2880 -8054 2886 -7254
rect 2994 -8054 3000 -7254
rect 3036 -8054 3042 -7254
rect 3150 -8054 3156 -7254
rect 3196 -8054 3202 -7254
rect 3310 -8054 3316 -7254
rect 3364 -8086 3370 -7906
rect 2500 -8092 3370 -8086
rect 2500 -8158 2512 -8092
rect 3212 -8158 3370 -8092
rect 2500 -8166 3370 -8158
rect 3478 -8086 3484 -7906
rect 3478 -8166 3486 -8086
rect 3614 -8176 3620 -7916
rect 3728 -8096 3734 -7916
rect 3782 -8054 3790 -7254
rect 3894 -8054 3902 -7254
rect 3940 -8054 3946 -7254
rect 4054 -8054 4060 -7254
rect 4098 -8054 4104 -7254
rect 4212 -8054 4218 -7254
rect 4256 -8054 4262 -7254
rect 4370 -8054 4376 -7254
rect 4414 -8054 4420 -7254
rect 4528 -8054 4534 -7254
rect 4572 -8054 4578 -7254
rect 4686 -8054 4692 -7254
rect 3728 -8102 4600 -8096
rect 3728 -8168 3888 -8102
rect 4588 -8168 4600 -8102
rect 3728 -8176 4600 -8168
rect 2312 -23296 2512 -23096
rect 24708 -23294 24908 -23094
<< via1 >>
rect 3370 -7222 3478 -6962
rect 3620 -7214 3728 -6954
rect 2412 -7266 2520 -7254
rect 2412 -8042 2420 -7266
rect 2420 -8042 2512 -7266
rect 2512 -8042 2520 -7266
rect 2412 -8054 2520 -8042
rect 2570 -7266 2678 -7254
rect 2570 -8042 2578 -7266
rect 2578 -8042 2670 -7266
rect 2670 -8042 2678 -7266
rect 2570 -8054 2678 -8042
rect 2728 -7266 2836 -7254
rect 2728 -8042 2736 -7266
rect 2736 -8042 2828 -7266
rect 2828 -8042 2836 -7266
rect 2728 -8054 2836 -8042
rect 2886 -7266 2994 -7254
rect 2886 -8042 2894 -7266
rect 2894 -8042 2986 -7266
rect 2986 -8042 2994 -7266
rect 2886 -8054 2994 -8042
rect 3042 -7266 3150 -7254
rect 3042 -8042 3050 -7266
rect 3050 -8042 3142 -7266
rect 3142 -8042 3150 -7266
rect 3042 -8054 3150 -8042
rect 3202 -7266 3310 -7254
rect 3202 -8042 3210 -7266
rect 3210 -8042 3302 -7266
rect 3302 -8042 3310 -7266
rect 3202 -8054 3310 -8042
rect 3370 -8166 3478 -7906
rect 3620 -8176 3728 -7916
rect 3790 -7266 3894 -7254
rect 3790 -8044 3796 -7266
rect 3796 -8044 3888 -7266
rect 3888 -8044 3894 -7266
rect 3790 -8054 3894 -8044
rect 3946 -7266 4054 -7254
rect 3946 -8044 3954 -7266
rect 3954 -8044 4046 -7266
rect 4046 -8044 4054 -7266
rect 3946 -8054 4054 -8044
rect 4104 -7266 4212 -7254
rect 4104 -8044 4112 -7266
rect 4112 -8044 4204 -7266
rect 4204 -8044 4212 -7266
rect 4104 -8054 4212 -8044
rect 4262 -7266 4370 -7254
rect 4262 -8044 4270 -7266
rect 4270 -8044 4362 -7266
rect 4362 -8044 4370 -7266
rect 4262 -8054 4370 -8044
rect 4420 -7266 4528 -7254
rect 4420 -8044 4428 -7266
rect 4428 -8044 4520 -7266
rect 4520 -8044 4528 -7266
rect 4420 -8054 4528 -8044
rect 4578 -7266 4686 -7254
rect 4578 -8044 4586 -7266
rect 4586 -8044 4678 -7266
rect 4678 -8044 4686 -7266
rect 4578 -8054 4686 -8044
<< metal2 >>
rect 2610 -6860 3484 -6740
rect 3364 -6962 3484 -6860
rect 2406 -7174 3158 -6974
rect 2406 -7254 2526 -7174
rect 2722 -7254 2842 -7174
rect 3036 -7254 3158 -7174
rect 3364 -7222 3370 -6962
rect 3478 -7222 3484 -6962
rect 2406 -8054 2412 -7254
rect 2520 -8054 2526 -7254
rect 2564 -8054 2570 -7254
rect 2678 -8054 2684 -7254
rect 2722 -8054 2728 -7254
rect 2836 -8054 2842 -7254
rect 2880 -8054 2886 -7254
rect 2994 -8054 3000 -7254
rect 3036 -8054 3042 -7254
rect 3150 -7554 3158 -7254
rect 3150 -8054 3156 -7554
rect 3196 -8054 3202 -7254
rect 3310 -8054 3316 -7254
rect 2564 -8134 2684 -8054
rect 2880 -8134 3000 -8054
rect 3196 -8134 3316 -8054
rect 2564 -8334 3316 -8134
rect 3364 -7906 3484 -7222
rect 3364 -8166 3370 -7906
rect 3478 -8166 3484 -7906
rect 3614 -6954 3734 -6750
rect 3614 -7214 3620 -6954
rect 3728 -7214 3734 -6954
rect 3614 -7916 3734 -7214
rect 3940 -7174 4692 -6974
rect 3940 -7254 4060 -7174
rect 4256 -7254 4376 -7174
rect 4572 -7254 4692 -7174
rect 3614 -8176 3620 -7916
rect 3728 -8176 3734 -7916
rect 3782 -8054 3790 -7254
rect 3894 -8054 3902 -7254
rect 3940 -8054 3946 -7254
rect 4054 -8054 4060 -7254
rect 4098 -8054 4104 -7254
rect 4212 -8054 4218 -7254
rect 4256 -8054 4262 -7254
rect 4370 -8054 4376 -7254
rect 4414 -8054 4420 -7254
rect 4528 -8054 4534 -7254
rect 4572 -8054 4578 -7254
rect 4686 -8054 4692 -7254
rect 3782 -8134 3902 -8054
rect 4098 -8134 4218 -8054
rect 4414 -8134 4534 -8054
rect 3782 -8334 4534 -8134
use sky130_fd_pr__cap_mim_m3_1_67RTNB  amp_XC1
timestamp 1712954147
transform 0 1 12008 -1 0 -4844
box -3798 -4640 3798 4640
use sky130_fd_pr__nfet_g5v0d10v5_554GUR  amp_XM1_2
timestamp 1712954147
transform 1 0 12505 0 1 -5164
box -2031 -458 2031 458
use sky130_fd_pr__pfet_g5v0d10v5_7FQJL7  amp_XM3_5
timestamp 1712954147
transform 1 0 16085 0 1 -6505
box -1145 -697 1145 697
use sky130_fd_pr__nfet_01v8_8DG47J  amp_XM4_18
timestamp 1712954147
transform 1 0 16055 0 1 -5128
box -1083 -610 1083 610
use sky130_fd_pr__pfet_01v8_EDYT7U  amp_XM6
timestamp 1712954147
transform -1 0 18932 0 -1 -6739
box -996 -269 996 269
use sky130_fd_pr__nfet_01v8_UY343Z  amp_XM7
timestamp 1712954147
transform -1 0 18944 0 -1 -5460
box -996 -260 996 260
use sky130_fd_pr__pfet_01v8_EDYT7U  amp_XM8
timestamp 1712954147
transform 0 1 9837 -1 0 -6412
box -996 -269 996 269
use sky130_fd_pr__nfet_01v8_UY343Z  amp_XM9
timestamp 1712954147
transform 0 1 9846 -1 0 -8530
box -996 -260 996 260
use sky130_fd_pr__pfet_01v8_8D4V8N  amp_XM10_12
timestamp 1712954147
transform 1 0 21031 0 1 -6579
box -425 -383 425 383
use sky130_fd_pr__nfet_01v8_U59KY9  amp_XM11_13
timestamp 1712954147
transform 1 0 21015 0 1 -5503
box -425 -365 425 365
use sky130_fd_pr__pfet_01v8_LXFDKK  amp_XM16_17
timestamp 1712954147
transform 1 0 12485 0 1 -6453
box -1999 -683 1999 683
use sky130_fd_pr__res_xhigh_po_0p35_WHP78W  amp_XR1
timestamp 1712954147
transform 0 1 17636 -1 0 -8635
box -1363 -7182 1363 7182
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  ant_diode_ena
timestamp 1712954147
transform 1 0 2997 0 1 -857
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  ant_diode_standby
timestamp 1712954147
transform 1 0 5363 0 1 -861
box -183 -183 183 183
use sky130_fd_pr__cap_mim_m3_1_VMUSDZ  bias_XC1
timestamp 1712954147
transform 0 -1 13568 1 0 -21238
box -2386 -11800 2386 11800
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  bias_XC2
timestamp 1712954147
transform 1 0 4162 0 1 -11318
box -2186 -2040 2186 2040
use sky130_fd_pr__cap_mim_m3_1_F5PPB9  bias_XC3
timestamp 1712954147
transform 0 1 9756 -1 0 -16322
box -1986 -7840 1986 7840
use sky130_fd_pr__nfet_g5v0d10v5_QNESWN  bias_XM1_2
timestamp 1712954147
transform 0 1 20676 -1 0 -14124
box -1802 -658 1802 658
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  bias_XM5
timestamp 1712954147
transform 1 0 7432 0 1 -12402
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_H6M2KM  bias_XM6_7_8
timestamp 1712954147
transform -1 0 10760 0 -1 -12398
box -2686 -300 2686 300
use sky130_fd_pr__res_xhigh_po_0p35_M35ED8  bias_XR2
timestamp 1712954147
transform 0 1 10752 -1 0 -15996
box -2276 -8782 2276 8782
use sky130_fd_pr__res_xhigh_po_0p35_VTNT3C  bias_XR3
timestamp 1712954147
transform 0 1 10090 -1 0 -13244
box -450 -8082 450 8082
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  esd_n_xin
timestamp 1712954147
transform 1 0 2149 0 1 -22841
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  esd_n_xout
timestamp 1712954147
transform 1 0 24941 0 1 -22845
box -183 -183 183 183
use sky130_fd_pr__diode_pd2nw_05v5_K4SERG  esd_p_xin
timestamp 1712954147
transform 1 0 2919 0 1 -22979
box -321 -321 321 321
use sky130_fd_pr__diode_pd2nw_05v5_K4SERG  esd_p_xout
timestamp 1712954147
transform 1 0 24293 0 1 -22977
box -321 -321 321 321
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712954147
transform 0 -1 5522 1 0 -1300
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1712954147
transform 0 1 2814 -1 0 -1208
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712954147
transform 0 1 2814 -1 0 -1300
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x2
timestamp 1712954147
transform 0 -1 5522 -1 0 -1300
box -38 -48 314 592
use level_shift  x3
timestamp 1712954147
transform 0 1 4250 -1 0 -1190
box 652 -1950 5670 -128
use level_shift  x4
timestamp 1712954147
transform 0 -1 4086 -1 0 -1190
box 652 -1950 5670 -128
use ripl_dly_clk_buf  x7
timestamp 1712954147
transform 1 0 13462 0 1 -828
box 216 -2416 8990 -156
use sky130_fd_pr__cap_mim_m3_1_KAF84V  XC1
timestamp 1712954147
transform 0 -1 13336 1 0 -12986
box -886 -3440 886 3440
use sky130_fd_pr__cap_mim_m3_1_43FTN9  XC2
timestamp 1712954147
transform 1 0 21712 0 1 -10212
box -3798 -8120 3798 8120
use sky130_fd_pr__cap_mim_m3_1_3DMTNZ  XC3
timestamp 1712954147
transform 1 0 4198 0 1 -5146
box -2492 -2320 2492 2320
use sky130_fd_pr__cap_mim_m3_1_4HHTN9  XC4
timestamp 1712954147
transform 0 -1 11980 1 0 -10184
box -1186 -4640 1186 4640
use sky130_fd_pr__nfet_g5v0d10v5_AB4DGB  XM1
timestamp 1712954147
transform 0 1 20676 -1 0 -17063
box -1147 -658 1147 658
use sky130_fd_pr__pfet_g5v0d10v5_V6TMVM  XM2_bias_XM3_4
timestamp 1712954147
transform 0 1 22801 -1 0 -15907
box -2061 -1161 2061 1161
use sky130_fd_pr__nfet_01v8_AHZR5K  XM3
timestamp 1712954147
transform 0 1 12824 -1 0 -2652
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_HZ6WG7  XM4
timestamp 1712954147
transform 0 1 23127 -1 0 -5526
box -296 -285 296 285
use sky130_fd_pr__nfet_g5v0d10v5_ZPGQJT  XM5
timestamp 1712954147
transform -1 0 2862 0 1 -7654
box -594 -658 594 658
use sky130_fd_pr__pfet_g5v0d10v5_KLKQZ5  XM6
timestamp 1712954147
transform 1 0 4238 0 -1 -7655
box -624 -697 624 697
use sky130_fd_pr__pfet_01v8_3H68VM  XM7
timestamp 1712954147
transform 0 -1 23133 1 0 -6552
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_EDP4SU  XM8
timestamp 1712954147
transform 1 0 9853 0 1 -2647
box -957 -619 957 619
use sky130_fd_pr__pfet_g5v0d10v5_KL3SY6  XM9
timestamp 1712954147
transform -1 0 11530 0 -1 -2569
box -308 -697 308 697
use sky130_fd_pr__nfet_01v8_MLR4K3  XM11
timestamp 1712954147
transform 1 0 7747 0 1 -2664
box -957 -610 957 610
use sky130_fd_pr__res_xhigh_po_0p35_68VL2P  XR2
timestamp 1712954147
transform 0 1 13546 -1 0 -20477
box -2193 -11582 2193 11582
<< labels >>
flabel metal1 11378 -950 11578 -750 0 FreeSans 256 0 0 0 ibias
port 4 nsew
flabel metal1 7066 -1128 7266 -928 0 FreeSans 256 0 0 0 dvss
port 3 nsew
flabel metal1 9806 -958 10006 -758 0 FreeSans 256 0 0 0 dvdd
port 2 nsew
flabel metal1 2242 -1202 2442 -1002 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 1890 -1200 2090 -1000 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal1 3264 -872 3464 -672 0 FreeSans 256 0 0 0 ena
port 5 nsew
flabel metal1 4922 -872 5122 -672 0 FreeSans 256 0 0 0 standby
port 6 nsew
flabel metal1 24708 -23294 24908 -23094 0 FreeSans 256 0 0 0 xout
port 9 nsew
flabel metal1 2312 -23296 2512 -23096 0 FreeSans 256 0 0 0 xin
port 8 nsew
flabel metal1 23862 -1102 24062 -902 0 FreeSans 256 0 0 0 dout
port 7 nsew
<< end >>
