magic
tech sky130A
magscale 1 2
timestamp 1713042744
<< dnwell >>
rect 1932 -9000 6418 -3442
rect 8780 -10312 25248 -4220
rect 1706 -23624 25490 -11618
<< nwell >>
rect 1852 -3648 6498 -3362
rect 1852 -8794 2138 -3648
rect 6212 -8794 6498 -3648
rect 1852 -9080 6498 -8794
rect 8700 -4426 25328 -4140
rect 8700 -10106 8986 -4426
rect 25042 -10106 25328 -4426
rect 8700 -10392 25328 -10106
rect 1626 -11824 25570 -11538
rect 1626 -23418 1912 -11824
rect 25284 -23418 25570 -11824
rect 1626 -23704 25570 -23418
<< pwell >>
rect 10652 -5358 11064 -4958
rect 12592 -5420 12844 -4896
rect 14698 -5358 15110 -4958
<< nsubdiff >>
rect 1889 -3419 6461 -3399
rect 1889 -3453 1969 -3419
rect 6381 -3453 6461 -3419
rect 1889 -3473 6461 -3453
rect 1889 -3479 1963 -3473
rect 1889 -8963 1909 -3479
rect 1943 -8963 1963 -3479
rect 1889 -8969 1963 -8963
rect 6387 -3479 6461 -3473
rect 6387 -8963 6407 -3479
rect 6441 -8963 6461 -3479
rect 6387 -8969 6461 -8963
rect 1889 -8989 6461 -8969
rect 1889 -9023 1969 -8989
rect 6381 -9023 6461 -8989
rect 1889 -9043 6461 -9023
rect 8737 -4197 25291 -4177
rect 8737 -4231 8817 -4197
rect 25211 -4231 25291 -4197
rect 8737 -4251 25291 -4231
rect 8737 -4257 8811 -4251
rect 8737 -10275 8757 -4257
rect 8791 -10275 8811 -4257
rect 8737 -10281 8811 -10275
rect 25217 -4257 25291 -4251
rect 25217 -10275 25237 -4257
rect 25271 -10275 25291 -4257
rect 25217 -10281 25291 -10275
rect 8737 -10301 25291 -10281
rect 8737 -10335 8817 -10301
rect 25211 -10335 25291 -10301
rect 8737 -10355 25291 -10335
rect 1663 -11595 25533 -11575
rect 1663 -11629 1743 -11595
rect 25453 -11629 25533 -11595
rect 1663 -11649 25533 -11629
rect 1663 -11655 1737 -11649
rect 1663 -23587 1683 -11655
rect 1717 -23587 1737 -11655
rect 1663 -23593 1737 -23587
rect 25459 -11655 25533 -11649
rect 25459 -23587 25479 -11655
rect 25513 -23587 25533 -11655
rect 25459 -23593 25533 -23587
rect 1663 -23613 25533 -23593
rect 1663 -23647 1743 -23613
rect 25453 -23647 25533 -23613
rect 1663 -23667 25533 -23647
<< nsubdiffcont >>
rect 1969 -3453 6381 -3419
rect 1909 -8963 1943 -3479
rect 6407 -8963 6441 -3479
rect 1969 -9023 6381 -8989
rect 8817 -4231 25211 -4197
rect 8757 -10275 8791 -4257
rect 25237 -10275 25271 -4257
rect 8817 -10335 25211 -10301
rect 1743 -11629 25453 -11595
rect 1683 -23587 1717 -11655
rect 25479 -23587 25513 -11655
rect 1743 -23647 25453 -23613
<< locali >>
rect 3146 -956 3246 -946
rect 3146 -1180 3156 -956
rect 3236 -1180 3246 -956
rect 3146 -1194 3246 -1180
rect 5086 -958 5186 -948
rect 5086 -1180 5096 -958
rect 5176 -1180 5186 -958
rect 5086 -1192 5186 -1180
rect 3146 -1358 3210 -1194
rect 5120 -1350 5184 -1192
rect 11300 -2180 11474 -2164
rect 11300 -2958 11310 -2180
rect 11468 -2958 11474 -2180
rect 12600 -2212 13048 -2092
rect 11300 -2974 11474 -2958
rect 1909 -3453 1969 -3419
rect 6381 -3453 6441 -3419
rect 1909 -3479 1943 -3453
rect 6407 -3479 6441 -3453
rect 3872 -7142 4600 -7134
rect 2500 -7152 3228 -7142
rect 2500 -7216 2512 -7152
rect 3872 -7208 3888 -7142
rect 4588 -7208 4600 -7142
rect 2406 -7266 2526 -7254
rect 2406 -8042 2420 -7266
rect 2512 -8042 2526 -7266
rect 2406 -8054 2526 -8042
rect 2564 -7266 2684 -7254
rect 2564 -8042 2578 -7266
rect 2670 -8042 2684 -7266
rect 2564 -8054 2684 -8042
rect 2722 -7266 2842 -7254
rect 2722 -8042 2736 -7266
rect 2828 -8042 2842 -7266
rect 2722 -8054 2842 -8042
rect 2880 -7266 3000 -7254
rect 2880 -8042 2894 -7266
rect 2986 -8042 3000 -7266
rect 2880 -8054 3000 -8042
rect 3036 -7266 3156 -7254
rect 3036 -8042 3050 -7266
rect 3142 -8042 3156 -7266
rect 3036 -8054 3156 -8042
rect 3196 -7266 3316 -7254
rect 3196 -8042 3210 -7266
rect 3302 -8042 3316 -7266
rect 3196 -8054 3316 -8042
rect 3782 -7266 3902 -7254
rect 3782 -8044 3796 -7266
rect 3888 -8044 3902 -7266
rect 3782 -8054 3902 -8044
rect 3940 -7266 4060 -7254
rect 3940 -8044 3954 -7266
rect 4046 -8044 4060 -7266
rect 3940 -8054 4060 -8044
rect 4098 -7266 4218 -7254
rect 4098 -8044 4112 -7266
rect 4204 -8044 4218 -7266
rect 4098 -8054 4218 -8044
rect 4256 -7266 4376 -7254
rect 4256 -8044 4270 -7266
rect 4362 -8044 4376 -7266
rect 4256 -8054 4376 -8044
rect 4414 -7266 4534 -7254
rect 4414 -8044 4428 -7266
rect 4520 -8044 4534 -7266
rect 4414 -8054 4534 -8044
rect 4572 -7266 4692 -7254
rect 4572 -8044 4586 -7266
rect 4678 -8044 4692 -7266
rect 4572 -8054 4692 -8044
rect 2500 -8158 2512 -8092
rect 3212 -8158 3228 -8092
rect 2500 -8166 3228 -8158
rect 3872 -8168 3888 -8102
rect 4588 -8168 4600 -8102
rect 3872 -8176 4600 -8168
rect 1909 -8989 1943 -8963
rect 6407 -8989 6441 -8963
rect 1909 -9023 1969 -8989
rect 6381 -9023 6441 -8989
rect 8757 -4231 8817 -4197
rect 25211 -4231 25271 -4197
rect 8757 -4257 8791 -4231
rect 25237 -4257 25271 -4231
rect 16946 -4382 17342 -4372
rect 16946 -4556 16958 -4382
rect 17330 -4556 17342 -4382
rect 16946 -4566 17342 -4556
rect 16260 -4700 18034 -4640
rect 16648 -4744 16924 -4700
rect 10486 -4970 11230 -4958
rect 10486 -5346 10612 -4970
rect 11224 -5346 11230 -4970
rect 10486 -5358 11230 -5346
rect 12104 -4970 12504 -4958
rect 12104 -5346 12122 -4970
rect 12488 -5346 12504 -4970
rect 12104 -5358 12504 -5346
rect 12918 -4970 13178 -4958
rect 12918 -5346 12924 -4970
rect 13168 -5346 13178 -4970
rect 12918 -5358 13178 -5346
rect 13260 -4970 13660 -4958
rect 13260 -5346 13276 -4970
rect 13642 -5346 13660 -4970
rect 13260 -5358 13660 -5346
rect 14532 -4970 15276 -4958
rect 14532 -5346 14538 -4970
rect 15150 -5346 15276 -4970
rect 14532 -5358 15276 -5346
rect 9612 -5572 10060 -5450
rect 16648 -5530 16666 -4744
rect 16878 -5530 16924 -4744
rect 16648 -5576 16924 -5530
rect 17026 -4750 17266 -4734
rect 17026 -5526 17044 -4750
rect 17246 -5526 17266 -4750
rect 17026 -5542 17266 -5526
rect 17500 -4750 17712 -4734
rect 17500 -5526 17520 -4750
rect 17692 -5526 17712 -4750
rect 17500 -5542 17712 -5526
rect 16260 -5636 18034 -5576
rect 18788 -5808 18912 -5360
rect 21254 -5508 21400 -5402
rect 23260 -5414 23758 -5288
rect 10682 -5908 15086 -5888
rect 10682 -5948 12924 -5908
rect 11088 -5988 11248 -5984
rect 10522 -6000 11248 -5988
rect 10522 -6378 11092 -6000
rect 11242 -6378 11248 -6000
rect 10522 -6388 11248 -6378
rect 11088 -6394 11248 -6388
rect 11294 -6430 11612 -5948
rect 11660 -6000 11820 -5984
rect 11660 -6378 11666 -6000
rect 11814 -6378 11820 -6000
rect 11660 -6394 11820 -6378
rect 11866 -6430 12184 -5948
rect 12234 -6000 12850 -5984
rect 12234 -6378 12238 -6000
rect 12388 -6378 12850 -6000
rect 12234 -6394 12850 -6378
rect 12916 -6430 12924 -5948
rect 10682 -6470 12924 -6430
rect 13318 -5948 15086 -5908
rect 13318 -6430 13330 -5948
rect 13376 -6000 13536 -5984
rect 13376 -6378 13382 -6000
rect 13530 -6378 13536 -6000
rect 13376 -6394 13536 -6378
rect 13584 -6430 13900 -5948
rect 13948 -6000 14108 -5984
rect 13948 -6378 13954 -6000
rect 14102 -6378 14108 -6000
rect 13948 -6394 14108 -6378
rect 14156 -6430 14472 -5948
rect 16156 -5960 17118 -5950
rect 14520 -5988 14680 -5984
rect 14520 -6000 15248 -5988
rect 14520 -6378 14526 -6000
rect 14674 -6378 15248 -6000
rect 16156 -6050 16162 -5960
rect 16608 -6050 17118 -5960
rect 17176 -5960 18138 -5950
rect 17176 -6050 17686 -5960
rect 18132 -6050 18138 -5960
rect 14520 -6388 15248 -6378
rect 16600 -6108 16770 -6092
rect 14520 -6394 14680 -6388
rect 13318 -6470 15086 -6430
rect 10682 -6476 15086 -6470
rect 11088 -6518 11248 -6512
rect 10522 -6528 11248 -6518
rect 10522 -6906 11092 -6528
rect 11242 -6906 11248 -6528
rect 10522 -6918 11248 -6906
rect 11088 -6922 11248 -6918
rect 11294 -6958 11612 -6476
rect 11660 -6528 11820 -6512
rect 11660 -6906 11666 -6528
rect 11814 -6906 11820 -6528
rect 11660 -6922 11820 -6906
rect 11866 -6958 12184 -6476
rect 12234 -6528 12394 -6512
rect 12234 -6906 12238 -6528
rect 12388 -6906 12394 -6528
rect 12234 -6922 12394 -6906
rect 12440 -6958 12756 -6476
rect 12804 -6528 12964 -6512
rect 12804 -6906 12810 -6528
rect 12958 -6906 12964 -6528
rect 12804 -6922 12964 -6906
rect 13012 -6958 13328 -6476
rect 13376 -6528 13536 -6512
rect 13376 -6906 13382 -6528
rect 13530 -6906 13536 -6528
rect 13376 -6922 13536 -6906
rect 13584 -6958 13900 -6476
rect 13948 -6528 14108 -6512
rect 13948 -6906 13954 -6528
rect 14102 -6906 14108 -6528
rect 13948 -6922 14108 -6906
rect 14156 -6958 14472 -6476
rect 14522 -6518 14682 -6512
rect 14522 -6528 15248 -6518
rect 14522 -6906 14526 -6528
rect 14674 -6906 15248 -6528
rect 16600 -6886 16612 -6108
rect 16758 -6886 16770 -6108
rect 16600 -6902 16770 -6886
rect 16998 -6106 17298 -6092
rect 16998 -6890 17014 -6106
rect 17280 -6890 17298 -6106
rect 16998 -6902 17298 -6890
rect 17520 -6108 17690 -6092
rect 17520 -6886 17532 -6108
rect 17678 -6886 17690 -6108
rect 18768 -6830 18892 -6364
rect 21254 -6742 21400 -6636
rect 22948 -6810 24114 -6686
rect 17520 -6902 17690 -6886
rect 14522 -6918 15248 -6906
rect 14522 -6922 14682 -6918
rect 10682 -7018 15086 -6958
rect 16156 -7034 16162 -6944
rect 16608 -7034 17118 -6944
rect 16156 -7044 17118 -7034
rect 17176 -7034 17686 -6944
rect 18132 -7034 18138 -6944
rect 17176 -7044 18138 -7034
rect 10618 -7674 11048 -7438
rect 10620 -8006 11050 -7770
rect 24220 -7840 24650 -7604
rect 10620 -8338 11050 -8102
rect 24220 -8172 24650 -7936
rect 10620 -8670 11050 -8434
rect 24220 -8502 24650 -8266
rect 10620 -9002 11050 -8766
rect 24220 -8834 24650 -8598
rect 10620 -9334 11050 -9098
rect 24220 -9166 24650 -8930
rect 9614 -9488 10062 -9366
rect 10620 -9664 11050 -9428
rect 24220 -9500 24650 -9264
rect 24220 -9832 24650 -9596
rect 8757 -10301 8791 -10275
rect 25237 -10301 25271 -10275
rect 8757 -10335 8817 -10301
rect 25211 -10335 25271 -10301
rect 1683 -11629 1743 -11595
rect 25453 -11629 25513 -11595
rect 1683 -11655 1717 -11629
rect 25479 -11655 25513 -11629
rect 7146 -12454 7314 -12246
rect 8090 -12304 8232 -12102
rect 8086 -12400 8256 -12304
rect 8090 -12602 8232 -12400
rect 3134 -12982 3568 -12810
rect 3134 -13314 3566 -13098
rect 17762 -13154 19094 -12794
rect 19790 -13190 21916 -12568
rect 18532 -13242 18968 -13228
rect 18532 -13338 18544 -13242
rect 18954 -13338 18968 -13242
rect 18532 -13350 18968 -13338
rect 19994 -13242 21712 -13228
rect 19994 -13244 20918 -13242
rect 19994 -13352 20008 -13244
rect 20788 -13286 20918 -13244
rect 20788 -13352 20802 -13286
rect 19994 -13368 20802 -13352
rect 20904 -13350 20918 -13286
rect 21698 -13350 21712 -13242
rect 20904 -13368 21712 -13350
rect 3132 -13602 3566 -13430
rect 18532 -13600 18966 -13428
rect 19924 -13452 21780 -13426
rect 19924 -13600 19998 -13452
rect 20798 -13600 20908 -13452
rect 21708 -13600 21780 -13452
rect 19924 -13626 21780 -13600
rect 22452 -13486 22554 -12794
rect 22596 -13138 23404 -12574
rect 22596 -13344 22612 -13138
rect 23390 -13344 23404 -13138
rect 22596 -13362 23404 -13344
rect 23448 -13486 23482 -12794
rect 23524 -13136 24332 -12574
rect 23524 -13342 23540 -13136
rect 24318 -13342 24332 -13136
rect 23524 -13362 24332 -13342
rect 24376 -13486 24478 -12794
rect 22452 -13586 24478 -13486
rect 19994 -13702 20802 -13680
rect 2134 -13922 2562 -13746
rect 18932 -13920 19360 -13744
rect 19994 -13802 20010 -13702
rect 20786 -13760 20802 -13702
rect 20904 -13700 21712 -13680
rect 20904 -13760 20920 -13700
rect 20786 -13800 20920 -13760
rect 21696 -13800 21712 -13700
rect 20786 -13802 21712 -13800
rect 19994 -13820 21712 -13802
rect 21816 -13758 21956 -13746
rect 19994 -13896 20802 -13820
rect 20200 -13952 20600 -13896
rect 18932 -13994 19366 -13978
rect 2132 -14254 2564 -14038
rect 18932 -14132 18946 -13994
rect 19348 -14132 19366 -13994
rect 18932 -14146 19366 -14132
rect 2134 -14584 2566 -14368
rect 18932 -14418 19364 -14202
rect 20200 -14262 20242 -13952
rect 20556 -14262 20600 -13952
rect 20904 -13952 20920 -13856
rect 21696 -13952 21712 -13856
rect 21816 -13874 21828 -13758
rect 21944 -13874 21956 -13758
rect 21816 -13886 21956 -13874
rect 20904 -13966 21712 -13952
rect 20200 -14308 20600 -14262
rect 20854 -14052 21764 -14008
rect 20854 -14266 20916 -14052
rect 21698 -14266 21764 -14052
rect 19994 -14384 20802 -14308
rect 20854 -14330 21764 -14266
rect 22452 -14056 22554 -13586
rect 22596 -13718 23404 -13702
rect 22596 -13924 22612 -13718
rect 23390 -13924 23404 -13718
rect 22596 -13942 23404 -13924
rect 23448 -14056 23482 -13586
rect 23522 -13716 24330 -13702
rect 23522 -13922 23540 -13716
rect 24318 -13744 24330 -13716
rect 24318 -13898 24332 -13744
rect 24318 -13922 24330 -13898
rect 23522 -13942 24330 -13922
rect 24376 -14056 24478 -13586
rect 22452 -14156 24478 -14056
rect 19994 -14400 21712 -14384
rect 19994 -14500 20010 -14400
rect 20786 -14404 21712 -14400
rect 20786 -14444 20920 -14404
rect 20786 -14500 20802 -14444
rect 19994 -14524 20802 -14500
rect 20904 -14504 20920 -14444
rect 21696 -14504 21712 -14404
rect 20904 -14524 21712 -14504
rect 2132 -14916 2564 -14700
rect 18932 -14750 19364 -14534
rect 19926 -14600 21782 -14576
rect 19926 -14602 20908 -14600
rect 19926 -14750 19998 -14602
rect 20798 -14748 20908 -14602
rect 21708 -14748 21782 -14600
rect 20798 -14750 21782 -14748
rect 19926 -14776 21782 -14750
rect 22452 -14632 22554 -14156
rect 22596 -14298 23404 -14280
rect 22596 -14504 22612 -14298
rect 23390 -14504 23404 -14298
rect 22596 -14520 23404 -14504
rect 23448 -14632 23482 -14156
rect 23524 -14298 24332 -14280
rect 23524 -14504 23540 -14298
rect 24318 -14504 24332 -14298
rect 23524 -14520 24332 -14504
rect 24376 -14632 24478 -14156
rect 22452 -14732 24478 -14632
rect 19994 -14854 20802 -14838
rect 2132 -15248 2564 -15032
rect 18932 -15082 19364 -14866
rect 19994 -14962 20008 -14854
rect 20788 -14920 20802 -14854
rect 20904 -14854 21712 -14838
rect 20904 -14920 20920 -14854
rect 20788 -14962 20920 -14920
rect 21700 -14962 21712 -14854
rect 19994 -14978 21712 -14962
rect 2130 -15578 2562 -15362
rect 18932 -15414 19364 -15198
rect 2132 -15912 2564 -15696
rect 18932 -15746 19364 -15530
rect 19788 -15636 21914 -15014
rect 22452 -15590 22554 -14732
rect 22596 -14816 23404 -14802
rect 22596 -14966 22612 -14816
rect 23390 -14966 23404 -14816
rect 22596 -14982 23404 -14966
rect 22598 -15512 23404 -15020
rect 23448 -15590 23482 -14732
rect 22452 -15598 23482 -15590
rect 2132 -16242 2564 -16026
rect 18932 -16078 19364 -15862
rect 22452 -15872 22612 -15598
rect 23390 -15788 23482 -15598
rect 23524 -15100 24332 -14900
rect 23524 -15432 23630 -15100
rect 24228 -15432 24332 -15100
rect 23524 -15632 24332 -15432
rect 24376 -15788 24478 -14732
rect 23390 -15872 24478 -15788
rect 22452 -15888 24478 -15872
rect 19854 -16020 20254 -15994
rect 2132 -16576 2564 -16360
rect 18932 -16410 19364 -16194
rect 2130 -16908 2562 -16692
rect 18932 -16742 19364 -16526
rect 2130 -17240 2562 -17024
rect 18932 -17074 19364 -16858
rect 2132 -17570 2564 -17354
rect 18932 -17406 19364 -17190
rect 2132 -17904 2564 -17688
rect 18932 -17738 19364 -17522
rect 18930 -17816 19376 -17798
rect 18930 -17944 18944 -17816
rect 19354 -17944 19376 -17816
rect 18930 -17958 19376 -17944
rect 19854 -17992 19884 -16020
rect 20222 -17992 20254 -16020
rect 20462 -16008 21266 -15934
rect 20462 -16236 20474 -16008
rect 21252 -16236 21266 -16008
rect 22452 -16366 22554 -15888
rect 22596 -16032 23404 -16014
rect 22596 -16238 22612 -16032
rect 23390 -16238 23404 -16032
rect 22596 -16254 23404 -16238
rect 23448 -16366 23482 -15888
rect 23522 -16030 24330 -16014
rect 23522 -16236 23540 -16030
rect 24318 -16056 24330 -16030
rect 24318 -16210 24332 -16056
rect 24318 -16236 24330 -16210
rect 23522 -16254 24330 -16236
rect 24376 -16366 24478 -15888
rect 22452 -16466 24478 -16366
rect 22452 -16940 22554 -16466
rect 22596 -16606 23404 -16590
rect 22596 -16812 22612 -16606
rect 23390 -16812 23404 -16606
rect 22596 -16830 23404 -16812
rect 23448 -16940 23482 -16466
rect 23524 -16606 24332 -16590
rect 23524 -16812 23540 -16606
rect 24318 -16812 24332 -16606
rect 23524 -16830 24332 -16812
rect 24376 -16940 24478 -16466
rect 22452 -17040 24478 -16940
rect 22452 -17736 22554 -17040
rect 22596 -17186 23404 -17170
rect 22596 -17392 22612 -17186
rect 23390 -17392 23404 -17186
rect 2134 -18194 2562 -18018
rect 18932 -18192 19360 -18016
rect 19854 -18022 20254 -17992
rect 20462 -18010 20474 -17782
rect 21252 -18010 21266 -17782
rect 22596 -17958 23404 -17392
rect 23448 -17736 23482 -17040
rect 23524 -17186 24332 -17170
rect 23524 -17392 23540 -17186
rect 24318 -17392 24332 -17186
rect 23524 -17958 24332 -17392
rect 24376 -17736 24478 -17040
rect 20462 -18084 21266 -18010
rect 2130 -18518 2564 -18338
rect 24528 -18520 24962 -18340
rect 2130 -18850 2564 -18616
rect 2130 -19184 2564 -18950
rect 24530 -19016 24964 -18782
rect 2130 -19514 2564 -19280
rect 24530 -19348 24964 -19114
rect 2130 -19846 2564 -19612
rect 24530 -19680 24964 -19446
rect 2130 -20180 2564 -19946
rect 24530 -20012 24964 -19778
rect 2130 -20510 2564 -20276
rect 24530 -20344 24964 -20110
rect 2130 -20842 2564 -20608
rect 24530 -20676 24964 -20442
rect 2128 -21174 2562 -20940
rect 24530 -21008 24964 -20774
rect 2130 -21506 2564 -21272
rect 24528 -21342 24962 -21108
rect 2130 -21838 2564 -21604
rect 24530 -21672 24964 -21438
rect 2128 -22170 2562 -21936
rect 24528 -22004 24962 -21770
rect 24528 -22338 24962 -22104
rect 2130 -22624 2564 -22444
rect 24530 -22622 24964 -22442
rect 1683 -23613 1717 -23587
rect 25479 -23613 25513 -23587
rect 1683 -23647 1743 -23613
rect 25453 -23647 25513 -23613
<< viali >>
rect 3156 -1180 3236 -956
rect 5096 -1180 5176 -958
rect 11310 -2958 11468 -2180
rect 2512 -7216 3230 -7152
rect 3888 -7208 4588 -7142
rect 2420 -8042 2512 -7266
rect 2578 -8042 2670 -7266
rect 2736 -8042 2828 -7266
rect 2894 -8042 2986 -7266
rect 3050 -8042 3142 -7266
rect 3210 -8042 3302 -7266
rect 3796 -8044 3888 -7266
rect 3954 -8044 4046 -7266
rect 4112 -8044 4204 -7266
rect 4270 -8044 4362 -7266
rect 4428 -8044 4520 -7266
rect 4586 -8044 4678 -7266
rect 2512 -8158 3212 -8092
rect 3888 -8168 4588 -8102
rect 16958 -4556 17330 -4382
rect 10612 -5346 11224 -4970
rect 12122 -5346 12488 -4970
rect 12924 -5346 13168 -4970
rect 13276 -5346 13642 -4970
rect 14538 -5346 15150 -4970
rect 16666 -5530 16878 -4744
rect 17044 -5526 17246 -4750
rect 17520 -5526 17692 -4750
rect 11092 -6378 11242 -6000
rect 11666 -6378 11814 -6000
rect 12238 -6378 12388 -6000
rect 12924 -6470 13318 -5908
rect 13382 -6378 13530 -6000
rect 13954 -6378 14102 -6000
rect 14526 -6378 14674 -6000
rect 16162 -6050 16608 -5960
rect 17686 -6050 18132 -5960
rect 11092 -6906 11242 -6528
rect 11666 -6906 11814 -6528
rect 12238 -6906 12388 -6528
rect 12810 -6906 12958 -6528
rect 13382 -6906 13530 -6528
rect 13954 -6906 14102 -6528
rect 14526 -6906 14674 -6528
rect 16612 -6886 16758 -6108
rect 17014 -6890 17280 -6106
rect 17532 -6886 17678 -6108
rect 16162 -7034 16608 -6944
rect 17686 -7034 18132 -6944
rect 18544 -13338 18954 -13242
rect 20008 -13352 20788 -13244
rect 20918 -13350 21698 -13242
rect 19998 -13600 20798 -13452
rect 20908 -13600 21708 -13452
rect 22612 -13344 23390 -13138
rect 23540 -13342 24318 -13136
rect 20010 -13802 20786 -13702
rect 20920 -13800 21696 -13700
rect 18946 -14132 19348 -13994
rect 20242 -14262 20556 -13952
rect 20920 -13952 21696 -13856
rect 21828 -13874 21944 -13758
rect 20916 -14266 21698 -14052
rect 22612 -13924 23390 -13718
rect 23540 -13922 24318 -13716
rect 20010 -14500 20786 -14400
rect 20920 -14504 21696 -14404
rect 19998 -14750 20798 -14602
rect 20908 -14748 21708 -14600
rect 22612 -14504 23390 -14298
rect 23540 -14504 24318 -14298
rect 20008 -14962 20788 -14854
rect 20920 -14962 21700 -14854
rect 22612 -14966 23390 -14816
rect 22612 -15872 23390 -15598
rect 23630 -15432 24228 -15100
rect 18944 -17944 19354 -17816
rect 19884 -17992 20222 -16020
rect 20474 -16242 21252 -16008
rect 22612 -16238 23390 -16032
rect 23540 -16236 24318 -16030
rect 22612 -16812 23390 -16606
rect 23540 -16812 24318 -16606
rect 22612 -17392 23390 -17186
rect 20474 -18010 21252 -17776
rect 23540 -17392 24318 -17186
<< metal1 >>
rect 3592 -826 3992 -812
rect 3592 -946 3606 -826
rect 2882 -956 3606 -946
rect 1890 -1200 2090 -1000
rect 2242 -1202 2442 -1002
rect 2882 -1046 3156 -956
rect 3146 -1180 3156 -1046
rect 3236 -1046 3606 -956
rect 3236 -1180 3246 -1046
rect 3146 -1194 3246 -1180
rect 3592 -1200 3606 -1046
rect 3980 -1200 3992 -826
rect 3592 -1212 3992 -1200
rect 4338 -824 4738 -812
rect 4338 -1198 4350 -824
rect 4724 -948 4738 -824
rect 4724 -958 5454 -948
rect 4724 -1048 5096 -958
rect 4724 -1198 4738 -1048
rect 5086 -1180 5096 -1048
rect 5176 -1048 5454 -958
rect 5176 -1180 5186 -1048
rect 7066 -1128 7266 -928
rect 9798 -1130 9998 -930
rect 5086 -1192 5186 -1180
rect 11388 -1196 11588 -996
rect 23862 -1102 24062 -902
rect 4338 -1212 4738 -1198
rect 11300 -2180 11474 -2164
rect 11300 -2958 11310 -2180
rect 11468 -2958 11474 -2180
rect 11300 -2974 11474 -2958
rect 11504 -3012 11550 -2082
rect 11592 -2968 11980 -2170
rect 12600 -2224 13048 -2092
rect 11772 -2980 11980 -2968
rect 11480 -3198 11580 -3012
rect 11772 -3164 11780 -2980
rect 11972 -3164 11980 -2980
rect 11772 -3172 11980 -3164
rect 12772 -3176 12874 -3062
rect 11416 -3208 11616 -3198
rect 11416 -3386 11426 -3208
rect 11604 -3386 11616 -3208
rect 12772 -3294 13942 -3176
rect 11416 -3398 11616 -3386
rect 16946 -4382 17342 -4372
rect 16946 -4556 16958 -4382
rect 17330 -4556 17342 -4382
rect 16946 -4566 17342 -4556
rect 11772 -4626 11980 -4616
rect 11772 -4810 11780 -4626
rect 11972 -4810 11980 -4626
rect 16260 -4700 17076 -4640
rect 11772 -4816 11980 -4810
rect 16648 -4744 16924 -4700
rect 17106 -4734 17186 -4566
rect 17218 -4700 18034 -4640
rect 17266 -4706 17486 -4700
rect 10662 -4896 15100 -4816
rect 10466 -4970 11230 -4958
rect 10466 -5346 10478 -4970
rect 11224 -5346 11230 -4970
rect 10466 -5358 11230 -5346
rect 11436 -5420 12014 -4896
rect 12104 -4970 12504 -4958
rect 12104 -5346 12122 -4970
rect 12488 -5346 12504 -4970
rect 12104 -5358 12504 -5346
rect 12592 -5420 12844 -4896
rect 12918 -4970 13178 -4958
rect 12918 -5346 12924 -4970
rect 13168 -5346 13178 -4970
rect 12918 -5358 13178 -5346
rect 13260 -4970 13660 -4958
rect 13260 -5346 13276 -4970
rect 13642 -5346 13660 -4970
rect 13260 -5358 13660 -5346
rect 13748 -5420 14326 -4896
rect 16648 -4912 16666 -4744
rect 14532 -4970 15296 -4958
rect 14532 -5346 14538 -4970
rect 15284 -5346 15296 -4970
rect 16248 -5212 16666 -4912
rect 14532 -5358 15296 -5346
rect 9612 -5582 10060 -5452
rect 10662 -5500 15100 -5420
rect 16648 -5530 16666 -5212
rect 16878 -5530 16924 -4744
rect 16648 -5576 16924 -5530
rect 17026 -4750 17266 -4734
rect 17026 -5526 17044 -4750
rect 17246 -5526 17266 -4750
rect 17026 -5542 17266 -5526
rect 17328 -5570 17424 -4706
rect 17500 -4750 17712 -4734
rect 17500 -5526 17520 -4750
rect 17692 -4932 17712 -4750
rect 17692 -5232 18044 -4932
rect 17692 -5526 17712 -5232
rect 20942 -5250 21570 -5150
rect 17500 -5538 17712 -5526
rect 17266 -5576 17486 -5570
rect 16648 -5636 17534 -5576
rect 3364 -7142 3370 -6962
rect 2500 -7152 3370 -7142
rect 2500 -7216 2512 -7152
rect 3230 -7216 3370 -7152
rect 2500 -7222 3370 -7216
rect 3478 -7222 3484 -6962
rect 3614 -7214 3620 -6954
rect 3728 -7134 3734 -6954
rect 3728 -7142 4600 -7134
rect 3728 -7208 3888 -7142
rect 4588 -7208 4600 -7142
rect 3728 -7214 4600 -7208
rect 2406 -8054 2412 -7254
rect 2520 -8054 2526 -7254
rect 2564 -8054 2570 -7254
rect 2678 -8054 2684 -7254
rect 2722 -8054 2728 -7254
rect 2836 -8054 2842 -7254
rect 2880 -8054 2886 -7254
rect 2994 -8054 3000 -7254
rect 3036 -8054 3042 -7254
rect 3150 -8054 3156 -7254
rect 3196 -8054 3202 -7254
rect 3310 -8054 3316 -7254
rect 3364 -8086 3370 -7906
rect 2500 -8092 3370 -8086
rect 2500 -8158 2512 -8092
rect 3212 -8158 3370 -8092
rect 2500 -8166 3370 -8158
rect 3478 -8086 3484 -7906
rect 3478 -8166 3486 -8086
rect 3614 -8176 3620 -7916
rect 3728 -8096 3734 -7916
rect 3782 -8054 3790 -7254
rect 3894 -8054 3902 -7254
rect 3940 -8054 3946 -7254
rect 4054 -8054 4060 -7254
rect 4098 -8054 4104 -7254
rect 4212 -8054 4218 -7254
rect 4256 -8054 4262 -7254
rect 4370 -8054 4376 -7254
rect 4414 -8054 4420 -7254
rect 4528 -8054 4534 -7254
rect 4572 -8054 4578 -7254
rect 4686 -8054 4692 -7254
rect 9732 -7411 9948 -5678
rect 10682 -5906 15086 -5888
rect 10682 -5948 12924 -5906
rect 10522 -6000 11248 -5988
rect 10522 -6378 11092 -6000
rect 11242 -6378 11248 -6000
rect 10522 -6388 11248 -6378
rect 11088 -6518 11248 -6388
rect 10522 -6528 11248 -6518
rect 10522 -6906 11092 -6528
rect 11242 -6906 11248 -6528
rect 10522 -6918 11248 -6906
rect 11088 -7056 11248 -6918
rect 11294 -6958 11612 -5948
rect 11660 -5990 11820 -5984
rect 11660 -6388 11666 -5990
rect 11814 -6388 11820 -5990
rect 11660 -6518 11820 -6388
rect 11660 -6916 11666 -6518
rect 11814 -6916 11820 -6518
rect 11660 -6922 11820 -6916
rect 11866 -6958 12184 -5948
rect 11294 -7018 12184 -6958
rect 12234 -5988 12392 -5984
rect 12234 -6000 12850 -5988
rect 12234 -6378 12238 -6000
rect 12388 -6378 12850 -6000
rect 12234 -6394 12850 -6378
rect 12234 -6528 12394 -6394
rect 12234 -6906 12238 -6528
rect 12388 -6906 12394 -6528
rect 12234 -7056 12394 -6906
rect 12440 -6958 12756 -6430
rect 12912 -6470 12924 -5948
rect 13318 -5948 15086 -5906
rect 13318 -6470 13330 -5948
rect 12912 -6482 13330 -6470
rect 13376 -6000 13536 -5984
rect 13376 -6378 13382 -6000
rect 13530 -6378 13536 -6000
rect 12804 -6518 12964 -6512
rect 12804 -6916 12810 -6518
rect 12958 -6916 12964 -6518
rect 12804 -6922 12964 -6916
rect 13012 -6958 13328 -6482
rect 13376 -6528 13536 -6378
rect 13376 -6906 13382 -6528
rect 13530 -6906 13536 -6528
rect 12440 -7018 13330 -6958
rect 13376 -7056 13536 -6906
rect 13584 -6958 13900 -5948
rect 13948 -5990 14108 -5984
rect 13948 -6388 13954 -5990
rect 14102 -6388 14108 -5990
rect 13948 -6518 14108 -6388
rect 13948 -6916 13954 -6518
rect 14102 -6916 14108 -6518
rect 13948 -6922 14108 -6916
rect 14156 -6958 14472 -5948
rect 16036 -5960 16620 -5950
rect 14520 -6000 15248 -5988
rect 14520 -6378 14526 -6000
rect 14674 -6378 15248 -6000
rect 14520 -6388 15248 -6378
rect 16036 -6050 16162 -5960
rect 16608 -6050 16620 -5960
rect 16036 -6056 16602 -6050
rect 14520 -6518 14680 -6388
rect 14520 -6528 15248 -6518
rect 14520 -6906 14526 -6528
rect 14674 -6906 15248 -6528
rect 14520 -6918 15248 -6906
rect 16036 -6554 16156 -6056
rect 16648 -6092 16728 -5636
rect 16768 -6056 16954 -6048
rect 16600 -6108 16770 -6092
rect 16600 -6392 16612 -6108
rect 13584 -7018 14474 -6958
rect 14520 -7056 14680 -6918
rect 16036 -7036 16044 -6554
rect 16148 -6938 16156 -6554
rect 16248 -6692 16612 -6392
rect 16600 -6886 16612 -6692
rect 16758 -6886 16770 -6108
rect 16600 -6902 16770 -6886
rect 16830 -6938 16954 -6056
rect 17340 -6056 17526 -6050
rect 16998 -6106 17298 -6092
rect 16998 -6890 17014 -6106
rect 17280 -6890 17298 -6106
rect 16998 -6902 17298 -6890
rect 17340 -6938 17464 -6056
rect 17564 -6092 17644 -5538
rect 18788 -5808 18920 -5360
rect 19616 -5452 19796 -5446
rect 17674 -5960 18258 -5950
rect 17674 -6050 17686 -5960
rect 18132 -6050 18258 -5960
rect 17780 -6056 18258 -6050
rect 17520 -6108 17690 -6092
rect 17520 -6886 17532 -6108
rect 17678 -6382 17690 -6108
rect 17678 -6682 18044 -6382
rect 18138 -6554 18258 -6056
rect 17678 -6886 17690 -6682
rect 17520 -6902 17690 -6886
rect 18138 -6938 18146 -6554
rect 16148 -6944 17118 -6938
rect 16148 -7034 16162 -6944
rect 16608 -7034 17118 -6944
rect 16148 -7036 17118 -7034
rect 16036 -7044 17118 -7036
rect 16160 -7046 17118 -7044
rect 17176 -6944 18146 -6938
rect 17176 -7034 17686 -6944
rect 18132 -7034 18146 -6944
rect 17176 -7036 18146 -7034
rect 18250 -7036 18258 -6554
rect 18768 -6830 18898 -6364
rect 19432 -6734 19978 -5452
rect 20574 -6030 20674 -5530
rect 20942 -6030 21042 -5250
rect 20574 -6130 21042 -6030
rect 20574 -6654 20674 -6130
rect 17176 -7046 18258 -7036
rect 11088 -7256 14680 -7056
rect 19616 -7380 19796 -6734
rect 20942 -6864 21042 -6130
rect 21290 -6010 21390 -5610
rect 21470 -5792 21570 -5250
rect 21620 -5274 21820 -5074
rect 21620 -5716 21662 -5274
rect 21718 -6010 21818 -5328
rect 21290 -6110 21818 -6010
rect 21290 -6516 21390 -6110
rect 21454 -6864 21554 -6326
rect 20940 -6964 21554 -6864
rect 21620 -6878 21662 -6412
rect 21718 -6828 21818 -6110
rect 21900 -5990 22000 -5406
rect 23260 -5424 23758 -5288
rect 22914 -5594 23666 -5494
rect 22914 -5842 23014 -5594
rect 22714 -5852 23014 -5842
rect 21900 -5996 22308 -5990
rect 21900 -6124 22006 -5996
rect 22302 -6124 22308 -5996
rect 21900 -6130 22308 -6124
rect 21900 -6738 22000 -6130
rect 22714 -6132 22726 -5852
rect 23002 -6132 23014 -5852
rect 22714 -6142 23014 -6132
rect 23434 -5930 23584 -5654
rect 24010 -5930 24210 -5924
rect 23434 -6130 24010 -5930
rect 22714 -6496 22814 -6142
rect 23434 -6438 23584 -6130
rect 24010 -6136 24210 -6130
rect 22714 -6596 24016 -6496
rect 22948 -6810 24114 -6676
rect 21620 -7078 21820 -6878
rect 9732 -7533 10357 -7411
rect 3728 -8102 4600 -8096
rect 3728 -8168 3888 -8102
rect 4588 -8168 4600 -8102
rect 3728 -8176 4600 -8168
rect 9732 -9268 9948 -7533
rect 9614 -9488 10062 -9356
rect 10235 -9748 10357 -7533
rect 10618 -7674 11048 -7438
rect 19616 -7560 24652 -7380
rect 10620 -8006 11050 -7770
rect 24220 -7840 24650 -7604
rect 10620 -8338 11050 -8102
rect 24220 -8172 24650 -7936
rect 10620 -8670 11050 -8434
rect 24220 -8502 24650 -8266
rect 10620 -9002 11050 -8766
rect 24220 -8834 24650 -8598
rect 10620 -9334 11050 -9098
rect 24220 -9166 24650 -8930
rect 10620 -9664 11050 -9428
rect 24220 -9500 24650 -9264
rect 10234 -9870 11052 -9748
rect 24220 -9832 24650 -9596
rect 7370 -12501 7478 -12200
rect 7534 -12270 7714 -12260
rect 7534 -12430 7542 -12270
rect 7704 -12430 7714 -12270
rect 7534 -12440 7714 -12430
rect 8336 -12264 9798 -12262
rect 8336 -12442 9886 -12264
rect 9978 -12268 11464 -12252
rect 9978 -12434 9998 -12268
rect 11440 -12434 11464 -12268
rect 9978 -12452 11464 -12434
rect 11640 -12268 13126 -12252
rect 11640 -12434 11662 -12268
rect 13104 -12434 13126 -12268
rect 20278 -12298 20478 -12284
rect 20278 -12302 20292 -12298
rect 13236 -12306 20292 -12302
rect 13190 -12398 20292 -12306
rect 13236 -12402 20292 -12398
rect 11640 -12452 13126 -12434
rect 20278 -12468 20292 -12402
rect 20464 -12468 20478 -12298
rect 20278 -12484 20478 -12468
rect 7339 -12620 7514 -12501
rect 7339 -12910 7346 -12620
rect 7506 -12910 7514 -12620
rect 7339 -12916 7514 -12910
rect 22452 -13070 24376 -12794
rect 3134 -13314 3566 -13098
rect 18532 -13242 21712 -13228
rect 18532 -13338 18544 -13242
rect 18954 -13244 20918 -13242
rect 18954 -13322 20008 -13244
rect 18954 -13338 19822 -13322
rect 18532 -13350 19822 -13338
rect 19460 -13368 19822 -13350
rect 19994 -13352 20008 -13322
rect 20788 -13330 20918 -13244
rect 20788 -13352 20802 -13330
rect 19994 -13368 20802 -13352
rect 20904 -13350 20918 -13330
rect 21698 -13350 21712 -13242
rect 20904 -13368 21712 -13350
rect 16048 -13986 19366 -13978
rect 2132 -14254 2564 -14038
rect 16048 -14136 16062 -13986
rect 16542 -13994 19366 -13986
rect 16542 -14132 18946 -13994
rect 19348 -14132 19366 -13994
rect 16542 -14136 19366 -14132
rect 16048 -14146 19366 -14136
rect 2134 -14584 2566 -14368
rect 18932 -14418 19364 -14202
rect 2132 -14916 2564 -14700
rect 18932 -14750 19364 -14534
rect 19460 -14838 19640 -13368
rect 19698 -13440 21780 -13426
rect 19698 -14762 19712 -13440
rect 19844 -13452 21780 -13440
rect 19844 -13600 19998 -13452
rect 20798 -13600 20908 -13452
rect 21708 -13600 21780 -13452
rect 19844 -13626 21780 -13600
rect 22452 -13450 22554 -13070
rect 22596 -13138 23404 -13122
rect 22596 -13344 22612 -13138
rect 23390 -13160 23404 -13138
rect 23524 -13136 24332 -13122
rect 23524 -13160 23540 -13136
rect 23390 -13326 23540 -13160
rect 23390 -13344 23404 -13326
rect 22596 -13362 23404 -13344
rect 23524 -13342 23540 -13326
rect 24318 -13160 24332 -13136
rect 24318 -13326 25176 -13160
rect 24318 -13342 24332 -13326
rect 23524 -13362 24332 -13342
rect 24376 -13450 24478 -13374
rect 22452 -13618 24478 -13450
rect 19844 -14576 19858 -13626
rect 19994 -13702 20802 -13680
rect 19994 -13802 20010 -13702
rect 20786 -13718 20802 -13702
rect 20904 -13700 21712 -13680
rect 20904 -13718 20920 -13700
rect 20786 -13800 20920 -13718
rect 21696 -13800 21712 -13700
rect 21816 -13758 21956 -13746
rect 20786 -13802 21712 -13800
rect 19994 -13820 21712 -13802
rect 19994 -13896 20802 -13820
rect 21748 -13848 21828 -13758
rect 20908 -13856 21828 -13848
rect 20200 -13906 20600 -13896
rect 20200 -14296 20214 -13906
rect 20590 -14296 20600 -13906
rect 20908 -13952 20920 -13856
rect 21696 -13874 21828 -13856
rect 21944 -13874 21956 -13758
rect 21696 -13908 21956 -13874
rect 21696 -13952 21708 -13908
rect 20908 -13964 21708 -13952
rect 20200 -14308 20600 -14296
rect 20854 -14030 21764 -14008
rect 20854 -14306 20882 -14030
rect 21736 -14170 21764 -14030
rect 22452 -14022 22554 -13618
rect 22596 -13716 23404 -13702
rect 22596 -13924 22612 -13716
rect 23390 -13738 23404 -13716
rect 23522 -13714 24330 -13702
rect 23522 -13738 23540 -13714
rect 23390 -13904 23540 -13738
rect 23390 -13924 23404 -13904
rect 22596 -13942 23404 -13924
rect 23522 -13922 23540 -13904
rect 24318 -13922 24330 -13714
rect 23522 -13942 24330 -13922
rect 24376 -14022 24478 -13618
rect 21736 -14306 22400 -14170
rect 19994 -14384 20802 -14308
rect 20854 -14330 22400 -14306
rect 19994 -14400 22156 -14384
rect 19994 -14500 20010 -14400
rect 20786 -14404 22156 -14400
rect 20786 -14486 20920 -14404
rect 20786 -14500 20802 -14486
rect 19994 -14524 20802 -14500
rect 20904 -14504 20920 -14486
rect 21696 -14482 22156 -14404
rect 21696 -14504 21712 -14482
rect 20904 -14524 21712 -14504
rect 19844 -14600 21782 -14576
rect 19844 -14602 20908 -14600
rect 19844 -14750 19998 -14602
rect 20798 -14748 20908 -14602
rect 21708 -14748 21782 -14600
rect 20798 -14750 21782 -14748
rect 19844 -14762 21782 -14750
rect 19698 -14776 21782 -14762
rect 2132 -15248 2564 -15032
rect 18932 -15082 19364 -14866
rect 19460 -14884 19822 -14838
rect 19994 -14854 20802 -14838
rect 19994 -14884 20008 -14854
rect 19460 -14962 20008 -14884
rect 20788 -14876 20802 -14854
rect 20904 -14854 21712 -14838
rect 20904 -14876 20920 -14854
rect 20788 -14962 20920 -14876
rect 21700 -14962 21712 -14854
rect 19460 -14978 21712 -14962
rect 18402 -15164 18802 -15148
rect 2130 -15578 2562 -15362
rect 18402 -15530 18420 -15164
rect 18784 -15530 18802 -15164
rect 18932 -15414 19364 -15198
rect 18402 -15548 18802 -15530
rect 2132 -15912 2564 -15696
rect 2132 -16242 2564 -16026
rect 2132 -16576 2564 -16360
rect 2130 -16908 2562 -16692
rect 2130 -17240 2562 -17024
rect 2132 -17570 2564 -17354
rect 2132 -17904 2564 -17688
rect 18560 -17798 18660 -15548
rect 18932 -15746 19364 -15530
rect 21956 -15590 22156 -14482
rect 22240 -14884 22400 -14330
rect 22452 -14190 24478 -14022
rect 22452 -14598 22554 -14190
rect 24376 -14268 24478 -14190
rect 22596 -14298 23404 -14280
rect 22596 -14504 22612 -14298
rect 23390 -14316 23404 -14298
rect 23524 -14298 24332 -14280
rect 23524 -14316 23540 -14298
rect 23390 -14482 23540 -14316
rect 23390 -14504 23404 -14482
rect 22596 -14520 23404 -14504
rect 23524 -14504 23540 -14482
rect 24318 -14316 24332 -14298
rect 24576 -14316 25176 -13326
rect 24318 -14482 25176 -14316
rect 24318 -14504 24332 -14482
rect 23524 -14520 24332 -14504
rect 24376 -14598 24478 -14532
rect 22452 -14766 24478 -14598
rect 22452 -14834 22554 -14766
rect 22596 -14816 23404 -14802
rect 22596 -14884 22612 -14816
rect 22240 -14966 22612 -14884
rect 23390 -14966 23404 -14816
rect 22240 -14982 23404 -14966
rect 23600 -14938 24258 -14900
rect 22452 -15184 22554 -15040
rect 22452 -15352 23448 -15184
rect 22452 -15590 22554 -15352
rect 21956 -15598 23486 -15590
rect 21956 -15750 22612 -15598
rect 18932 -16078 19364 -15862
rect 22452 -15872 22612 -15750
rect 23390 -15752 23486 -15598
rect 23600 -15592 23628 -14938
rect 24228 -15592 24258 -14938
rect 23600 -15634 24258 -15592
rect 24376 -15752 24478 -14766
rect 23390 -15872 24478 -15752
rect 22452 -15920 24478 -15872
rect 22452 -15946 23486 -15920
rect 19854 -16020 20254 -15994
rect 18932 -16410 19364 -16194
rect 18932 -16742 19364 -16526
rect 18932 -17074 19364 -16858
rect 18932 -17406 19364 -17190
rect 18932 -17738 19364 -17522
rect 18560 -17816 19376 -17798
rect 18560 -17944 18944 -17816
rect 19354 -17944 19376 -17816
rect 18560 -17958 19376 -17944
rect 19854 -17992 19884 -16020
rect 20222 -17992 20254 -16020
rect 20464 -16008 21264 -15994
rect 19854 -18022 20254 -17992
rect 20332 -18116 20432 -16094
rect 20464 -16242 20474 -16008
rect 21252 -16242 21264 -16008
rect 20464 -16268 20476 -16242
rect 21250 -16268 21264 -16242
rect 20464 -16284 21264 -16268
rect 20464 -16324 21264 -16312
rect 20464 -16430 20474 -16324
rect 21252 -16430 21264 -16324
rect 20464 -16442 21264 -16430
rect 20464 -16482 21264 -16470
rect 20464 -16588 20474 -16482
rect 21252 -16588 21264 -16482
rect 20464 -16600 21264 -16588
rect 20464 -16640 21264 -16628
rect 20464 -16746 20474 -16640
rect 21252 -16746 21264 -16640
rect 20464 -16758 21264 -16746
rect 20464 -16798 21264 -16786
rect 20464 -16904 20474 -16798
rect 21252 -16904 21264 -16798
rect 20464 -16916 21264 -16904
rect 20464 -16956 21264 -16944
rect 20464 -17062 20474 -16956
rect 21252 -17062 21264 -16956
rect 20464 -17074 21264 -17062
rect 20464 -17114 21264 -17102
rect 20464 -17220 20476 -17114
rect 21254 -17220 21264 -17114
rect 20464 -17232 21264 -17220
rect 20464 -17272 21264 -17260
rect 20464 -17378 20474 -17272
rect 21252 -17378 21264 -17272
rect 20464 -17390 21264 -17378
rect 20464 -17430 21264 -17418
rect 20464 -17536 20474 -17430
rect 21252 -17536 21264 -17430
rect 20464 -17548 21264 -17536
rect 20464 -17588 21264 -17576
rect 20464 -17694 20474 -17588
rect 21252 -17694 21264 -17588
rect 20464 -17706 21264 -17694
rect 20464 -17750 21264 -17734
rect 20464 -17776 20476 -17750
rect 21250 -17776 21264 -17750
rect 20464 -18010 20474 -17776
rect 21252 -18010 21264 -17776
rect 20464 -18022 21264 -18010
rect 21296 -18116 21396 -16094
rect 22452 -16332 22554 -15946
rect 24376 -16000 24478 -15920
rect 22596 -16032 23404 -16014
rect 22596 -16238 22612 -16032
rect 23390 -16050 23404 -16032
rect 23522 -16030 24330 -16014
rect 23522 -16050 23540 -16030
rect 23390 -16216 23540 -16050
rect 23390 -16238 23404 -16216
rect 22596 -16254 23404 -16238
rect 23522 -16236 23540 -16216
rect 24318 -16050 24330 -16030
rect 24576 -16050 25176 -14482
rect 24318 -16216 25176 -16050
rect 24318 -16236 24330 -16216
rect 23522 -16254 24330 -16236
rect 24376 -16332 24478 -16264
rect 22452 -16500 24478 -16332
rect 21704 -16590 22104 -16576
rect 21704 -17098 21718 -16590
rect 22090 -17098 22104 -16590
rect 21704 -17112 22104 -17098
rect 22452 -16906 22554 -16500
rect 22596 -16604 23404 -16590
rect 22596 -16812 22610 -16604
rect 23388 -16606 23404 -16604
rect 23390 -16628 23404 -16606
rect 23524 -16604 24332 -16590
rect 23524 -16628 23540 -16604
rect 23390 -16794 23540 -16628
rect 23390 -16812 23404 -16794
rect 22596 -16830 23404 -16812
rect 23524 -16812 23540 -16794
rect 24318 -16812 24332 -16604
rect 23524 -16830 24332 -16812
rect 24376 -16906 24478 -16500
rect 22452 -17074 24478 -16906
rect 20332 -18216 21396 -18116
rect 2130 -18850 2564 -18616
rect 2130 -19184 2564 -18950
rect 2130 -19514 2564 -19280
rect 2130 -19846 2564 -19612
rect 2130 -20180 2564 -19946
rect 2130 -20510 2564 -20276
rect 20776 -20592 20936 -18216
rect 21830 -18388 21990 -17112
rect 22452 -17460 22554 -17074
rect 24376 -17158 24478 -17074
rect 22596 -17186 23404 -17170
rect 22596 -17392 22612 -17186
rect 23390 -17206 23404 -17186
rect 23524 -17186 24332 -17170
rect 23524 -17206 23540 -17186
rect 23390 -17372 23540 -17206
rect 23390 -17392 23404 -17372
rect 22596 -17410 23404 -17392
rect 23524 -17392 23540 -17372
rect 24318 -17206 24332 -17186
rect 24576 -17206 25176 -16216
rect 24318 -17372 25176 -17206
rect 24318 -17392 24332 -17372
rect 23524 -17410 24332 -17392
rect 22452 -17736 24376 -17460
rect 21830 -18548 23334 -18388
rect 23174 -18572 23334 -18548
rect 23174 -18732 24982 -18572
rect 23174 -19970 23334 -18732
rect 24530 -19016 24964 -18782
rect 24530 -19348 24964 -19114
rect 24530 -19680 24964 -19446
rect 23102 -19984 23402 -19970
rect 23102 -20260 23114 -19984
rect 23386 -20260 23402 -19984
rect 24530 -20012 24964 -19778
rect 23102 -20270 23402 -20260
rect 20704 -20606 21004 -20592
rect 2130 -20842 2564 -20608
rect 20704 -20882 20718 -20606
rect 20990 -20882 21004 -20606
rect 20704 -20892 21004 -20882
rect 2128 -21174 2562 -20940
rect 2130 -21506 2564 -21272
rect 2130 -21838 2564 -21604
rect 2128 -22170 2562 -21936
rect 20776 -22222 20936 -20892
rect 2136 -22382 20936 -22222
rect 20776 -22932 20936 -22382
rect 23174 -22932 23334 -20270
rect 24530 -20344 24964 -20110
rect 24530 -20676 24964 -20442
rect 24530 -21008 24964 -20774
rect 24528 -21342 24962 -21108
rect 24530 -21672 24964 -21438
rect 24528 -22004 24962 -21770
rect 24528 -22338 24962 -22104
rect 20458 -23032 21408 -22932
rect 22740 -23032 23658 -22932
rect 20776 -23304 20936 -23032
rect 23174 -23304 23334 -23032
rect 20656 -23312 21056 -23304
rect 20656 -23696 20664 -23312
rect 21048 -23696 21056 -23312
rect 20656 -23704 21056 -23696
rect 23054 -23316 23454 -23304
rect 23054 -23690 23070 -23316
rect 23440 -23690 23454 -23316
rect 23054 -23704 23454 -23690
<< via1 >>
rect 3606 -1200 3980 -826
rect 4350 -1198 4724 -824
rect 11780 -3164 11972 -2980
rect 11426 -3386 11604 -3208
rect 13942 -3470 14128 -3124
rect 14344 -3464 14520 -3152
rect 11780 -4810 11972 -4626
rect 10478 -5346 10612 -4970
rect 10612 -5346 11224 -4970
rect 12122 -5346 12488 -4970
rect 12924 -5346 13168 -4970
rect 13276 -5346 13642 -4970
rect 14538 -5346 15150 -4970
rect 15150 -5346 15284 -4970
rect 3370 -7222 3478 -6962
rect 3620 -7214 3728 -6954
rect 2412 -7266 2520 -7254
rect 2412 -8042 2420 -7266
rect 2420 -8042 2512 -7266
rect 2512 -8042 2520 -7266
rect 2412 -8054 2520 -8042
rect 2570 -7266 2678 -7254
rect 2570 -8042 2578 -7266
rect 2578 -8042 2670 -7266
rect 2670 -8042 2678 -7266
rect 2570 -8054 2678 -8042
rect 2728 -7266 2836 -7254
rect 2728 -8042 2736 -7266
rect 2736 -8042 2828 -7266
rect 2828 -8042 2836 -7266
rect 2728 -8054 2836 -8042
rect 2886 -7266 2994 -7254
rect 2886 -8042 2894 -7266
rect 2894 -8042 2986 -7266
rect 2986 -8042 2994 -7266
rect 2886 -8054 2994 -8042
rect 3042 -7266 3150 -7254
rect 3042 -8042 3050 -7266
rect 3050 -8042 3142 -7266
rect 3142 -8042 3150 -7266
rect 3042 -8054 3150 -8042
rect 3202 -7266 3310 -7254
rect 3202 -8042 3210 -7266
rect 3210 -8042 3302 -7266
rect 3302 -8042 3310 -7266
rect 3202 -8054 3310 -8042
rect 3370 -8166 3478 -7906
rect 3620 -8176 3728 -7916
rect 3790 -7266 3894 -7254
rect 3790 -8044 3796 -7266
rect 3796 -8044 3888 -7266
rect 3888 -8044 3894 -7266
rect 3790 -8054 3894 -8044
rect 3946 -7266 4054 -7254
rect 3946 -8044 3954 -7266
rect 3954 -8044 4046 -7266
rect 4046 -8044 4054 -7266
rect 3946 -8054 4054 -8044
rect 4104 -7266 4212 -7254
rect 4104 -8044 4112 -7266
rect 4112 -8044 4204 -7266
rect 4204 -8044 4212 -7266
rect 4104 -8054 4212 -8044
rect 4262 -7266 4370 -7254
rect 4262 -8044 4270 -7266
rect 4270 -8044 4362 -7266
rect 4362 -8044 4370 -7266
rect 4262 -8054 4370 -8044
rect 4420 -7266 4528 -7254
rect 4420 -8044 4428 -7266
rect 4428 -8044 4520 -7266
rect 4520 -8044 4528 -7266
rect 4420 -8054 4528 -8044
rect 4578 -7266 4686 -7254
rect 4578 -8044 4586 -7266
rect 4586 -8044 4678 -7266
rect 4678 -8044 4686 -7266
rect 4578 -8054 4686 -8044
rect 12924 -5908 13318 -5906
rect 11666 -6000 11814 -5990
rect 11666 -6378 11814 -6000
rect 11666 -6388 11814 -6378
rect 11666 -6528 11814 -6518
rect 11666 -6906 11814 -6528
rect 11666 -6916 11814 -6906
rect 12924 -6468 13318 -5908
rect 12810 -6528 12958 -6518
rect 12810 -6906 12958 -6528
rect 12810 -6916 12958 -6906
rect 13954 -6000 14102 -5990
rect 13954 -6378 14102 -6000
rect 13954 -6388 14102 -6378
rect 13954 -6528 14102 -6518
rect 13954 -6906 14102 -6528
rect 13954 -6916 14102 -6906
rect 16044 -7036 16148 -6554
rect 17014 -6890 17280 -6106
rect 18146 -7036 18250 -6554
rect 22006 -6124 22302 -5996
rect 22726 -6132 23002 -5852
rect 24010 -6130 24210 -5930
rect 7542 -12430 7704 -12270
rect 9998 -12434 11440 -12268
rect 11662 -12434 13104 -12268
rect 20292 -12468 20464 -12298
rect 7346 -12910 7506 -12620
rect 16062 -14136 16542 -13986
rect 18946 -14132 19348 -13994
rect 19712 -14762 19844 -13440
rect 20214 -13952 20590 -13906
rect 20214 -14262 20242 -13952
rect 20242 -14262 20556 -13952
rect 20556 -14262 20590 -13952
rect 20214 -14296 20590 -14262
rect 20882 -14052 21736 -14030
rect 20882 -14266 20916 -14052
rect 20916 -14266 21698 -14052
rect 21698 -14266 21736 -14052
rect 22612 -13718 23390 -13716
rect 22612 -13924 23390 -13718
rect 23540 -13716 24318 -13714
rect 23540 -13922 24318 -13716
rect 20882 -14306 21736 -14266
rect 18420 -15530 18784 -15164
rect 23628 -15100 24228 -14938
rect 23628 -15432 23630 -15100
rect 23630 -15432 24228 -15100
rect 23628 -15592 24228 -15432
rect 19884 -17992 20222 -16020
rect 20476 -16242 21250 -16010
rect 20476 -16268 21250 -16242
rect 20474 -16430 21252 -16324
rect 20474 -16588 21252 -16482
rect 20474 -16746 21252 -16640
rect 20474 -16904 21252 -16798
rect 20474 -17062 21252 -16956
rect 20476 -17220 21254 -17114
rect 20474 -17378 21252 -17272
rect 20474 -17536 21252 -17430
rect 20474 -17694 21252 -17588
rect 20476 -17776 21250 -17750
rect 20476 -18008 21250 -17776
rect 21718 -17098 22090 -16590
rect 22610 -16606 23388 -16604
rect 22610 -16812 22612 -16606
rect 22612 -16812 23388 -16606
rect 23540 -16606 24318 -16604
rect 23540 -16812 24318 -16606
rect 23114 -20260 23386 -19984
rect 20718 -20882 20990 -20606
rect 20664 -23696 21048 -23312
rect 23070 -23690 23440 -23316
<< metal2 >>
rect 3592 -826 3992 -812
rect 3592 -1200 3606 -826
rect 3980 -1200 3992 -826
rect 3592 -1212 3992 -1200
rect 4338 -824 4738 -812
rect 4338 -1198 4350 -824
rect 4724 -1198 4738 -824
rect 4338 -1212 4738 -1198
rect 11772 -2980 11980 -2972
rect 11772 -3164 11780 -2980
rect 11972 -3164 11980 -2980
rect 11772 -3172 11980 -3164
rect 13934 -3124 14136 -3116
rect 11416 -3208 11616 -3198
rect 11416 -3386 11426 -3208
rect 11604 -3386 11616 -3208
rect 11416 -3398 11616 -3386
rect 11466 -3808 11566 -3398
rect 7582 -3908 11566 -3808
rect 5526 -6710 5726 -6660
rect 7582 -6710 7682 -3908
rect 11826 -4616 11926 -3172
rect 13934 -3470 13942 -3124
rect 14128 -3470 14136 -3124
rect 13934 -3476 14136 -3470
rect 14332 -3152 14532 -3140
rect 14332 -3464 14344 -3152
rect 14520 -3464 14532 -3152
rect 14332 -3476 14532 -3464
rect 13962 -3882 14102 -3476
rect 14360 -3512 14500 -3476
rect 14360 -3652 22856 -3512
rect 13962 -4022 22308 -3882
rect 11772 -4626 11980 -4616
rect 11772 -4810 11780 -4626
rect 11972 -4810 11980 -4626
rect 11772 -4816 11980 -4810
rect 12104 -4758 13660 -4558
rect 12104 -4958 12504 -4758
rect 13260 -4958 13660 -4758
rect 10466 -4970 12504 -4958
rect 10466 -5346 10478 -4970
rect 11224 -5346 12122 -4970
rect 12488 -5346 12504 -4970
rect 10466 -5358 12504 -5346
rect 12918 -4970 13178 -4958
rect 12918 -5346 12924 -4970
rect 13168 -5346 13178 -4970
rect 12918 -5358 13178 -5346
rect 13260 -4970 15296 -4958
rect 13260 -5346 13276 -4970
rect 13642 -5346 14538 -4970
rect 15284 -5346 15296 -4970
rect 13260 -5358 15296 -5346
rect 12998 -5896 13098 -5358
rect 12912 -5906 13330 -5896
rect 2610 -6860 3484 -6740
rect 3364 -6962 3484 -6860
rect 2406 -7174 3158 -6974
rect 2406 -7254 2526 -7174
rect 2722 -7254 2842 -7174
rect 3036 -7254 3158 -7174
rect 3364 -7222 3370 -6962
rect 3478 -7222 3484 -6962
rect 2406 -8054 2412 -7254
rect 2520 -8054 2526 -7254
rect 2564 -8054 2570 -7254
rect 2678 -8054 2684 -7254
rect 2722 -8054 2728 -7254
rect 2836 -8054 2842 -7254
rect 2880 -8054 2886 -7254
rect 2994 -8054 3000 -7254
rect 3036 -8054 3042 -7254
rect 3150 -7554 3158 -7254
rect 3150 -8054 3156 -7554
rect 3196 -8054 3202 -7254
rect 3310 -8054 3316 -7254
rect 2564 -8134 2684 -8054
rect 2880 -8134 3000 -8054
rect 3196 -8134 3316 -8054
rect 2564 -8334 3316 -8134
rect 3364 -7906 3484 -7222
rect 3364 -8166 3370 -7906
rect 3478 -8166 3484 -7906
rect 3614 -6954 3734 -6750
rect 5526 -6810 7682 -6710
rect 11660 -5990 11820 -5984
rect 11660 -6388 11666 -5990
rect 11814 -6388 11820 -5990
rect 11660 -6512 11820 -6388
rect 12912 -6468 12924 -5906
rect 13318 -6468 13330 -5906
rect 12912 -6482 13330 -6468
rect 13948 -5990 14108 -5984
rect 22168 -5990 22308 -4022
rect 22716 -5842 22856 -3652
rect 13948 -6388 13954 -5990
rect 14102 -6388 14108 -5990
rect 22000 -5996 22308 -5990
rect 13948 -6402 14108 -6388
rect 16998 -6106 17298 -6092
rect 16998 -6402 17014 -6106
rect 13948 -6502 17014 -6402
rect 13948 -6512 14108 -6502
rect 11660 -6518 14108 -6512
rect 5526 -6860 5726 -6810
rect 11660 -6916 11666 -6518
rect 11814 -6916 12810 -6518
rect 12958 -6916 13954 -6518
rect 14102 -6916 14108 -6518
rect 11660 -6922 14108 -6916
rect 16036 -6554 16156 -6544
rect 3614 -7214 3620 -6954
rect 3728 -7214 3734 -6954
rect 3614 -7916 3734 -7214
rect 3940 -7174 4692 -6974
rect 3940 -7254 4060 -7174
rect 4256 -7254 4376 -7174
rect 4572 -7254 4692 -7174
rect 3614 -8176 3620 -7916
rect 3728 -8176 3734 -7916
rect 3782 -8054 3790 -7254
rect 3894 -8054 3902 -7254
rect 3940 -8054 3946 -7254
rect 4054 -8054 4060 -7254
rect 4098 -8054 4104 -7254
rect 4212 -8054 4218 -7254
rect 4256 -8054 4262 -7254
rect 4370 -8054 4376 -7254
rect 4414 -8054 4420 -7254
rect 4528 -8054 4534 -7254
rect 4572 -8054 4578 -7254
rect 4686 -8054 4692 -7254
rect 16036 -7036 16044 -6554
rect 16148 -7036 16156 -6554
rect 16998 -6890 17014 -6502
rect 17280 -6890 17298 -6106
rect 22000 -6124 22006 -5996
rect 22302 -6124 22308 -5996
rect 22000 -6130 22308 -6124
rect 22714 -5852 23014 -5842
rect 22714 -6132 22726 -5852
rect 23002 -6132 23014 -5852
rect 24010 -5930 24210 -1292
rect 24004 -6130 24010 -5930
rect 24210 -6130 24216 -5930
rect 22714 -6142 23014 -6132
rect 16998 -6902 17298 -6890
rect 18138 -6554 18258 -6546
rect 16036 -7424 16156 -7036
rect 18138 -7036 18146 -6554
rect 18250 -7036 18258 -6554
rect 16036 -7544 16904 -7424
rect 18138 -7426 18258 -7036
rect 3782 -8134 3902 -8054
rect 4098 -8134 4218 -8054
rect 4414 -8134 4534 -8054
rect 3782 -8334 4534 -8134
rect 7534 -12270 7714 -12260
rect 7534 -12430 7542 -12270
rect 7704 -12272 7714 -12270
rect 9978 -12268 13126 -12252
rect 9978 -12272 9998 -12268
rect 7704 -12428 9998 -12272
rect 7704 -12430 7714 -12428
rect 7534 -12440 7714 -12430
rect 9978 -12434 9998 -12428
rect 11440 -12434 11662 -12268
rect 13104 -12434 13126 -12268
rect 9978 -12452 13126 -12434
rect 7334 -12620 7520 -12612
rect 7334 -12910 7346 -12620
rect 7506 -12910 7520 -12620
rect 7334 -13976 7520 -12910
rect 7334 -13978 9618 -13976
rect 7334 -13986 16552 -13978
rect 7334 -14136 16062 -13986
rect 16542 -14136 16552 -13986
rect 7334 -14146 16552 -14136
rect 7334 -14148 9618 -14146
rect 7334 -14154 7520 -14148
rect 16784 -20684 16904 -7544
rect 17400 -7546 18258 -7426
rect 17400 -20062 17520 -7546
rect 20278 -12298 20478 -12284
rect 20278 -12468 20292 -12298
rect 20464 -12468 20478 -12298
rect 20278 -12484 20478 -12468
rect 19698 -13440 19858 -13426
rect 19698 -13978 19712 -13440
rect 18932 -13994 19712 -13978
rect 18932 -14132 18946 -13994
rect 19348 -14132 19712 -13994
rect 18932 -14146 19712 -14132
rect 19698 -14762 19712 -14146
rect 19844 -14762 19858 -13440
rect 20328 -13896 20478 -12484
rect 22596 -13714 24330 -13688
rect 22596 -13716 23540 -13714
rect 20200 -13906 20600 -13896
rect 20200 -14296 20214 -13906
rect 20590 -14296 20600 -13906
rect 22596 -13924 22612 -13716
rect 23390 -13922 23540 -13716
rect 24318 -13922 24330 -13714
rect 23390 -13924 24330 -13922
rect 22596 -13956 24330 -13924
rect 20200 -14308 20600 -14296
rect 20856 -14030 21760 -14010
rect 20856 -14306 20882 -14030
rect 21736 -14306 21760 -14030
rect 19698 -14776 19858 -14762
rect 20856 -14328 21760 -14306
rect 20856 -15148 20956 -14328
rect 18402 -15164 20956 -15148
rect 18402 -15530 18420 -15164
rect 18784 -15248 20956 -15164
rect 23584 -14938 24274 -13956
rect 18784 -15530 18802 -15248
rect 18402 -15548 18802 -15530
rect 23584 -15592 23628 -14938
rect 24228 -15592 24274 -14938
rect 19854 -16010 21264 -15994
rect 19854 -16020 20476 -16010
rect 19854 -17992 19884 -16020
rect 20222 -16268 20476 -16020
rect 21250 -16268 21264 -16010
rect 20222 -16284 21264 -16268
rect 20222 -16470 20432 -16284
rect 20464 -16324 21704 -16312
rect 20464 -16430 20474 -16324
rect 21252 -16430 21704 -16324
rect 20464 -16442 21704 -16430
rect 20222 -16482 21264 -16470
rect 20222 -16588 20474 -16482
rect 21252 -16588 21264 -16482
rect 20222 -16600 21264 -16588
rect 21296 -16576 21704 -16442
rect 23584 -16576 24274 -15592
rect 21296 -16590 24330 -16576
rect 20222 -16786 20432 -16600
rect 21296 -16628 21718 -16590
rect 20464 -16640 21718 -16628
rect 20464 -16746 20474 -16640
rect 21252 -16746 21718 -16640
rect 20464 -16758 21718 -16746
rect 20222 -16798 21264 -16786
rect 20222 -16904 20474 -16798
rect 21252 -16904 21264 -16798
rect 20222 -16916 21264 -16904
rect 20222 -17102 20432 -16916
rect 21296 -16944 21718 -16758
rect 20464 -16956 21718 -16944
rect 20464 -17062 20474 -16956
rect 21252 -17062 21718 -16956
rect 20464 -17074 21718 -17062
rect 21296 -17098 21718 -17074
rect 22090 -16604 24330 -16590
rect 22090 -16812 22610 -16604
rect 23388 -16812 23540 -16604
rect 24318 -16812 24330 -16604
rect 22090 -16844 24330 -16812
rect 22090 -17098 22104 -16844
rect 20222 -17114 21264 -17102
rect 20222 -17220 20476 -17114
rect 21254 -17220 21264 -17114
rect 20222 -17232 21264 -17220
rect 21296 -17112 22104 -17098
rect 20222 -17418 20432 -17232
rect 21296 -17260 21704 -17112
rect 20464 -17272 21704 -17260
rect 20464 -17378 20474 -17272
rect 21252 -17378 21704 -17272
rect 20464 -17390 21704 -17378
rect 20222 -17430 21264 -17418
rect 20222 -17536 20474 -17430
rect 21252 -17536 21264 -17430
rect 20222 -17548 21264 -17536
rect 20222 -17734 20432 -17548
rect 21296 -17576 21704 -17390
rect 20464 -17588 21704 -17576
rect 20464 -17694 20474 -17588
rect 21252 -17694 21704 -17588
rect 20464 -17706 21704 -17694
rect 20222 -17750 21264 -17734
rect 20222 -17992 20476 -17750
rect 19854 -18008 20476 -17992
rect 21250 -18008 21264 -17750
rect 19854 -18022 21264 -18008
rect 23102 -19984 23402 -19970
rect 23102 -20062 23114 -19984
rect 17400 -20182 23114 -20062
rect 23102 -20260 23114 -20182
rect 23386 -20260 23402 -19984
rect 23102 -20270 23402 -20260
rect 20704 -20606 21004 -20592
rect 20704 -20684 20718 -20606
rect 16784 -20804 20718 -20684
rect 20704 -20882 20718 -20804
rect 20990 -20882 21004 -20606
rect 20704 -20892 21004 -20882
rect 20656 -23312 21056 -23304
rect 20656 -23696 20664 -23312
rect 21048 -23696 21056 -23312
rect 20656 -23704 21056 -23696
rect 23054 -23316 23454 -23304
rect 23054 -23690 23070 -23316
rect 23440 -23690 23454 -23316
rect 23054 -23704 23454 -23690
use sky130_fd_pr__cap_mim_m3_1_67RTNB  amp_XC1
timestamp 1713017924
transform 0 1 12008 -1 0 -4844
box -3798 -4640 3798 4640
use sky130_fd_pr__nfet_g5v0d10v5_ZRJEUR  amp_XM1_2
timestamp 1713024033
transform 1 0 12881 0 1 -5158
box -2451 -458 2451 458
use sky130_fd_pr__pfet_g5v0d10v5_RE37LC  amp_XM3_5
timestamp 1713025933
transform 1 0 17147 0 1 -6497
box -1145 -697 1145 697
use sky130_fd_pr__nfet_01v8_MW6CRE  amp_XM4_18
timestamp 1713025933
transform 1 0 17147 0 1 -5138
box -1083 -610 1083 610
use sky130_fd_pr__pfet_01v8_EDYT7U  amp_XM6
timestamp 1713017924
transform -1 0 19728 0 -1 -6597
box -996 -269 996 269
use sky130_fd_pr__nfet_01v8_UY343Z  amp_XM7
timestamp 1713017924
transform -1 0 19748 0 -1 -5584
box -996 -260 996 260
use sky130_fd_pr__pfet_01v8_EDYT7U  amp_XM8
timestamp 1713017924
transform 0 1 9837 -1 0 -6412
box -996 -269 996 269
use sky130_fd_pr__nfet_01v8_UY343Z  amp_XM9
timestamp 1713017924
transform 0 1 9838 -1 0 -8530
box -996 -260 996 260
use sky130_fd_pr__pfet_01v8_M6QFHF  amp_XM10_12
timestamp 1713033850
transform 1 0 21641 0 1 -6575
box -425 -383 425 383
use sky130_fd_pr__nfet_01v8_6G4XAN  amp_XM11_13
timestamp 1713033850
transform 1 0 21641 0 1 -5561
box -425 -365 425 365
use sky130_fd_pr__pfet_01v8_SV8DF7  amp_XM16_17
timestamp 1713025933
transform 1 0 12884 0 1 -6453
box -2398 -683 2398 683
use sky130_fd_pr__res_xhigh_po_0p35_WHP78W  amp_XR1
timestamp 1713017924
transform 0 1 17636 -1 0 -8635
box -1363 -7182 1363 7182
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  ant_diode_ena
timestamp 1713017924
transform 1 0 2933 0 1 -997
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  ant_diode_standby
timestamp 1713017924
transform 1 0 5403 0 1 -997
box -183 -183 183 183
use sky130_fd_pr__cap_mim_m3_1_VMUSDZ  bias_XC1
timestamp 1713017924
transform 0 -1 13498 1 0 -21238
box -2386 -11800 2386 11800
use sky130_fd_pr__cap_mim_m3_1_WXTTNJ  bias_XC2
timestamp 1713017924
transform 1 0 4162 0 1 -11318
box -2186 -2040 2186 2040
use sky130_fd_pr__cap_mim_m3_1_F5PPB9  bias_XC3
timestamp 1713017924
transform 0 1 9766 -1 0 -16312
box -1986 -7840 1986 7840
use sky130_fd_pr__nfet_g5v0d10v5_RXJTU6  bias_XM1_2
timestamp 1713017924
transform 0 1 20853 -1 0 -14102
box -1584 -1113 1584 1113
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  bias_XM5
timestamp 1713017924
transform 1 0 7426 0 1 -12350
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_H6M2KM  bias_XM6_7_8
timestamp 1713017924
transform -1 0 10726 0 -1 -12352
box -2686 -300 2686 300
use sky130_fd_pr__res_xhigh_po_0p35_M35ED8  bias_XR2
timestamp 1713017924
transform 0 1 10748 -1 0 -15970
box -2276 -8782 2276 8782
use sky130_fd_pr__res_xhigh_po_0p35_VTNT3C  bias_XR3
timestamp 1713017924
transform 0 1 11050 -1 0 -13206
box -450 -8082 450 8082
use sky130_fd_sc_hd__tapvpwrvgnd_1  ena_buf_tap $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1713017924
transform 0 1 2950 -1 0 -1232
box -38 -48 130 592
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  esd_n_xin
timestamp 1713017924
transform 1 0 20505 0 1 -22985
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  esd_n_xout
timestamp 1713017924
transform 1 0 23613 0 1 -22987
box -183 -183 183 183
use sky130_fd_pr__diode_pd2nw_05v5_K4SERG  esd_p_xin
timestamp 1713017924
transform 1 0 21361 0 1 -22975
box -321 -321 321 321
use sky130_fd_pr__diode_pd2nw_05v5_K4SERG  esd_p_xout
timestamp 1713017924
transform 1 0 22787 0 1 -22977
box -321 -321 321 321
use sky130_fd_sc_hd__tapvpwrvgnd_1  standby_buf_tap
timestamp 1713017924
transform 0 -1 5380 1 0 -1324
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1713017924
transform 0 1 2950 -1 0 -1324
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x2
timestamp 1713017924
transform 0 -1 5380 -1 0 -1324
box -38 -48 314 592
use level_shift  x3
timestamp 1713017924
transform 0 1 4250 -1 0 -1190
box 652 -1950 5670 -128
use level_shift  x4
timestamp 1713017924
transform 0 -1 4086 -1 0 -1190
box 652 -1950 5670 -128
use ripl_dly_clk_buf  x7
timestamp 1713017924
transform 1 0 13446 0 1 -1060
box 216 -2416 8990 -156
use sky130_fd_pr__cap_mim_m3_1_KAF84V  XC1
timestamp 1713017924
transform 0 1 13336 -1 0 -12986
box -886 -3440 886 3440
use sky130_fd_pr__cap_mim_m3_1_43FTN9  XC2
timestamp 1713017924
transform 1 0 21712 0 1 -10212
box -3798 -8120 3798 8120
use sky130_fd_pr__cap_mim_m3_1_3DMTNZ  XC3
timestamp 1713017924
transform 1 0 4198 0 1 -5146
box -2492 -2320 2492 2320
use sky130_fd_pr__cap_mim_m3_1_4HHTN9  XC4
timestamp 1713024033
transform 0 -1 11980 1 0 -10184
box -1186 -4640 1186 4640
use sky130_fd_pr__nfet_g5v0d10v5_AB4DGB  XM1
timestamp 1713017924
transform 0 1 20864 -1 0 -17009
box -1147 -658 1147 658
use sky130_fd_pr__pfet_g5v0d10v5_9CUZEG  XM2_bias_XM3_4
timestamp 1713017924
transform 0 1 23465 -1 0 -15266
box -2770 -1161 2770 1161
use sky130_fd_pr__nfet_01v8_AHZR5K  XM3
timestamp 1713017924
transform 0 1 12824 -1 0 -2652
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_HZ6WG7  XM4
timestamp 1713017924
transform 0 1 23509 -1 0 -5548
box -296 -285 296 285
use sky130_fd_pr__nfet_g5v0d10v5_ZPGQJT  XM5
timestamp 1713017924
transform -1 0 2862 0 1 -7654
box -594 -658 594 658
use sky130_fd_pr__pfet_g5v0d10v5_KLKQZ5  XM6
timestamp 1713017924
transform 1 0 4238 0 -1 -7655
box -624 -697 624 697
use sky130_fd_pr__pfet_01v8_3H68VM  XM7
timestamp 1713017924
transform 0 -1 23531 1 0 -6550
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_EDP4SU  XM8
timestamp 1713017924
transform 1 0 8283 0 1 -2587
box -957 -619 957 619
use sky130_fd_pr__pfet_g5v0d10v5_KL3SY6  XM9
timestamp 1713017924
transform -1 0 11530 0 -1 -2569
box -308 -697 308 697
use sky130_fd_pr__nfet_01v8_MLR4K3  XM11
timestamp 1713017924
transform 1 0 10209 0 1 -2592
box -957 -610 957 610
use sky130_fd_pr__res_xhigh_po_0p35_68VL2P  XR2
timestamp 1713017924
transform 0 1 13546 -1 0 -20477
box -2193 -11582 2193 11582
<< labels >>
flabel metal1 7066 -1128 7266 -928 0 FreeSans 256 0 0 0 dvss
port 3 nsew
flabel metal1 2242 -1202 2442 -1002 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 1890 -1200 2090 -1000 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal1 23862 -1102 24062 -902 0 FreeSans 256 0 0 0 dout
port 7 nsew
flabel metal1 21956 -15750 22156 -14384 0 FreeSans 400 0 0 0 vbreg
flabel metal1 22240 -14982 22400 -14170 0 FreeSans 400 0 0 0 vg1
flabel dnwell 19658 -14776 19858 -13426 0 FreeSans 400 0 0 0 vg2
flabel metal1 19698 -14776 19858 -13426 0 FreeSans 400 0 0 0 vg2
flabel metal1 19460 -14978 19640 -13228 0 FreeSans 400 0 0 0 vrb
flabel metal1 24576 -17372 25176 -13160 0 FreeSans 400 0 0 0 avdd_ip
flabel metal2 19854 -18022 20254 -15994 0 FreeSans 400 0 0 0 avss_ip
flabel metal2 7704 -12428 9998 -12272 0 FreeSans 400 0 0 0 icnode
flabel metal2 12998 -5906 13098 -5346 0 FreeSans 400 0 0 0 vbp
flabel metal1 11088 -7256 14680 -7056 0 FreeSans 400 0 0 0 dvdd_ip
flabel metal2 12104 -4758 13660 -4558 0 FreeSans 400 0 0 0 dvss_ip
flabel metal2 13948 -6502 17014 -6402 0 FreeSans 400 0 0 0 tail
flabel metal1 19432 -6734 19978 -5452 0 FreeSans 400 0 0 0 inv_in
flabel metal1 20574 -6654 20674 -5530 0 FreeSans 400 0 0 0 inv_m1
flabel metal1 21290 -6516 21390 -5610 0 FreeSans 400 0 0 0 inv_m2
flabel metal1 16648 -6900 16728 -4734 0 FreeSans 400 0 0 0 vn
flabel metal1 17564 -6898 17644 -4734 0 FreeSans 400 0 0 0 xin_buf
flabel metal1 21900 -6738 22000 -5406 0 FreeSans 400 0 0 0 dout_ip
flabel metal2 20656 -23704 21056 -23304 0 FreeSans 1600 0 0 0 xin
port 10 nsew
flabel metal2 23054 -23704 23454 -23304 0 FreeSans 1600 0 0 0 xout
port 11 nsew
flabel metal2 22716 -5852 22856 -3512 0 FreeSans 400 0 0 0 dout_filt
flabel metal2 3614 -7916 3734 -7214 0 FreeSans 400 0 0 0 ena_b_33
flabel metal2 3364 -7906 3484 -7222 0 FreeSans 400 0 0 0 ena_33
flabel metal2 2564 -8334 3316 -8134 0 FreeSans 400 0 0 0 avss_ip
flabel metal2 3782 -8334 4534 -8134 0 FreeSans 400 0 0 0 avdd_ip
flabel metal2 7582 -6810 7682 -3808 0 FreeSans 400 0 0 0 standby_33
flabel metal1 9798 -1130 9998 -930 0 FreeSans 256 0 0 0 dvdd
port 2 nsew
flabel metal1 11388 -1196 11588 -996 0 FreeSans 256 0 0 0 ibias
port 4 nsew
flabel metal2 4338 -1212 4738 -812 0 FreeSans 1200 0 0 0 standby
port 9 nsew
flabel metal2 3592 -1212 3992 -812 0 FreeSans 1200 0 0 0 ena
port 8 nsew
<< end >>
