magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< pwell >>
rect -4268 -4582 4268 4582
<< psubdiff >>
rect -4232 4512 -4136 4546
rect 4136 4512 4232 4546
rect -4232 4450 -4198 4512
rect 4198 4450 4232 4512
rect -4232 -4512 -4198 -4450
rect 4198 -4512 4232 -4450
rect -4232 -4546 -4136 -4512
rect 4136 -4546 4232 -4512
<< psubdiffcont >>
rect -4136 4512 4136 4546
rect -4232 -4450 -4198 4450
rect 4198 -4450 4232 4450
rect -4136 -4546 4136 -4512
<< xpolycontact >>
rect -4102 3984 -4032 4416
rect -4102 -4416 -4032 -3984
rect -3936 3984 -3866 4416
rect -3936 -4416 -3866 -3984
rect -3770 3984 -3700 4416
rect -3770 -4416 -3700 -3984
rect -3604 3984 -3534 4416
rect -3604 -4416 -3534 -3984
rect -3438 3984 -3368 4416
rect -3438 -4416 -3368 -3984
rect -3272 3984 -3202 4416
rect -3272 -4416 -3202 -3984
rect -3106 3984 -3036 4416
rect -3106 -4416 -3036 -3984
rect -2940 3984 -2870 4416
rect -2940 -4416 -2870 -3984
rect -2774 3984 -2704 4416
rect -2774 -4416 -2704 -3984
rect -2608 3984 -2538 4416
rect -2608 -4416 -2538 -3984
rect -2442 3984 -2372 4416
rect -2442 -4416 -2372 -3984
rect -2276 3984 -2206 4416
rect -2276 -4416 -2206 -3984
rect -2110 3984 -2040 4416
rect -2110 -4416 -2040 -3984
rect -1944 3984 -1874 4416
rect -1944 -4416 -1874 -3984
rect -1778 3984 -1708 4416
rect -1778 -4416 -1708 -3984
rect -1612 3984 -1542 4416
rect -1612 -4416 -1542 -3984
rect -1446 3984 -1376 4416
rect -1446 -4416 -1376 -3984
rect -1280 3984 -1210 4416
rect -1280 -4416 -1210 -3984
rect -1114 3984 -1044 4416
rect -1114 -4416 -1044 -3984
rect -948 3984 -878 4416
rect -948 -4416 -878 -3984
rect -782 3984 -712 4416
rect -782 -4416 -712 -3984
rect -616 3984 -546 4416
rect -616 -4416 -546 -3984
rect -450 3984 -380 4416
rect -450 -4416 -380 -3984
rect -284 3984 -214 4416
rect -284 -4416 -214 -3984
rect -118 3984 -48 4416
rect -118 -4416 -48 -3984
rect 48 3984 118 4416
rect 48 -4416 118 -3984
rect 214 3984 284 4416
rect 214 -4416 284 -3984
rect 380 3984 450 4416
rect 380 -4416 450 -3984
rect 546 3984 616 4416
rect 546 -4416 616 -3984
rect 712 3984 782 4416
rect 712 -4416 782 -3984
rect 878 3984 948 4416
rect 878 -4416 948 -3984
rect 1044 3984 1114 4416
rect 1044 -4416 1114 -3984
rect 1210 3984 1280 4416
rect 1210 -4416 1280 -3984
rect 1376 3984 1446 4416
rect 1376 -4416 1446 -3984
rect 1542 3984 1612 4416
rect 1542 -4416 1612 -3984
rect 1708 3984 1778 4416
rect 1708 -4416 1778 -3984
rect 1874 3984 1944 4416
rect 1874 -4416 1944 -3984
rect 2040 3984 2110 4416
rect 2040 -4416 2110 -3984
rect 2206 3984 2276 4416
rect 2206 -4416 2276 -3984
rect 2372 3984 2442 4416
rect 2372 -4416 2442 -3984
rect 2538 3984 2608 4416
rect 2538 -4416 2608 -3984
rect 2704 3984 2774 4416
rect 2704 -4416 2774 -3984
rect 2870 3984 2940 4416
rect 2870 -4416 2940 -3984
rect 3036 3984 3106 4416
rect 3036 -4416 3106 -3984
rect 3202 3984 3272 4416
rect 3202 -4416 3272 -3984
rect 3368 3984 3438 4416
rect 3368 -4416 3438 -3984
rect 3534 3984 3604 4416
rect 3534 -4416 3604 -3984
rect 3700 3984 3770 4416
rect 3700 -4416 3770 -3984
rect 3866 3984 3936 4416
rect 3866 -4416 3936 -3984
rect 4032 3984 4102 4416
rect 4032 -4416 4102 -3984
<< xpolyres >>
rect -4102 -3984 -4032 3984
rect -3936 -3984 -3866 3984
rect -3770 -3984 -3700 3984
rect -3604 -3984 -3534 3984
rect -3438 -3984 -3368 3984
rect -3272 -3984 -3202 3984
rect -3106 -3984 -3036 3984
rect -2940 -3984 -2870 3984
rect -2774 -3984 -2704 3984
rect -2608 -3984 -2538 3984
rect -2442 -3984 -2372 3984
rect -2276 -3984 -2206 3984
rect -2110 -3984 -2040 3984
rect -1944 -3984 -1874 3984
rect -1778 -3984 -1708 3984
rect -1612 -3984 -1542 3984
rect -1446 -3984 -1376 3984
rect -1280 -3984 -1210 3984
rect -1114 -3984 -1044 3984
rect -948 -3984 -878 3984
rect -782 -3984 -712 3984
rect -616 -3984 -546 3984
rect -450 -3984 -380 3984
rect -284 -3984 -214 3984
rect -118 -3984 -48 3984
rect 48 -3984 118 3984
rect 214 -3984 284 3984
rect 380 -3984 450 3984
rect 546 -3984 616 3984
rect 712 -3984 782 3984
rect 878 -3984 948 3984
rect 1044 -3984 1114 3984
rect 1210 -3984 1280 3984
rect 1376 -3984 1446 3984
rect 1542 -3984 1612 3984
rect 1708 -3984 1778 3984
rect 1874 -3984 1944 3984
rect 2040 -3984 2110 3984
rect 2206 -3984 2276 3984
rect 2372 -3984 2442 3984
rect 2538 -3984 2608 3984
rect 2704 -3984 2774 3984
rect 2870 -3984 2940 3984
rect 3036 -3984 3106 3984
rect 3202 -3984 3272 3984
rect 3368 -3984 3438 3984
rect 3534 -3984 3604 3984
rect 3700 -3984 3770 3984
rect 3866 -3984 3936 3984
rect 4032 -3984 4102 3984
<< locali >>
rect -4232 4512 -4136 4546
rect 4136 4512 4232 4546
rect -4232 4450 -4198 4512
rect 4198 4450 4232 4512
rect -4232 -4512 -4198 -4450
rect 4198 -4512 4232 -4450
rect -4232 -4546 -4136 -4512
rect 4136 -4546 4232 -4512
<< viali >>
rect -4086 4001 -4048 4398
rect -3920 4001 -3882 4398
rect -3754 4001 -3716 4398
rect -3588 4001 -3550 4398
rect -3422 4001 -3384 4398
rect -3256 4001 -3218 4398
rect -3090 4001 -3052 4398
rect -2924 4001 -2886 4398
rect -2758 4001 -2720 4398
rect -2592 4001 -2554 4398
rect -2426 4001 -2388 4398
rect -2260 4001 -2222 4398
rect -2094 4001 -2056 4398
rect -1928 4001 -1890 4398
rect -1762 4001 -1724 4398
rect -1596 4001 -1558 4398
rect -1430 4001 -1392 4398
rect -1264 4001 -1226 4398
rect -1098 4001 -1060 4398
rect -932 4001 -894 4398
rect -766 4001 -728 4398
rect -600 4001 -562 4398
rect -434 4001 -396 4398
rect -268 4001 -230 4398
rect -102 4001 -64 4398
rect 64 4001 102 4398
rect 230 4001 268 4398
rect 396 4001 434 4398
rect 562 4001 600 4398
rect 728 4001 766 4398
rect 894 4001 932 4398
rect 1060 4001 1098 4398
rect 1226 4001 1264 4398
rect 1392 4001 1430 4398
rect 1558 4001 1596 4398
rect 1724 4001 1762 4398
rect 1890 4001 1928 4398
rect 2056 4001 2094 4398
rect 2222 4001 2260 4398
rect 2388 4001 2426 4398
rect 2554 4001 2592 4398
rect 2720 4001 2758 4398
rect 2886 4001 2924 4398
rect 3052 4001 3090 4398
rect 3218 4001 3256 4398
rect 3384 4001 3422 4398
rect 3550 4001 3588 4398
rect 3716 4001 3754 4398
rect 3882 4001 3920 4398
rect 4048 4001 4086 4398
rect -4086 -4398 -4048 -4001
rect -3920 -4398 -3882 -4001
rect -3754 -4398 -3716 -4001
rect -3588 -4398 -3550 -4001
rect -3422 -4398 -3384 -4001
rect -3256 -4398 -3218 -4001
rect -3090 -4398 -3052 -4001
rect -2924 -4398 -2886 -4001
rect -2758 -4398 -2720 -4001
rect -2592 -4398 -2554 -4001
rect -2426 -4398 -2388 -4001
rect -2260 -4398 -2222 -4001
rect -2094 -4398 -2056 -4001
rect -1928 -4398 -1890 -4001
rect -1762 -4398 -1724 -4001
rect -1596 -4398 -1558 -4001
rect -1430 -4398 -1392 -4001
rect -1264 -4398 -1226 -4001
rect -1098 -4398 -1060 -4001
rect -932 -4398 -894 -4001
rect -766 -4398 -728 -4001
rect -600 -4398 -562 -4001
rect -434 -4398 -396 -4001
rect -268 -4398 -230 -4001
rect -102 -4398 -64 -4001
rect 64 -4398 102 -4001
rect 230 -4398 268 -4001
rect 396 -4398 434 -4001
rect 562 -4398 600 -4001
rect 728 -4398 766 -4001
rect 894 -4398 932 -4001
rect 1060 -4398 1098 -4001
rect 1226 -4398 1264 -4001
rect 1392 -4398 1430 -4001
rect 1558 -4398 1596 -4001
rect 1724 -4398 1762 -4001
rect 1890 -4398 1928 -4001
rect 2056 -4398 2094 -4001
rect 2222 -4398 2260 -4001
rect 2388 -4398 2426 -4001
rect 2554 -4398 2592 -4001
rect 2720 -4398 2758 -4001
rect 2886 -4398 2924 -4001
rect 3052 -4398 3090 -4001
rect 3218 -4398 3256 -4001
rect 3384 -4398 3422 -4001
rect 3550 -4398 3588 -4001
rect 3716 -4398 3754 -4001
rect 3882 -4398 3920 -4001
rect 4048 -4398 4086 -4001
<< metal1 >>
rect -4092 4398 -4042 4410
rect -4092 4001 -4086 4398
rect -4048 4001 -4042 4398
rect -4092 3989 -4042 4001
rect -3926 4398 -3876 4410
rect -3926 4001 -3920 4398
rect -3882 4001 -3876 4398
rect -3926 3989 -3876 4001
rect -3760 4398 -3710 4410
rect -3760 4001 -3754 4398
rect -3716 4001 -3710 4398
rect -3760 3989 -3710 4001
rect -3594 4398 -3544 4410
rect -3594 4001 -3588 4398
rect -3550 4001 -3544 4398
rect -3594 3989 -3544 4001
rect -3428 4398 -3378 4410
rect -3428 4001 -3422 4398
rect -3384 4001 -3378 4398
rect -3428 3989 -3378 4001
rect -3262 4398 -3212 4410
rect -3262 4001 -3256 4398
rect -3218 4001 -3212 4398
rect -3262 3989 -3212 4001
rect -3096 4398 -3046 4410
rect -3096 4001 -3090 4398
rect -3052 4001 -3046 4398
rect -3096 3989 -3046 4001
rect -2930 4398 -2880 4410
rect -2930 4001 -2924 4398
rect -2886 4001 -2880 4398
rect -2930 3989 -2880 4001
rect -2764 4398 -2714 4410
rect -2764 4001 -2758 4398
rect -2720 4001 -2714 4398
rect -2764 3989 -2714 4001
rect -2598 4398 -2548 4410
rect -2598 4001 -2592 4398
rect -2554 4001 -2548 4398
rect -2598 3989 -2548 4001
rect -2432 4398 -2382 4410
rect -2432 4001 -2426 4398
rect -2388 4001 -2382 4398
rect -2432 3989 -2382 4001
rect -2266 4398 -2216 4410
rect -2266 4001 -2260 4398
rect -2222 4001 -2216 4398
rect -2266 3989 -2216 4001
rect -2100 4398 -2050 4410
rect -2100 4001 -2094 4398
rect -2056 4001 -2050 4398
rect -2100 3989 -2050 4001
rect -1934 4398 -1884 4410
rect -1934 4001 -1928 4398
rect -1890 4001 -1884 4398
rect -1934 3989 -1884 4001
rect -1768 4398 -1718 4410
rect -1768 4001 -1762 4398
rect -1724 4001 -1718 4398
rect -1768 3989 -1718 4001
rect -1602 4398 -1552 4410
rect -1602 4001 -1596 4398
rect -1558 4001 -1552 4398
rect -1602 3989 -1552 4001
rect -1436 4398 -1386 4410
rect -1436 4001 -1430 4398
rect -1392 4001 -1386 4398
rect -1436 3989 -1386 4001
rect -1270 4398 -1220 4410
rect -1270 4001 -1264 4398
rect -1226 4001 -1220 4398
rect -1270 3989 -1220 4001
rect -1104 4398 -1054 4410
rect -1104 4001 -1098 4398
rect -1060 4001 -1054 4398
rect -1104 3989 -1054 4001
rect -938 4398 -888 4410
rect -938 4001 -932 4398
rect -894 4001 -888 4398
rect -938 3989 -888 4001
rect -772 4398 -722 4410
rect -772 4001 -766 4398
rect -728 4001 -722 4398
rect -772 3989 -722 4001
rect -606 4398 -556 4410
rect -606 4001 -600 4398
rect -562 4001 -556 4398
rect -606 3989 -556 4001
rect -440 4398 -390 4410
rect -440 4001 -434 4398
rect -396 4001 -390 4398
rect -440 3989 -390 4001
rect -274 4398 -224 4410
rect -274 4001 -268 4398
rect -230 4001 -224 4398
rect -274 3989 -224 4001
rect -108 4398 -58 4410
rect -108 4001 -102 4398
rect -64 4001 -58 4398
rect -108 3989 -58 4001
rect 58 4398 108 4410
rect 58 4001 64 4398
rect 102 4001 108 4398
rect 58 3989 108 4001
rect 224 4398 274 4410
rect 224 4001 230 4398
rect 268 4001 274 4398
rect 224 3989 274 4001
rect 390 4398 440 4410
rect 390 4001 396 4398
rect 434 4001 440 4398
rect 390 3989 440 4001
rect 556 4398 606 4410
rect 556 4001 562 4398
rect 600 4001 606 4398
rect 556 3989 606 4001
rect 722 4398 772 4410
rect 722 4001 728 4398
rect 766 4001 772 4398
rect 722 3989 772 4001
rect 888 4398 938 4410
rect 888 4001 894 4398
rect 932 4001 938 4398
rect 888 3989 938 4001
rect 1054 4398 1104 4410
rect 1054 4001 1060 4398
rect 1098 4001 1104 4398
rect 1054 3989 1104 4001
rect 1220 4398 1270 4410
rect 1220 4001 1226 4398
rect 1264 4001 1270 4398
rect 1220 3989 1270 4001
rect 1386 4398 1436 4410
rect 1386 4001 1392 4398
rect 1430 4001 1436 4398
rect 1386 3989 1436 4001
rect 1552 4398 1602 4410
rect 1552 4001 1558 4398
rect 1596 4001 1602 4398
rect 1552 3989 1602 4001
rect 1718 4398 1768 4410
rect 1718 4001 1724 4398
rect 1762 4001 1768 4398
rect 1718 3989 1768 4001
rect 1884 4398 1934 4410
rect 1884 4001 1890 4398
rect 1928 4001 1934 4398
rect 1884 3989 1934 4001
rect 2050 4398 2100 4410
rect 2050 4001 2056 4398
rect 2094 4001 2100 4398
rect 2050 3989 2100 4001
rect 2216 4398 2266 4410
rect 2216 4001 2222 4398
rect 2260 4001 2266 4398
rect 2216 3989 2266 4001
rect 2382 4398 2432 4410
rect 2382 4001 2388 4398
rect 2426 4001 2432 4398
rect 2382 3989 2432 4001
rect 2548 4398 2598 4410
rect 2548 4001 2554 4398
rect 2592 4001 2598 4398
rect 2548 3989 2598 4001
rect 2714 4398 2764 4410
rect 2714 4001 2720 4398
rect 2758 4001 2764 4398
rect 2714 3989 2764 4001
rect 2880 4398 2930 4410
rect 2880 4001 2886 4398
rect 2924 4001 2930 4398
rect 2880 3989 2930 4001
rect 3046 4398 3096 4410
rect 3046 4001 3052 4398
rect 3090 4001 3096 4398
rect 3046 3989 3096 4001
rect 3212 4398 3262 4410
rect 3212 4001 3218 4398
rect 3256 4001 3262 4398
rect 3212 3989 3262 4001
rect 3378 4398 3428 4410
rect 3378 4001 3384 4398
rect 3422 4001 3428 4398
rect 3378 3989 3428 4001
rect 3544 4398 3594 4410
rect 3544 4001 3550 4398
rect 3588 4001 3594 4398
rect 3544 3989 3594 4001
rect 3710 4398 3760 4410
rect 3710 4001 3716 4398
rect 3754 4001 3760 4398
rect 3710 3989 3760 4001
rect 3876 4398 3926 4410
rect 3876 4001 3882 4398
rect 3920 4001 3926 4398
rect 3876 3989 3926 4001
rect 4042 4398 4092 4410
rect 4042 4001 4048 4398
rect 4086 4001 4092 4398
rect 4042 3989 4092 4001
rect -4092 -4001 -4042 -3989
rect -4092 -4398 -4086 -4001
rect -4048 -4398 -4042 -4001
rect -4092 -4410 -4042 -4398
rect -3926 -4001 -3876 -3989
rect -3926 -4398 -3920 -4001
rect -3882 -4398 -3876 -4001
rect -3926 -4410 -3876 -4398
rect -3760 -4001 -3710 -3989
rect -3760 -4398 -3754 -4001
rect -3716 -4398 -3710 -4001
rect -3760 -4410 -3710 -4398
rect -3594 -4001 -3544 -3989
rect -3594 -4398 -3588 -4001
rect -3550 -4398 -3544 -4001
rect -3594 -4410 -3544 -4398
rect -3428 -4001 -3378 -3989
rect -3428 -4398 -3422 -4001
rect -3384 -4398 -3378 -4001
rect -3428 -4410 -3378 -4398
rect -3262 -4001 -3212 -3989
rect -3262 -4398 -3256 -4001
rect -3218 -4398 -3212 -4001
rect -3262 -4410 -3212 -4398
rect -3096 -4001 -3046 -3989
rect -3096 -4398 -3090 -4001
rect -3052 -4398 -3046 -4001
rect -3096 -4410 -3046 -4398
rect -2930 -4001 -2880 -3989
rect -2930 -4398 -2924 -4001
rect -2886 -4398 -2880 -4001
rect -2930 -4410 -2880 -4398
rect -2764 -4001 -2714 -3989
rect -2764 -4398 -2758 -4001
rect -2720 -4398 -2714 -4001
rect -2764 -4410 -2714 -4398
rect -2598 -4001 -2548 -3989
rect -2598 -4398 -2592 -4001
rect -2554 -4398 -2548 -4001
rect -2598 -4410 -2548 -4398
rect -2432 -4001 -2382 -3989
rect -2432 -4398 -2426 -4001
rect -2388 -4398 -2382 -4001
rect -2432 -4410 -2382 -4398
rect -2266 -4001 -2216 -3989
rect -2266 -4398 -2260 -4001
rect -2222 -4398 -2216 -4001
rect -2266 -4410 -2216 -4398
rect -2100 -4001 -2050 -3989
rect -2100 -4398 -2094 -4001
rect -2056 -4398 -2050 -4001
rect -2100 -4410 -2050 -4398
rect -1934 -4001 -1884 -3989
rect -1934 -4398 -1928 -4001
rect -1890 -4398 -1884 -4001
rect -1934 -4410 -1884 -4398
rect -1768 -4001 -1718 -3989
rect -1768 -4398 -1762 -4001
rect -1724 -4398 -1718 -4001
rect -1768 -4410 -1718 -4398
rect -1602 -4001 -1552 -3989
rect -1602 -4398 -1596 -4001
rect -1558 -4398 -1552 -4001
rect -1602 -4410 -1552 -4398
rect -1436 -4001 -1386 -3989
rect -1436 -4398 -1430 -4001
rect -1392 -4398 -1386 -4001
rect -1436 -4410 -1386 -4398
rect -1270 -4001 -1220 -3989
rect -1270 -4398 -1264 -4001
rect -1226 -4398 -1220 -4001
rect -1270 -4410 -1220 -4398
rect -1104 -4001 -1054 -3989
rect -1104 -4398 -1098 -4001
rect -1060 -4398 -1054 -4001
rect -1104 -4410 -1054 -4398
rect -938 -4001 -888 -3989
rect -938 -4398 -932 -4001
rect -894 -4398 -888 -4001
rect -938 -4410 -888 -4398
rect -772 -4001 -722 -3989
rect -772 -4398 -766 -4001
rect -728 -4398 -722 -4001
rect -772 -4410 -722 -4398
rect -606 -4001 -556 -3989
rect -606 -4398 -600 -4001
rect -562 -4398 -556 -4001
rect -606 -4410 -556 -4398
rect -440 -4001 -390 -3989
rect -440 -4398 -434 -4001
rect -396 -4398 -390 -4001
rect -440 -4410 -390 -4398
rect -274 -4001 -224 -3989
rect -274 -4398 -268 -4001
rect -230 -4398 -224 -4001
rect -274 -4410 -224 -4398
rect -108 -4001 -58 -3989
rect -108 -4398 -102 -4001
rect -64 -4398 -58 -4001
rect -108 -4410 -58 -4398
rect 58 -4001 108 -3989
rect 58 -4398 64 -4001
rect 102 -4398 108 -4001
rect 58 -4410 108 -4398
rect 224 -4001 274 -3989
rect 224 -4398 230 -4001
rect 268 -4398 274 -4001
rect 224 -4410 274 -4398
rect 390 -4001 440 -3989
rect 390 -4398 396 -4001
rect 434 -4398 440 -4001
rect 390 -4410 440 -4398
rect 556 -4001 606 -3989
rect 556 -4398 562 -4001
rect 600 -4398 606 -4001
rect 556 -4410 606 -4398
rect 722 -4001 772 -3989
rect 722 -4398 728 -4001
rect 766 -4398 772 -4001
rect 722 -4410 772 -4398
rect 888 -4001 938 -3989
rect 888 -4398 894 -4001
rect 932 -4398 938 -4001
rect 888 -4410 938 -4398
rect 1054 -4001 1104 -3989
rect 1054 -4398 1060 -4001
rect 1098 -4398 1104 -4001
rect 1054 -4410 1104 -4398
rect 1220 -4001 1270 -3989
rect 1220 -4398 1226 -4001
rect 1264 -4398 1270 -4001
rect 1220 -4410 1270 -4398
rect 1386 -4001 1436 -3989
rect 1386 -4398 1392 -4001
rect 1430 -4398 1436 -4001
rect 1386 -4410 1436 -4398
rect 1552 -4001 1602 -3989
rect 1552 -4398 1558 -4001
rect 1596 -4398 1602 -4001
rect 1552 -4410 1602 -4398
rect 1718 -4001 1768 -3989
rect 1718 -4398 1724 -4001
rect 1762 -4398 1768 -4001
rect 1718 -4410 1768 -4398
rect 1884 -4001 1934 -3989
rect 1884 -4398 1890 -4001
rect 1928 -4398 1934 -4001
rect 1884 -4410 1934 -4398
rect 2050 -4001 2100 -3989
rect 2050 -4398 2056 -4001
rect 2094 -4398 2100 -4001
rect 2050 -4410 2100 -4398
rect 2216 -4001 2266 -3989
rect 2216 -4398 2222 -4001
rect 2260 -4398 2266 -4001
rect 2216 -4410 2266 -4398
rect 2382 -4001 2432 -3989
rect 2382 -4398 2388 -4001
rect 2426 -4398 2432 -4001
rect 2382 -4410 2432 -4398
rect 2548 -4001 2598 -3989
rect 2548 -4398 2554 -4001
rect 2592 -4398 2598 -4001
rect 2548 -4410 2598 -4398
rect 2714 -4001 2764 -3989
rect 2714 -4398 2720 -4001
rect 2758 -4398 2764 -4001
rect 2714 -4410 2764 -4398
rect 2880 -4001 2930 -3989
rect 2880 -4398 2886 -4001
rect 2924 -4398 2930 -4001
rect 2880 -4410 2930 -4398
rect 3046 -4001 3096 -3989
rect 3046 -4398 3052 -4001
rect 3090 -4398 3096 -4001
rect 3046 -4410 3096 -4398
rect 3212 -4001 3262 -3989
rect 3212 -4398 3218 -4001
rect 3256 -4398 3262 -4001
rect 3212 -4410 3262 -4398
rect 3378 -4001 3428 -3989
rect 3378 -4398 3384 -4001
rect 3422 -4398 3428 -4001
rect 3378 -4410 3428 -4398
rect 3544 -4001 3594 -3989
rect 3544 -4398 3550 -4001
rect 3588 -4398 3594 -4001
rect 3544 -4410 3594 -4398
rect 3710 -4001 3760 -3989
rect 3710 -4398 3716 -4001
rect 3754 -4398 3760 -4001
rect 3710 -4410 3760 -4398
rect 3876 -4001 3926 -3989
rect 3876 -4398 3882 -4001
rect 3920 -4398 3926 -4001
rect 3876 -4410 3926 -4398
rect 4042 -4001 4092 -3989
rect 4042 -4398 4048 -4001
rect 4086 -4398 4092 -4001
rect 4042 -4410 4092 -4398
<< properties >>
string FIXED_BBOX -4215 -4529 4215 4529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 40.0 m 1 nx 50 wmin 0.350 lmin 0.50 rho 2000 val 229.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
