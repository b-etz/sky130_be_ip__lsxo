magic
tech sky130A
magscale 1 2
timestamp 1712854380
<< metal3 >>
rect -2492 6812 -120 6840
rect -2492 4788 -204 6812
rect -140 4788 -120 6812
rect -2492 4760 -120 4788
rect 120 6812 2492 6840
rect 120 4788 2408 6812
rect 2472 4788 2492 6812
rect 120 4760 2492 4788
rect -2492 4492 -120 4520
rect -2492 2468 -204 4492
rect -140 2468 -120 4492
rect -2492 2440 -120 2468
rect 120 4492 2492 4520
rect 120 2468 2408 4492
rect 2472 2468 2492 4492
rect 120 2440 2492 2468
rect -2492 2172 -120 2200
rect -2492 148 -204 2172
rect -140 148 -120 2172
rect -2492 120 -120 148
rect 120 2172 2492 2200
rect 120 148 2408 2172
rect 2472 148 2492 2172
rect 120 120 2492 148
rect -2492 -148 -120 -120
rect -2492 -2172 -204 -148
rect -140 -2172 -120 -148
rect -2492 -2200 -120 -2172
rect 120 -148 2492 -120
rect 120 -2172 2408 -148
rect 2472 -2172 2492 -148
rect 120 -2200 2492 -2172
rect -2492 -2468 -120 -2440
rect -2492 -4492 -204 -2468
rect -140 -4492 -120 -2468
rect -2492 -4520 -120 -4492
rect 120 -2468 2492 -2440
rect 120 -4492 2408 -2468
rect 2472 -4492 2492 -2468
rect 120 -4520 2492 -4492
rect -2492 -4788 -120 -4760
rect -2492 -6812 -204 -4788
rect -140 -6812 -120 -4788
rect -2492 -6840 -120 -6812
rect 120 -4788 2492 -4760
rect 120 -6812 2408 -4788
rect 2472 -6812 2492 -4788
rect 120 -6840 2492 -6812
<< via3 >>
rect -204 4788 -140 6812
rect 2408 4788 2472 6812
rect -204 2468 -140 4492
rect 2408 2468 2472 4492
rect -204 148 -140 2172
rect 2408 148 2472 2172
rect -204 -2172 -140 -148
rect 2408 -2172 2472 -148
rect -204 -4492 -140 -2468
rect 2408 -4492 2472 -2468
rect -204 -6812 -140 -4788
rect 2408 -6812 2472 -4788
<< mimcap >>
rect -2452 6760 -452 6800
rect -2452 4840 -2412 6760
rect -492 4840 -452 6760
rect -2452 4800 -452 4840
rect 160 6760 2160 6800
rect 160 4840 200 6760
rect 2120 4840 2160 6760
rect 160 4800 2160 4840
rect -2452 4440 -452 4480
rect -2452 2520 -2412 4440
rect -492 2520 -452 4440
rect -2452 2480 -452 2520
rect 160 4440 2160 4480
rect 160 2520 200 4440
rect 2120 2520 2160 4440
rect 160 2480 2160 2520
rect -2452 2120 -452 2160
rect -2452 200 -2412 2120
rect -492 200 -452 2120
rect -2452 160 -452 200
rect 160 2120 2160 2160
rect 160 200 200 2120
rect 2120 200 2160 2120
rect 160 160 2160 200
rect -2452 -200 -452 -160
rect -2452 -2120 -2412 -200
rect -492 -2120 -452 -200
rect -2452 -2160 -452 -2120
rect 160 -200 2160 -160
rect 160 -2120 200 -200
rect 2120 -2120 2160 -200
rect 160 -2160 2160 -2120
rect -2452 -2520 -452 -2480
rect -2452 -4440 -2412 -2520
rect -492 -4440 -452 -2520
rect -2452 -4480 -452 -4440
rect 160 -2520 2160 -2480
rect 160 -4440 200 -2520
rect 2120 -4440 2160 -2520
rect 160 -4480 2160 -4440
rect -2452 -4840 -452 -4800
rect -2452 -6760 -2412 -4840
rect -492 -6760 -452 -4840
rect -2452 -6800 -452 -6760
rect 160 -4840 2160 -4800
rect 160 -6760 200 -4840
rect 2120 -6760 2160 -4840
rect 160 -6800 2160 -6760
<< mimcapcontact >>
rect -2412 4840 -492 6760
rect 200 4840 2120 6760
rect -2412 2520 -492 4440
rect 200 2520 2120 4440
rect -2412 200 -492 2120
rect 200 200 2120 2120
rect -2412 -2120 -492 -200
rect 200 -2120 2120 -200
rect -2412 -4440 -492 -2520
rect 200 -4440 2120 -2520
rect -2412 -6760 -492 -4840
rect 200 -6760 2120 -4840
<< metal4 >>
rect -1504 6761 -1400 6960
rect -224 6812 -120 6960
rect -2413 6760 -491 6761
rect -2413 4840 -2412 6760
rect -492 4840 -491 6760
rect -2413 4839 -491 4840
rect -1504 4441 -1400 4839
rect -224 4788 -204 6812
rect -140 4788 -120 6812
rect 1108 6761 1212 6960
rect 2388 6812 2492 6960
rect 199 6760 2121 6761
rect 199 4840 200 6760
rect 2120 4840 2121 6760
rect 199 4839 2121 4840
rect -224 4492 -120 4788
rect -2413 4440 -491 4441
rect -2413 2520 -2412 4440
rect -492 2520 -491 4440
rect -2413 2519 -491 2520
rect -1504 2121 -1400 2519
rect -224 2468 -204 4492
rect -140 2468 -120 4492
rect 1108 4441 1212 4839
rect 2388 4788 2408 6812
rect 2472 4788 2492 6812
rect 2388 4492 2492 4788
rect 199 4440 2121 4441
rect 199 2520 200 4440
rect 2120 2520 2121 4440
rect 199 2519 2121 2520
rect -224 2172 -120 2468
rect -2413 2120 -491 2121
rect -2413 200 -2412 2120
rect -492 200 -491 2120
rect -2413 199 -491 200
rect -1504 -199 -1400 199
rect -224 148 -204 2172
rect -140 148 -120 2172
rect 1108 2121 1212 2519
rect 2388 2468 2408 4492
rect 2472 2468 2492 4492
rect 2388 2172 2492 2468
rect 199 2120 2121 2121
rect 199 200 200 2120
rect 2120 200 2121 2120
rect 199 199 2121 200
rect -224 -148 -120 148
rect -2413 -200 -491 -199
rect -2413 -2120 -2412 -200
rect -492 -2120 -491 -200
rect -2413 -2121 -491 -2120
rect -1504 -2519 -1400 -2121
rect -224 -2172 -204 -148
rect -140 -2172 -120 -148
rect 1108 -199 1212 199
rect 2388 148 2408 2172
rect 2472 148 2492 2172
rect 2388 -148 2492 148
rect 199 -200 2121 -199
rect 199 -2120 200 -200
rect 2120 -2120 2121 -200
rect 199 -2121 2121 -2120
rect -224 -2468 -120 -2172
rect -2413 -2520 -491 -2519
rect -2413 -4440 -2412 -2520
rect -492 -4440 -491 -2520
rect -2413 -4441 -491 -4440
rect -1504 -4839 -1400 -4441
rect -224 -4492 -204 -2468
rect -140 -4492 -120 -2468
rect 1108 -2519 1212 -2121
rect 2388 -2172 2408 -148
rect 2472 -2172 2492 -148
rect 2388 -2468 2492 -2172
rect 199 -2520 2121 -2519
rect 199 -4440 200 -2520
rect 2120 -4440 2121 -2520
rect 199 -4441 2121 -4440
rect -224 -4788 -120 -4492
rect -2413 -4840 -491 -4839
rect -2413 -6760 -2412 -4840
rect -492 -6760 -491 -4840
rect -2413 -6761 -491 -6760
rect -1504 -6960 -1400 -6761
rect -224 -6812 -204 -4788
rect -140 -6812 -120 -4788
rect 1108 -4839 1212 -4441
rect 2388 -4492 2408 -2468
rect 2472 -4492 2492 -2468
rect 2388 -4788 2492 -4492
rect 199 -4840 2121 -4839
rect 199 -6760 200 -4840
rect 2120 -6760 2121 -4840
rect 199 -6761 2121 -6760
rect -224 -6960 -120 -6812
rect 1108 -6960 1212 -6761
rect 2388 -6812 2408 -4788
rect 2472 -6812 2492 -4788
rect 2388 -6960 2492 -6812
<< properties >>
string FIXED_BBOX 120 4760 2200 6840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10 l 10 val 207.6 carea 2.00 cperi 0.19 nx 2 ny 6 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
