magic
tech sky130A
magscale 1 2
timestamp 1713210209
<< metal3 >>
rect -3546 7146 -1464 8004
rect -1186 7146 896 8000
rect 1580 7146 3672 8000
rect -3546 6746 3672 7146
rect -3546 5924 -1464 6746
rect -2734 5684 -2332 5924
rect -1186 5920 896 6746
rect 1580 5920 3672 6746
rect -3546 4892 -1464 5684
rect -376 5680 26 5920
rect 2416 5680 2818 5920
rect -1186 4892 896 5680
rect 1580 4892 3672 5680
rect -3546 4492 3672 4892
rect -3546 3604 -1464 4492
rect -2734 3364 -2332 3604
rect -1186 3600 896 4492
rect 1580 3600 3672 4492
rect -3546 2546 -1464 3364
rect -376 3360 26 3600
rect 2416 3360 2818 3600
rect -1186 2546 896 3360
rect 1580 2546 3672 3360
rect -3546 2146 3672 2546
rect -3546 1284 -1464 2146
rect -2734 1044 -2332 1284
rect -1186 1280 896 2146
rect 1580 1280 3672 2146
rect -3546 224 -1464 1044
rect -376 1040 26 1280
rect 2416 1040 2818 1280
rect -1186 224 896 1040
rect 1580 224 3672 1040
rect -3546 -176 3672 224
rect -3546 -1036 -1464 -176
rect -2734 -1276 -2332 -1036
rect -1186 -1040 896 -176
rect 1580 -1040 3672 -176
rect -3546 -2160 -1464 -1276
rect -376 -1280 26 -1040
rect 2416 -1280 2818 -1040
rect -1186 -2160 896 -1280
rect 1580 -2160 3672 -1280
rect -3546 -2560 3672 -2160
rect -3546 -3356 -1464 -2560
rect -2734 -3596 -2332 -3356
rect -1186 -3360 896 -2560
rect 1580 -3360 3672 -2560
rect -3546 -4396 -1464 -3596
rect -376 -3600 26 -3360
rect 2416 -3600 2818 -3360
rect -1186 -4396 896 -3600
rect 1580 -4396 3672 -3600
rect -3546 -4796 3672 -4396
rect -3546 -5676 -1464 -4796
rect -2734 -5916 -2332 -5676
rect -1186 -5680 896 -4796
rect 1580 -5680 3672 -4796
rect -3546 -6778 -1464 -5916
rect -376 -5920 26 -5680
rect 2416 -5920 2818 -5680
rect -1186 -6778 896 -5920
rect 1580 -6778 3672 -5920
rect -3546 -7178 3672 -6778
rect -3546 -7996 -1464 -7178
rect -1186 -8000 896 -7178
rect 1580 -8000 3672 -7178
<< mimcap >>
rect -3506 7924 -1506 7964
rect -3506 6004 -3466 7924
rect -1546 6004 -1506 7924
rect -3506 5964 -1506 6004
rect -1146 7920 854 7960
rect -1146 6000 -1106 7920
rect 814 6000 854 7920
rect -1146 5960 854 6000
rect 1620 7920 3620 7960
rect 1620 6000 1660 7920
rect 3580 6000 3620 7920
rect 1620 5960 3620 6000
rect -3506 5604 -1506 5644
rect -3506 3684 -3466 5604
rect -1546 3684 -1506 5604
rect -3506 3644 -1506 3684
rect -1146 5600 854 5640
rect -1146 3680 -1106 5600
rect 814 3680 854 5600
rect -1146 3640 854 3680
rect 1620 5600 3620 5640
rect 1620 3680 1660 5600
rect 3580 3680 3620 5600
rect 1620 3640 3620 3680
rect -3506 3284 -1506 3324
rect -3506 1364 -3466 3284
rect -1546 1364 -1506 3284
rect -3506 1324 -1506 1364
rect -1146 3280 854 3320
rect -1146 1360 -1106 3280
rect 814 1360 854 3280
rect -1146 1320 854 1360
rect 1620 3280 3620 3320
rect 1620 1360 1660 3280
rect 3580 1360 3620 3280
rect 1620 1320 3620 1360
rect -3506 964 -1506 1004
rect -3506 -956 -3466 964
rect -1546 -956 -1506 964
rect -3506 -996 -1506 -956
rect -1146 960 854 1000
rect -1146 -960 -1106 960
rect 814 -960 854 960
rect -1146 -1000 854 -960
rect 1620 960 3620 1000
rect 1620 -960 1660 960
rect 3580 -960 3620 960
rect 1620 -1000 3620 -960
rect -3506 -1356 -1506 -1316
rect -3506 -3276 -3466 -1356
rect -1546 -3276 -1506 -1356
rect -3506 -3316 -1506 -3276
rect -1146 -1360 854 -1320
rect -1146 -3280 -1106 -1360
rect 814 -3280 854 -1360
rect -1146 -3320 854 -3280
rect 1620 -1360 3620 -1320
rect 1620 -3280 1660 -1360
rect 3580 -3280 3620 -1360
rect 1620 -3320 3620 -3280
rect -3506 -3676 -1506 -3636
rect -3506 -5596 -3466 -3676
rect -1546 -5596 -1506 -3676
rect -3506 -5636 -1506 -5596
rect -1146 -3680 854 -3640
rect -1146 -5600 -1106 -3680
rect 814 -5600 854 -3680
rect -1146 -5640 854 -5600
rect 1620 -3680 3620 -3640
rect 1620 -5600 1660 -3680
rect 3580 -5600 3620 -3680
rect 1620 -5640 3620 -5600
rect -3506 -5996 -1506 -5956
rect -3506 -7916 -3466 -5996
rect -1546 -7916 -1506 -5996
rect -3506 -7956 -1506 -7916
rect -1146 -6000 854 -5960
rect -1146 -7920 -1106 -6000
rect 814 -7920 854 -6000
rect -1146 -7960 854 -7920
rect 1620 -6000 3620 -5960
rect 1620 -7920 1660 -6000
rect 3580 -7920 3620 -6000
rect 1620 -7960 3620 -7920
<< mimcapcontact >>
rect -3466 6004 -1546 7924
rect -1106 6000 814 7920
rect 1660 6000 3580 7920
rect -3466 3684 -1546 5604
rect -1106 3680 814 5600
rect 1660 3680 3580 5600
rect -3466 1364 -1546 3284
rect -1106 1360 814 3280
rect 1660 1360 3580 3280
rect -3466 -956 -1546 964
rect -1106 -960 814 960
rect 1660 -960 3580 960
rect -3466 -3276 -1546 -1356
rect -1106 -3280 814 -1360
rect 1660 -3280 3580 -1360
rect -3466 -5596 -1546 -3676
rect -1106 -5600 814 -3680
rect 1660 -5600 3580 -3680
rect -3466 -7916 -1546 -5996
rect -1106 -7920 814 -6000
rect 1660 -7920 3580 -6000
<< metal4 >>
rect -2558 7925 -2454 8020
rect -3467 7924 -1545 7925
rect -3467 6004 -3466 7924
rect -1546 7146 -1545 7924
rect -198 7921 -94 8016
rect 2568 7921 2672 8016
rect -1107 7920 815 7921
rect -1107 7146 -1106 7920
rect -1546 6746 -1106 7146
rect -1546 6004 -1545 6746
rect -3467 6003 -1545 6004
rect -2734 5605 -2332 6003
rect -1107 6000 -1106 6746
rect 814 7146 815 7920
rect 1659 7920 3581 7921
rect 1659 7146 1660 7920
rect 814 6746 1660 7146
rect 814 6000 815 6746
rect -1107 5999 815 6000
rect 1659 6000 1660 6746
rect 3580 6000 3581 7920
rect 1659 5999 3581 6000
rect -3467 5604 -1545 5605
rect -3467 3684 -3466 5604
rect -1546 4892 -1545 5604
rect -376 5601 26 5999
rect 2416 5601 2818 5999
rect -1107 5600 815 5601
rect -1107 4892 -1106 5600
rect -1546 4492 -1106 4892
rect -1546 3684 -1545 4492
rect -3467 3683 -1545 3684
rect -2734 3285 -2332 3683
rect -1107 3680 -1106 4492
rect 814 4892 815 5600
rect 1659 5600 3581 5601
rect 1659 4892 1660 5600
rect 814 4492 1660 4892
rect 814 3680 815 4492
rect -1107 3679 815 3680
rect 1659 3680 1660 4492
rect 3580 3680 3581 5600
rect 1659 3679 3581 3680
rect -3467 3284 -1545 3285
rect -3467 1364 -3466 3284
rect -1546 2546 -1545 3284
rect -376 3281 26 3679
rect 2416 3281 2818 3679
rect -1107 3280 815 3281
rect -1107 2546 -1106 3280
rect -1546 2146 -1106 2546
rect -1546 1364 -1545 2146
rect -3467 1363 -1545 1364
rect -2734 965 -2332 1363
rect -1107 1360 -1106 2146
rect 814 2546 815 3280
rect 1659 3280 3581 3281
rect 1659 2546 1660 3280
rect 814 2146 1660 2546
rect 814 1360 815 2146
rect -1107 1359 815 1360
rect 1659 1360 1660 2146
rect 3580 1360 3581 3280
rect 1659 1359 3581 1360
rect -3467 964 -1545 965
rect -3467 -956 -3466 964
rect -1546 224 -1545 964
rect -376 961 26 1359
rect 2416 961 2818 1359
rect -1107 960 815 961
rect -1107 224 -1106 960
rect -1546 -176 -1106 224
rect -1546 -956 -1545 -176
rect -3467 -957 -1545 -956
rect -2734 -1355 -2332 -957
rect -1107 -960 -1106 -176
rect 814 224 815 960
rect 1659 960 3581 961
rect 1659 224 1660 960
rect 814 -176 1660 224
rect 814 -960 815 -176
rect -1107 -961 815 -960
rect 1659 -960 1660 -176
rect 3580 -960 3581 960
rect 1659 -961 3581 -960
rect -3467 -1356 -1545 -1355
rect -3467 -3276 -3466 -1356
rect -1546 -2160 -1545 -1356
rect -376 -1359 26 -961
rect 2416 -1359 2818 -961
rect -1107 -1360 815 -1359
rect -1107 -2160 -1106 -1360
rect -1546 -2560 -1106 -2160
rect -1546 -3276 -1545 -2560
rect -3467 -3277 -1545 -3276
rect -2734 -3675 -2332 -3277
rect -1107 -3280 -1106 -2560
rect 814 -2160 815 -1360
rect 1659 -1360 3581 -1359
rect 1659 -2160 1660 -1360
rect 814 -2560 1660 -2160
rect 814 -3280 815 -2560
rect -1107 -3281 815 -3280
rect 1659 -3280 1660 -2560
rect 3580 -3280 3581 -1360
rect 1659 -3281 3581 -3280
rect -3467 -3676 -1545 -3675
rect -3467 -5596 -3466 -3676
rect -1546 -4396 -1545 -3676
rect -376 -3679 26 -3281
rect 2416 -3679 2818 -3281
rect -1107 -3680 815 -3679
rect -1107 -4396 -1106 -3680
rect -1546 -4796 -1106 -4396
rect -1546 -5596 -1545 -4796
rect -3467 -5597 -1545 -5596
rect -2734 -5995 -2332 -5597
rect -1107 -5600 -1106 -4796
rect 814 -4396 815 -3680
rect 1659 -3680 3581 -3679
rect 1659 -4396 1660 -3680
rect 814 -4796 1660 -4396
rect 814 -5600 815 -4796
rect -1107 -5601 815 -5600
rect 1659 -5600 1660 -4796
rect 3580 -5600 3581 -3680
rect 1659 -5601 3581 -5600
rect -3467 -5996 -1545 -5995
rect -3467 -7916 -3466 -5996
rect -1546 -6778 -1545 -5996
rect -376 -5999 26 -5601
rect 2416 -5999 2818 -5601
rect -1107 -6000 815 -5999
rect -1107 -6778 -1106 -6000
rect -1546 -7178 -1106 -6778
rect -1546 -7916 -1545 -7178
rect -3467 -7917 -1545 -7916
rect -2558 -8004 -2454 -7917
rect -1107 -7920 -1106 -7178
rect 814 -6778 815 -6000
rect 1659 -6000 3581 -5999
rect 1659 -6778 1660 -6000
rect 814 -7178 1660 -6778
rect 814 -7920 815 -7178
rect -1107 -7921 815 -7920
rect 1659 -7920 1660 -7178
rect 3580 -7920 3581 -6000
rect 1659 -7921 3581 -7920
rect -198 -8008 -94 -7921
rect 2568 -8008 2672 -7921
<< properties >>
string FIXED_BBOX 1426 5920 3506 8000
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 3 ny 7 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
