magic
tech sky130A
magscale 1 2
timestamp 1712782684
<< nwell >>
rect -1374 -1161 1374 1161
<< mvpmos >>
rect -1116 64 -716 864
rect -658 64 -258 864
rect -200 64 200 864
rect 258 64 658 864
rect 716 64 1116 864
rect -1116 -864 -716 -64
rect -658 -864 -258 -64
rect -200 -864 200 -64
rect 258 -864 658 -64
rect 716 -864 1116 -64
<< mvpdiff >>
rect -1174 852 -1116 864
rect -1174 76 -1162 852
rect -1128 76 -1116 852
rect -1174 64 -1116 76
rect -716 852 -658 864
rect -716 76 -704 852
rect -670 76 -658 852
rect -716 64 -658 76
rect -258 852 -200 864
rect -258 76 -246 852
rect -212 76 -200 852
rect -258 64 -200 76
rect 200 852 258 864
rect 200 76 212 852
rect 246 76 258 852
rect 200 64 258 76
rect 658 852 716 864
rect 658 76 670 852
rect 704 76 716 852
rect 658 64 716 76
rect 1116 852 1174 864
rect 1116 76 1128 852
rect 1162 76 1174 852
rect 1116 64 1174 76
rect -1174 -76 -1116 -64
rect -1174 -852 -1162 -76
rect -1128 -852 -1116 -76
rect -1174 -864 -1116 -852
rect -716 -76 -658 -64
rect -716 -852 -704 -76
rect -670 -852 -658 -76
rect -716 -864 -658 -852
rect -258 -76 -200 -64
rect -258 -852 -246 -76
rect -212 -852 -200 -76
rect -258 -864 -200 -852
rect 200 -76 258 -64
rect 200 -852 212 -76
rect 246 -852 258 -76
rect 200 -864 258 -852
rect 658 -76 716 -64
rect 658 -852 670 -76
rect 704 -852 716 -76
rect 658 -864 716 -852
rect 1116 -76 1174 -64
rect 1116 -852 1128 -76
rect 1162 -852 1174 -76
rect 1116 -864 1174 -852
<< mvpdiffc >>
rect -1162 76 -1128 852
rect -704 76 -670 852
rect -246 76 -212 852
rect 212 76 246 852
rect 670 76 704 852
rect 1128 76 1162 852
rect -1162 -852 -1128 -76
rect -704 -852 -670 -76
rect -246 -852 -212 -76
rect 212 -852 246 -76
rect 670 -852 704 -76
rect 1128 -852 1162 -76
<< mvnsubdiff >>
rect -1308 1083 1308 1095
rect -1308 1049 -1200 1083
rect 1200 1049 1308 1083
rect -1308 1037 1308 1049
rect -1308 987 -1250 1037
rect -1308 -987 -1296 987
rect -1262 -987 -1250 987
rect 1250 987 1308 1037
rect -1308 -1037 -1250 -987
rect 1250 -987 1262 987
rect 1296 -987 1308 987
rect 1250 -1037 1308 -987
rect -1308 -1049 1308 -1037
rect -1308 -1083 -1200 -1049
rect 1200 -1083 1308 -1049
rect -1308 -1095 1308 -1083
<< mvnsubdiffcont >>
rect -1200 1049 1200 1083
rect -1296 -987 -1262 987
rect 1262 -987 1296 987
rect -1200 -1083 1200 -1049
<< poly >>
rect -1116 945 -716 961
rect -1116 911 -1100 945
rect -732 911 -716 945
rect -1116 864 -716 911
rect -658 945 -258 961
rect -658 911 -642 945
rect -274 911 -258 945
rect -658 864 -258 911
rect -200 945 200 961
rect -200 911 -184 945
rect 184 911 200 945
rect -200 864 200 911
rect 258 945 658 961
rect 258 911 274 945
rect 642 911 658 945
rect 258 864 658 911
rect 716 945 1116 961
rect 716 911 732 945
rect 1100 911 1116 945
rect 716 864 1116 911
rect -1116 17 -716 64
rect -1116 -17 -1100 17
rect -732 -17 -716 17
rect -1116 -64 -716 -17
rect -658 17 -258 64
rect -658 -17 -642 17
rect -274 -17 -258 17
rect -658 -64 -258 -17
rect -200 17 200 64
rect -200 -17 -184 17
rect 184 -17 200 17
rect -200 -64 200 -17
rect 258 17 658 64
rect 258 -17 274 17
rect 642 -17 658 17
rect 258 -64 658 -17
rect 716 17 1116 64
rect 716 -17 732 17
rect 1100 -17 1116 17
rect 716 -64 1116 -17
rect -1116 -911 -716 -864
rect -1116 -945 -1100 -911
rect -732 -945 -716 -911
rect -1116 -961 -716 -945
rect -658 -911 -258 -864
rect -658 -945 -642 -911
rect -274 -945 -258 -911
rect -658 -961 -258 -945
rect -200 -911 200 -864
rect -200 -945 -184 -911
rect 184 -945 200 -911
rect -200 -961 200 -945
rect 258 -911 658 -864
rect 258 -945 274 -911
rect 642 -945 658 -911
rect 258 -961 658 -945
rect 716 -911 1116 -864
rect 716 -945 732 -911
rect 1100 -945 1116 -911
rect 716 -961 1116 -945
<< polycont >>
rect -1100 911 -732 945
rect -642 911 -274 945
rect -184 911 184 945
rect 274 911 642 945
rect 732 911 1100 945
rect -1100 -17 -732 17
rect -642 -17 -274 17
rect -184 -17 184 17
rect 274 -17 642 17
rect 732 -17 1100 17
rect -1100 -945 -732 -911
rect -642 -945 -274 -911
rect -184 -945 184 -911
rect 274 -945 642 -911
rect 732 -945 1100 -911
<< locali >>
rect -1296 1049 -1200 1083
rect 1200 1049 1296 1083
rect -1296 987 -1262 1049
rect 1262 987 1296 1049
rect -1116 911 -1100 945
rect -732 911 -716 945
rect -658 911 -642 945
rect -274 911 -258 945
rect -200 911 -184 945
rect 184 911 200 945
rect 258 911 274 945
rect 642 911 658 945
rect 716 911 732 945
rect 1100 911 1116 945
rect -1162 852 -1128 868
rect -1162 60 -1128 76
rect -704 852 -670 868
rect -704 60 -670 76
rect -246 852 -212 868
rect -246 60 -212 76
rect 212 852 246 868
rect 212 60 246 76
rect 670 852 704 868
rect 670 60 704 76
rect 1128 852 1162 868
rect 1128 60 1162 76
rect -1116 -17 -1100 17
rect -732 -17 -716 17
rect -658 -17 -642 17
rect -274 -17 -258 17
rect -200 -17 -184 17
rect 184 -17 200 17
rect 258 -17 274 17
rect 642 -17 658 17
rect 716 -17 732 17
rect 1100 -17 1116 17
rect -1162 -76 -1128 -60
rect -1162 -868 -1128 -852
rect -704 -76 -670 -60
rect -704 -868 -670 -852
rect -246 -76 -212 -60
rect -246 -868 -212 -852
rect 212 -76 246 -60
rect 212 -868 246 -852
rect 670 -76 704 -60
rect 670 -868 704 -852
rect 1128 -76 1162 -60
rect 1128 -868 1162 -852
rect -1116 -945 -1100 -911
rect -732 -945 -716 -911
rect -658 -945 -642 -911
rect -274 -945 -258 -911
rect -200 -945 -184 -911
rect 184 -945 200 -911
rect 258 -945 274 -911
rect 642 -945 658 -911
rect 716 -945 732 -911
rect 1100 -945 1116 -911
rect -1296 -1049 -1262 -987
rect 1262 -1049 1296 -987
rect -1296 -1083 -1200 -1049
rect 1200 -1083 1296 -1049
<< viali >>
rect -1100 911 -732 945
rect -642 911 -274 945
rect -184 911 184 945
rect 274 911 642 945
rect 732 911 1100 945
rect -1162 76 -1128 852
rect -704 76 -670 852
rect -246 76 -212 852
rect 212 76 246 852
rect 670 76 704 852
rect 1128 76 1162 852
rect -1100 -17 -732 17
rect -642 -17 -274 17
rect -184 -17 184 17
rect 274 -17 642 17
rect 732 -17 1100 17
rect -1162 -852 -1128 -76
rect -704 -852 -670 -76
rect -246 -852 -212 -76
rect 212 -852 246 -76
rect 670 -852 704 -76
rect 1128 -852 1162 -76
rect -1100 -945 -732 -911
rect -642 -945 -274 -911
rect -184 -945 184 -911
rect 274 -945 642 -911
rect 732 -945 1100 -911
<< metal1 >>
rect -1112 945 -720 951
rect -1112 911 -1100 945
rect -732 911 -720 945
rect -1112 905 -720 911
rect -654 945 -262 951
rect -654 911 -642 945
rect -274 911 -262 945
rect -654 905 -262 911
rect -196 945 196 951
rect -196 911 -184 945
rect 184 911 196 945
rect -196 905 196 911
rect 262 945 654 951
rect 262 911 274 945
rect 642 911 654 945
rect 262 905 654 911
rect 720 945 1112 951
rect 720 911 732 945
rect 1100 911 1112 945
rect 720 905 1112 911
rect -1168 852 -1122 864
rect -1168 76 -1162 852
rect -1128 76 -1122 852
rect -1168 64 -1122 76
rect -710 852 -664 864
rect -710 76 -704 852
rect -670 76 -664 852
rect -710 64 -664 76
rect -252 852 -206 864
rect -252 76 -246 852
rect -212 76 -206 852
rect -252 64 -206 76
rect 206 852 252 864
rect 206 76 212 852
rect 246 76 252 852
rect 206 64 252 76
rect 664 852 710 864
rect 664 76 670 852
rect 704 76 710 852
rect 664 64 710 76
rect 1122 852 1168 864
rect 1122 76 1128 852
rect 1162 76 1168 852
rect 1122 64 1168 76
rect -1112 17 -720 23
rect -1112 -17 -1100 17
rect -732 -17 -720 17
rect -1112 -23 -720 -17
rect -654 17 -262 23
rect -654 -17 -642 17
rect -274 -17 -262 17
rect -654 -23 -262 -17
rect -196 17 196 23
rect -196 -17 -184 17
rect 184 -17 196 17
rect -196 -23 196 -17
rect 262 17 654 23
rect 262 -17 274 17
rect 642 -17 654 17
rect 262 -23 654 -17
rect 720 17 1112 23
rect 720 -17 732 17
rect 1100 -17 1112 17
rect 720 -23 1112 -17
rect -1168 -76 -1122 -64
rect -1168 -852 -1162 -76
rect -1128 -852 -1122 -76
rect -1168 -864 -1122 -852
rect -710 -76 -664 -64
rect -710 -852 -704 -76
rect -670 -852 -664 -76
rect -710 -864 -664 -852
rect -252 -76 -206 -64
rect -252 -852 -246 -76
rect -212 -852 -206 -76
rect -252 -864 -206 -852
rect 206 -76 252 -64
rect 206 -852 212 -76
rect 246 -852 252 -76
rect 206 -864 252 -852
rect 664 -76 710 -64
rect 664 -852 670 -76
rect 704 -852 710 -76
rect 664 -864 710 -852
rect 1122 -76 1168 -64
rect 1122 -852 1128 -76
rect 1162 -852 1168 -76
rect 1122 -864 1168 -852
rect -1112 -911 -720 -905
rect -1112 -945 -1100 -911
rect -732 -945 -720 -911
rect -1112 -951 -720 -945
rect -654 -911 -262 -905
rect -654 -945 -642 -911
rect -274 -945 -262 -911
rect -654 -951 -262 -945
rect -196 -911 196 -905
rect -196 -945 -184 -911
rect 184 -945 196 -911
rect -196 -951 196 -945
rect 262 -911 654 -905
rect 262 -945 274 -911
rect 642 -945 654 -911
rect 262 -951 654 -945
rect 720 -911 1112 -905
rect 720 -945 732 -911
rect 1100 -945 1112 -911
rect 720 -951 1112 -945
<< properties >>
string FIXED_BBOX -1279 -1066 1279 1066
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 2.0 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
