magic
tech sky130A
magscale 1 2
timestamp 1713017924
<< metal3 >>
rect -2492 2172 -120 2200
rect -2492 148 -204 2172
rect -140 148 -120 2172
rect -2492 120 -120 148
rect 120 2172 2492 2200
rect 120 148 2408 2172
rect 2472 148 2492 2172
rect 120 120 2492 148
rect -2492 -148 -120 -120
rect -2492 -2172 -204 -148
rect -140 -2172 -120 -148
rect -2492 -2200 -120 -2172
rect 120 -148 2492 -120
rect 120 -2172 2408 -148
rect 2472 -2172 2492 -148
rect 120 -2200 2492 -2172
<< via3 >>
rect -204 148 -140 2172
rect 2408 148 2472 2172
rect -204 -2172 -140 -148
rect 2408 -2172 2472 -148
<< mimcap >>
rect -2452 2120 -452 2160
rect -2452 200 -2412 2120
rect -492 200 -452 2120
rect -2452 160 -452 200
rect 160 2120 2160 2160
rect 160 200 200 2120
rect 2120 200 2160 2120
rect 160 160 2160 200
rect -2452 -200 -452 -160
rect -2452 -2120 -2412 -200
rect -492 -2120 -452 -200
rect -2452 -2160 -452 -2120
rect 160 -200 2160 -160
rect 160 -2120 200 -200
rect 2120 -2120 2160 -200
rect 160 -2160 2160 -2120
<< mimcapcontact >>
rect -2412 200 -492 2120
rect 200 200 2120 2120
rect -2412 -2120 -492 -200
rect 200 -2120 2120 -200
<< metal4 >>
rect -1504 2121 -1400 2320
rect -224 2172 -120 2320
rect -2413 2120 -491 2121
rect -2413 200 -2412 2120
rect -492 200 -491 2120
rect -2413 199 -491 200
rect -1504 -199 -1400 199
rect -224 148 -204 2172
rect -140 148 -120 2172
rect 1108 2121 1212 2320
rect 2388 2172 2492 2320
rect 199 2120 2121 2121
rect 199 200 200 2120
rect 2120 200 2121 2120
rect 199 199 2121 200
rect -224 -148 -120 148
rect -2413 -200 -491 -199
rect -2413 -2120 -2412 -200
rect -492 -2120 -491 -200
rect -2413 -2121 -491 -2120
rect -1504 -2320 -1400 -2121
rect -224 -2172 -204 -148
rect -140 -2172 -120 -148
rect 1108 -199 1212 199
rect 2388 148 2408 2172
rect 2472 148 2492 2172
rect 2388 -148 2492 148
rect 199 -200 2121 -199
rect 199 -2120 200 -200
rect 2120 -2120 2121 -200
rect 199 -2121 2121 -2120
rect -224 -2320 -120 -2172
rect 1108 -2320 1212 -2121
rect 2388 -2172 2408 -148
rect 2472 -2172 2492 -148
rect 2388 -2320 2492 -2172
<< properties >>
string FIXED_BBOX 120 120 2200 2200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
