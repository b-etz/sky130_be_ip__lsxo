magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< nwell >>
rect -396 -2691 396 2691
<< pmos >>
rect -200 1672 200 2472
rect -200 636 200 1436
rect -200 -400 200 400
rect -200 -1436 200 -636
rect -200 -2472 200 -1672
<< pdiff >>
rect -258 2460 -200 2472
rect -258 1684 -246 2460
rect -212 1684 -200 2460
rect -258 1672 -200 1684
rect 200 2460 258 2472
rect 200 1684 212 2460
rect 246 1684 258 2460
rect 200 1672 258 1684
rect -258 1424 -200 1436
rect -258 648 -246 1424
rect -212 648 -200 1424
rect -258 636 -200 648
rect 200 1424 258 1436
rect 200 648 212 1424
rect 246 648 258 1424
rect 200 636 258 648
rect -258 388 -200 400
rect -258 -388 -246 388
rect -212 -388 -200 388
rect -258 -400 -200 -388
rect 200 388 258 400
rect 200 -388 212 388
rect 246 -388 258 388
rect 200 -400 258 -388
rect -258 -648 -200 -636
rect -258 -1424 -246 -648
rect -212 -1424 -200 -648
rect -258 -1436 -200 -1424
rect 200 -648 258 -636
rect 200 -1424 212 -648
rect 246 -1424 258 -648
rect 200 -1436 258 -1424
rect -258 -1684 -200 -1672
rect -258 -2460 -246 -1684
rect -212 -2460 -200 -1684
rect -258 -2472 -200 -2460
rect 200 -1684 258 -1672
rect 200 -2460 212 -1684
rect 246 -2460 258 -1684
rect 200 -2472 258 -2460
<< pdiffc >>
rect -246 1684 -212 2460
rect 212 1684 246 2460
rect -246 648 -212 1424
rect 212 648 246 1424
rect -246 -388 -212 388
rect 212 -388 246 388
rect -246 -1424 -212 -648
rect 212 -1424 246 -648
rect -246 -2460 -212 -1684
rect 212 -2460 246 -1684
<< nsubdiff >>
rect -360 2621 -264 2655
rect 264 2621 360 2655
rect -360 2559 -326 2621
rect 326 2559 360 2621
rect -360 -2621 -326 -2559
rect 326 -2621 360 -2559
rect -360 -2655 -264 -2621
rect 264 -2655 360 -2621
<< nsubdiffcont >>
rect -264 2621 264 2655
rect -360 -2559 -326 2559
rect 326 -2559 360 2559
rect -264 -2655 264 -2621
<< poly >>
rect -200 2553 200 2569
rect -200 2519 -184 2553
rect 184 2519 200 2553
rect -200 2472 200 2519
rect -200 1625 200 1672
rect -200 1591 -184 1625
rect 184 1591 200 1625
rect -200 1575 200 1591
rect -200 1517 200 1533
rect -200 1483 -184 1517
rect 184 1483 200 1517
rect -200 1436 200 1483
rect -200 589 200 636
rect -200 555 -184 589
rect 184 555 200 589
rect -200 539 200 555
rect -200 481 200 497
rect -200 447 -184 481
rect 184 447 200 481
rect -200 400 200 447
rect -200 -447 200 -400
rect -200 -481 -184 -447
rect 184 -481 200 -447
rect -200 -497 200 -481
rect -200 -555 200 -539
rect -200 -589 -184 -555
rect 184 -589 200 -555
rect -200 -636 200 -589
rect -200 -1483 200 -1436
rect -200 -1517 -184 -1483
rect 184 -1517 200 -1483
rect -200 -1533 200 -1517
rect -200 -1591 200 -1575
rect -200 -1625 -184 -1591
rect 184 -1625 200 -1591
rect -200 -1672 200 -1625
rect -200 -2519 200 -2472
rect -200 -2553 -184 -2519
rect 184 -2553 200 -2519
rect -200 -2569 200 -2553
<< polycont >>
rect -184 2519 184 2553
rect -184 1591 184 1625
rect -184 1483 184 1517
rect -184 555 184 589
rect -184 447 184 481
rect -184 -481 184 -447
rect -184 -589 184 -555
rect -184 -1517 184 -1483
rect -184 -1625 184 -1591
rect -184 -2553 184 -2519
<< locali >>
rect -360 2621 -264 2655
rect 264 2621 360 2655
rect -360 2559 -326 2621
rect 326 2559 360 2621
rect -200 2519 -184 2553
rect 184 2519 200 2553
rect -246 2460 -212 2476
rect -246 1668 -212 1684
rect 212 2460 246 2476
rect 212 1668 246 1684
rect -200 1591 -184 1625
rect 184 1591 200 1625
rect -200 1483 -184 1517
rect 184 1483 200 1517
rect -246 1424 -212 1440
rect -246 632 -212 648
rect 212 1424 246 1440
rect 212 632 246 648
rect -200 555 -184 589
rect 184 555 200 589
rect -200 447 -184 481
rect 184 447 200 481
rect -246 388 -212 404
rect -246 -404 -212 -388
rect 212 388 246 404
rect 212 -404 246 -388
rect -200 -481 -184 -447
rect 184 -481 200 -447
rect -200 -589 -184 -555
rect 184 -589 200 -555
rect -246 -648 -212 -632
rect -246 -1440 -212 -1424
rect 212 -648 246 -632
rect 212 -1440 246 -1424
rect -200 -1517 -184 -1483
rect 184 -1517 200 -1483
rect -200 -1625 -184 -1591
rect 184 -1625 200 -1591
rect -246 -1684 -212 -1668
rect -246 -2476 -212 -2460
rect 212 -1684 246 -1668
rect 212 -2476 246 -2460
rect -200 -2553 -184 -2519
rect 184 -2553 200 -2519
rect -360 -2621 -326 -2559
rect 326 -2621 360 -2559
rect -360 -2655 -264 -2621
rect 264 -2655 360 -2621
<< viali >>
rect -184 2519 184 2553
rect -246 1684 -212 2460
rect 212 1684 246 2460
rect -184 1591 184 1625
rect -184 1483 184 1517
rect -246 648 -212 1424
rect 212 648 246 1424
rect -184 555 184 589
rect -184 447 184 481
rect -246 -388 -212 388
rect 212 -388 246 388
rect -184 -481 184 -447
rect -184 -589 184 -555
rect -246 -1424 -212 -648
rect 212 -1424 246 -648
rect -184 -1517 184 -1483
rect -184 -1625 184 -1591
rect -246 -2460 -212 -1684
rect 212 -2460 246 -1684
rect -184 -2553 184 -2519
<< metal1 >>
rect -196 2553 196 2559
rect -196 2519 -184 2553
rect 184 2519 196 2553
rect -196 2513 196 2519
rect -252 2460 -206 2472
rect -252 1684 -246 2460
rect -212 1684 -206 2460
rect -252 1672 -206 1684
rect 206 2460 252 2472
rect 206 1684 212 2460
rect 246 1684 252 2460
rect 206 1672 252 1684
rect -196 1625 196 1631
rect -196 1591 -184 1625
rect 184 1591 196 1625
rect -196 1585 196 1591
rect -196 1517 196 1523
rect -196 1483 -184 1517
rect 184 1483 196 1517
rect -196 1477 196 1483
rect -252 1424 -206 1436
rect -252 648 -246 1424
rect -212 648 -206 1424
rect -252 636 -206 648
rect 206 1424 252 1436
rect 206 648 212 1424
rect 246 648 252 1424
rect 206 636 252 648
rect -196 589 196 595
rect -196 555 -184 589
rect 184 555 196 589
rect -196 549 196 555
rect -196 481 196 487
rect -196 447 -184 481
rect 184 447 196 481
rect -196 441 196 447
rect -252 388 -206 400
rect -252 -388 -246 388
rect -212 -388 -206 388
rect -252 -400 -206 -388
rect 206 388 252 400
rect 206 -388 212 388
rect 246 -388 252 388
rect 206 -400 252 -388
rect -196 -447 196 -441
rect -196 -481 -184 -447
rect 184 -481 196 -447
rect -196 -487 196 -481
rect -196 -555 196 -549
rect -196 -589 -184 -555
rect 184 -589 196 -555
rect -196 -595 196 -589
rect -252 -648 -206 -636
rect -252 -1424 -246 -648
rect -212 -1424 -206 -648
rect -252 -1436 -206 -1424
rect 206 -648 252 -636
rect 206 -1424 212 -648
rect 246 -1424 252 -648
rect 206 -1436 252 -1424
rect -196 -1483 196 -1477
rect -196 -1517 -184 -1483
rect 184 -1517 196 -1483
rect -196 -1523 196 -1517
rect -196 -1591 196 -1585
rect -196 -1625 -184 -1591
rect 184 -1625 196 -1591
rect -196 -1631 196 -1625
rect -252 -1684 -206 -1672
rect -252 -2460 -246 -1684
rect -212 -2460 -206 -1684
rect -252 -2472 -206 -2460
rect 206 -1684 252 -1672
rect 206 -2460 212 -1684
rect 246 -2460 252 -1684
rect 206 -2472 252 -2460
rect -196 -2519 196 -2513
rect -196 -2553 -184 -2519
rect 184 -2553 196 -2519
rect -196 -2559 196 -2553
<< properties >>
string FIXED_BBOX -343 -2638 343 2638
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.0 l 2.0 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
