magic
tech sky130A
timestamp 1712071977
<< pwell >>
rect -214 -847 214 847
<< mvnmos >>
rect -100 518 100 718
rect -100 209 100 409
rect -100 -100 100 100
rect -100 -409 100 -209
rect -100 -718 100 -518
<< mvndiff >>
rect -129 712 -100 718
rect -129 524 -123 712
rect -106 524 -100 712
rect -129 518 -100 524
rect 100 712 129 718
rect 100 524 106 712
rect 123 524 129 712
rect 100 518 129 524
rect -129 403 -100 409
rect -129 215 -123 403
rect -106 215 -100 403
rect -129 209 -100 215
rect 100 403 129 409
rect 100 215 106 403
rect 123 215 129 403
rect 100 209 129 215
rect -129 94 -100 100
rect -129 -94 -123 94
rect -106 -94 -100 94
rect -129 -100 -100 -94
rect 100 94 129 100
rect 100 -94 106 94
rect 123 -94 129 94
rect 100 -100 129 -94
rect -129 -215 -100 -209
rect -129 -403 -123 -215
rect -106 -403 -100 -215
rect -129 -409 -100 -403
rect 100 -215 129 -209
rect 100 -403 106 -215
rect 123 -403 129 -215
rect 100 -409 129 -403
rect -129 -524 -100 -518
rect -129 -712 -123 -524
rect -106 -712 -100 -524
rect -129 -718 -100 -712
rect 100 -524 129 -518
rect 100 -712 106 -524
rect 123 -712 129 -524
rect 100 -718 129 -712
<< mvndiffc >>
rect -123 524 -106 712
rect 106 524 123 712
rect -123 215 -106 403
rect 106 215 123 403
rect -123 -94 -106 94
rect 106 -94 123 94
rect -123 -403 -106 -215
rect 106 -403 123 -215
rect -123 -712 -106 -524
rect 106 -712 123 -524
<< mvpsubdiff >>
rect -196 823 196 829
rect -196 806 -142 823
rect 142 806 196 823
rect -196 800 196 806
rect -196 775 -167 800
rect -196 -775 -190 775
rect -173 -775 -167 775
rect 167 775 196 800
rect -196 -800 -167 -775
rect 167 -775 173 775
rect 190 -775 196 775
rect 167 -800 196 -775
rect -196 -806 196 -800
rect -196 -823 -142 -806
rect 142 -823 196 -806
rect -196 -829 196 -823
<< mvpsubdiffcont >>
rect -142 806 142 823
rect -190 -775 -173 775
rect 173 -775 190 775
rect -142 -823 142 -806
<< poly >>
rect -100 754 100 762
rect -100 737 -92 754
rect 92 737 100 754
rect -100 718 100 737
rect -100 499 100 518
rect -100 482 -92 499
rect 92 482 100 499
rect -100 474 100 482
rect -100 445 100 453
rect -100 428 -92 445
rect 92 428 100 445
rect -100 409 100 428
rect -100 190 100 209
rect -100 173 -92 190
rect 92 173 100 190
rect -100 165 100 173
rect -100 136 100 144
rect -100 119 -92 136
rect 92 119 100 136
rect -100 100 100 119
rect -100 -119 100 -100
rect -100 -136 -92 -119
rect 92 -136 100 -119
rect -100 -144 100 -136
rect -100 -173 100 -165
rect -100 -190 -92 -173
rect 92 -190 100 -173
rect -100 -209 100 -190
rect -100 -428 100 -409
rect -100 -445 -92 -428
rect 92 -445 100 -428
rect -100 -453 100 -445
rect -100 -482 100 -474
rect -100 -499 -92 -482
rect 92 -499 100 -482
rect -100 -518 100 -499
rect -100 -737 100 -718
rect -100 -754 -92 -737
rect 92 -754 100 -737
rect -100 -762 100 -754
<< polycont >>
rect -92 737 92 754
rect -92 482 92 499
rect -92 428 92 445
rect -92 173 92 190
rect -92 119 92 136
rect -92 -136 92 -119
rect -92 -190 92 -173
rect -92 -445 92 -428
rect -92 -499 92 -482
rect -92 -754 92 -737
<< locali >>
rect -190 806 -142 823
rect 142 806 190 823
rect -190 775 -173 806
rect 173 775 190 806
rect -100 737 -92 754
rect 92 737 100 754
rect -123 712 -106 720
rect -123 516 -106 524
rect 106 712 123 720
rect 106 516 123 524
rect -100 482 -92 499
rect 92 482 100 499
rect -100 428 -92 445
rect 92 428 100 445
rect -123 403 -106 411
rect -123 207 -106 215
rect 106 403 123 411
rect 106 207 123 215
rect -100 173 -92 190
rect 92 173 100 190
rect -100 119 -92 136
rect 92 119 100 136
rect -123 94 -106 102
rect -123 -102 -106 -94
rect 106 94 123 102
rect 106 -102 123 -94
rect -100 -136 -92 -119
rect 92 -136 100 -119
rect -100 -190 -92 -173
rect 92 -190 100 -173
rect -123 -215 -106 -207
rect -123 -411 -106 -403
rect 106 -215 123 -207
rect 106 -411 123 -403
rect -100 -445 -92 -428
rect 92 -445 100 -428
rect -100 -499 -92 -482
rect 92 -499 100 -482
rect -123 -524 -106 -516
rect -123 -720 -106 -712
rect 106 -524 123 -516
rect 106 -720 123 -712
rect -100 -754 -92 -737
rect 92 -754 100 -737
rect -190 -806 -173 -775
rect 173 -806 190 -775
rect -190 -823 -142 -806
rect 142 -823 190 -806
<< viali >>
rect -92 737 92 754
rect -123 524 -106 712
rect 106 524 123 712
rect -92 482 92 499
rect -92 428 92 445
rect -123 215 -106 403
rect 106 215 123 403
rect -92 173 92 190
rect -92 119 92 136
rect -123 -94 -106 94
rect 106 -94 123 94
rect -92 -136 92 -119
rect -92 -190 92 -173
rect -123 -403 -106 -215
rect 106 -403 123 -215
rect -92 -445 92 -428
rect -92 -499 92 -482
rect -123 -712 -106 -524
rect 106 -712 123 -524
rect -92 -754 92 -737
<< metal1 >>
rect -98 754 98 757
rect -98 737 -92 754
rect 92 737 98 754
rect -98 734 98 737
rect -126 712 -103 718
rect -126 524 -123 712
rect -106 524 -103 712
rect -126 518 -103 524
rect 103 712 126 718
rect 103 524 106 712
rect 123 524 126 712
rect 103 518 126 524
rect -98 499 98 502
rect -98 482 -92 499
rect 92 482 98 499
rect -98 479 98 482
rect -98 445 98 448
rect -98 428 -92 445
rect 92 428 98 445
rect -98 425 98 428
rect -126 403 -103 409
rect -126 215 -123 403
rect -106 215 -103 403
rect -126 209 -103 215
rect 103 403 126 409
rect 103 215 106 403
rect 123 215 126 403
rect 103 209 126 215
rect -98 190 98 193
rect -98 173 -92 190
rect 92 173 98 190
rect -98 170 98 173
rect -98 136 98 139
rect -98 119 -92 136
rect 92 119 98 136
rect -98 116 98 119
rect -126 94 -103 100
rect -126 -94 -123 94
rect -106 -94 -103 94
rect -126 -100 -103 -94
rect 103 94 126 100
rect 103 -94 106 94
rect 123 -94 126 94
rect 103 -100 126 -94
rect -98 -119 98 -116
rect -98 -136 -92 -119
rect 92 -136 98 -119
rect -98 -139 98 -136
rect -98 -173 98 -170
rect -98 -190 -92 -173
rect 92 -190 98 -173
rect -98 -193 98 -190
rect -126 -215 -103 -209
rect -126 -403 -123 -215
rect -106 -403 -103 -215
rect -126 -409 -103 -403
rect 103 -215 126 -209
rect 103 -403 106 -215
rect 123 -403 126 -215
rect 103 -409 126 -403
rect -98 -428 98 -425
rect -98 -445 -92 -428
rect 92 -445 98 -428
rect -98 -448 98 -445
rect -98 -482 98 -479
rect -98 -499 -92 -482
rect 92 -499 98 -482
rect -98 -502 98 -499
rect -126 -524 -103 -518
rect -126 -712 -123 -524
rect -106 -712 -103 -524
rect -126 -718 -103 -712
rect 103 -524 126 -518
rect 103 -712 106 -524
rect 123 -712 126 -524
rect 103 -718 126 -712
rect -98 -737 98 -734
rect -98 -754 -92 -737
rect 92 -754 98 -737
rect -98 -757 98 -754
<< properties >>
string FIXED_BBOX -181 -814 181 814
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.0 l 2.0 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
