magic
tech sky130A
magscale 1 2
timestamp 1712965163
<< nwell >>
rect -2061 -1161 2061 1161
<< mvpmos >>
rect -1803 64 -1403 864
rect -1345 64 -945 864
rect -887 64 -487 864
rect -429 64 -29 864
rect 29 64 429 864
rect 487 64 887 864
rect 945 64 1345 864
rect 1403 64 1803 864
rect -1803 -864 -1403 -64
rect -1345 -864 -945 -64
rect -887 -864 -487 -64
rect -429 -864 -29 -64
rect 29 -864 429 -64
rect 487 -864 887 -64
rect 945 -864 1345 -64
rect 1403 -864 1803 -64
<< mvpdiff >>
rect -1861 852 -1803 864
rect -1861 76 -1849 852
rect -1815 76 -1803 852
rect -1861 64 -1803 76
rect -1403 852 -1345 864
rect -1403 76 -1391 852
rect -1357 76 -1345 852
rect -1403 64 -1345 76
rect -945 852 -887 864
rect -945 76 -933 852
rect -899 76 -887 852
rect -945 64 -887 76
rect -487 852 -429 864
rect -487 76 -475 852
rect -441 76 -429 852
rect -487 64 -429 76
rect -29 852 29 864
rect -29 76 -17 852
rect 17 76 29 852
rect -29 64 29 76
rect 429 852 487 864
rect 429 76 441 852
rect 475 76 487 852
rect 429 64 487 76
rect 887 852 945 864
rect 887 76 899 852
rect 933 76 945 852
rect 887 64 945 76
rect 1345 852 1403 864
rect 1345 76 1357 852
rect 1391 76 1403 852
rect 1345 64 1403 76
rect 1803 852 1861 864
rect 1803 76 1815 852
rect 1849 76 1861 852
rect 1803 64 1861 76
rect -1861 -76 -1803 -64
rect -1861 -852 -1849 -76
rect -1815 -852 -1803 -76
rect -1861 -864 -1803 -852
rect -1403 -76 -1345 -64
rect -1403 -852 -1391 -76
rect -1357 -852 -1345 -76
rect -1403 -864 -1345 -852
rect -945 -76 -887 -64
rect -945 -852 -933 -76
rect -899 -852 -887 -76
rect -945 -864 -887 -852
rect -487 -76 -429 -64
rect -487 -852 -475 -76
rect -441 -852 -429 -76
rect -487 -864 -429 -852
rect -29 -76 29 -64
rect -29 -852 -17 -76
rect 17 -852 29 -76
rect -29 -864 29 -852
rect 429 -76 487 -64
rect 429 -852 441 -76
rect 475 -852 487 -76
rect 429 -864 487 -852
rect 887 -76 945 -64
rect 887 -852 899 -76
rect 933 -852 945 -76
rect 887 -864 945 -852
rect 1345 -76 1403 -64
rect 1345 -852 1357 -76
rect 1391 -852 1403 -76
rect 1345 -864 1403 -852
rect 1803 -76 1861 -64
rect 1803 -852 1815 -76
rect 1849 -852 1861 -76
rect 1803 -864 1861 -852
<< mvpdiffc >>
rect -1849 76 -1815 852
rect -1391 76 -1357 852
rect -933 76 -899 852
rect -475 76 -441 852
rect -17 76 17 852
rect 441 76 475 852
rect 899 76 933 852
rect 1357 76 1391 852
rect 1815 76 1849 852
rect -1849 -852 -1815 -76
rect -1391 -852 -1357 -76
rect -933 -852 -899 -76
rect -475 -852 -441 -76
rect -17 -852 17 -76
rect 441 -852 475 -76
rect 899 -852 933 -76
rect 1357 -852 1391 -76
rect 1815 -852 1849 -76
<< mvnsubdiff >>
rect -1995 1083 1995 1095
rect -1995 1049 -1887 1083
rect 1887 1049 1995 1083
rect -1995 1037 1995 1049
rect -1995 987 -1937 1037
rect -1995 -987 -1983 987
rect -1949 -987 -1937 987
rect 1937 987 1995 1037
rect -1995 -1037 -1937 -987
rect 1937 -987 1949 987
rect 1983 -987 1995 987
rect 1937 -1037 1995 -987
rect -1995 -1049 1995 -1037
rect -1995 -1083 -1887 -1049
rect 1887 -1083 1995 -1049
rect -1995 -1095 1995 -1083
<< mvnsubdiffcont >>
rect -1887 1049 1887 1083
rect -1983 -987 -1949 987
rect 1949 -987 1983 987
rect -1887 -1083 1887 -1049
<< poly >>
rect -1803 945 -1403 961
rect -1803 911 -1787 945
rect -1419 911 -1403 945
rect -1803 864 -1403 911
rect -1345 945 -945 961
rect -1345 911 -1329 945
rect -961 911 -945 945
rect -1345 864 -945 911
rect -887 945 -487 961
rect -887 911 -871 945
rect -503 911 -487 945
rect -887 864 -487 911
rect -429 945 -29 961
rect -429 911 -413 945
rect -45 911 -29 945
rect -429 864 -29 911
rect 29 945 429 961
rect 29 911 45 945
rect 413 911 429 945
rect 29 864 429 911
rect 487 945 887 961
rect 487 911 503 945
rect 871 911 887 945
rect 487 864 887 911
rect 945 945 1345 961
rect 945 911 961 945
rect 1329 911 1345 945
rect 945 864 1345 911
rect 1403 945 1803 961
rect 1403 911 1419 945
rect 1787 911 1803 945
rect 1403 864 1803 911
rect -1803 17 -1403 64
rect -1803 -17 -1787 17
rect -1419 -17 -1403 17
rect -1803 -64 -1403 -17
rect -1345 17 -945 64
rect -1345 -17 -1329 17
rect -961 -17 -945 17
rect -1345 -64 -945 -17
rect -887 17 -487 64
rect -887 -17 -871 17
rect -503 -17 -487 17
rect -887 -64 -487 -17
rect -429 17 -29 64
rect -429 -17 -413 17
rect -45 -17 -29 17
rect -429 -64 -29 -17
rect 29 17 429 64
rect 29 -17 45 17
rect 413 -17 429 17
rect 29 -64 429 -17
rect 487 17 887 64
rect 487 -17 503 17
rect 871 -17 887 17
rect 487 -64 887 -17
rect 945 17 1345 64
rect 945 -17 961 17
rect 1329 -17 1345 17
rect 945 -64 1345 -17
rect 1403 17 1803 64
rect 1403 -17 1419 17
rect 1787 -17 1803 17
rect 1403 -64 1803 -17
rect -1803 -911 -1403 -864
rect -1803 -945 -1787 -911
rect -1419 -945 -1403 -911
rect -1803 -961 -1403 -945
rect -1345 -911 -945 -864
rect -1345 -945 -1329 -911
rect -961 -945 -945 -911
rect -1345 -961 -945 -945
rect -887 -911 -487 -864
rect -887 -945 -871 -911
rect -503 -945 -487 -911
rect -887 -961 -487 -945
rect -429 -911 -29 -864
rect -429 -945 -413 -911
rect -45 -945 -29 -911
rect -429 -961 -29 -945
rect 29 -911 429 -864
rect 29 -945 45 -911
rect 413 -945 429 -911
rect 29 -961 429 -945
rect 487 -911 887 -864
rect 487 -945 503 -911
rect 871 -945 887 -911
rect 487 -961 887 -945
rect 945 -911 1345 -864
rect 945 -945 961 -911
rect 1329 -945 1345 -911
rect 945 -961 1345 -945
rect 1403 -911 1803 -864
rect 1403 -945 1419 -911
rect 1787 -945 1803 -911
rect 1403 -961 1803 -945
<< polycont >>
rect -1787 911 -1419 945
rect -1329 911 -961 945
rect -871 911 -503 945
rect -413 911 -45 945
rect 45 911 413 945
rect 503 911 871 945
rect 961 911 1329 945
rect 1419 911 1787 945
rect -1787 -17 -1419 17
rect -1329 -17 -961 17
rect -871 -17 -503 17
rect -413 -17 -45 17
rect 45 -17 413 17
rect 503 -17 871 17
rect 961 -17 1329 17
rect 1419 -17 1787 17
rect -1787 -945 -1419 -911
rect -1329 -945 -961 -911
rect -871 -945 -503 -911
rect -413 -945 -45 -911
rect 45 -945 413 -911
rect 503 -945 871 -911
rect 961 -945 1329 -911
rect 1419 -945 1787 -911
<< locali >>
rect -1983 1049 -1887 1083
rect 1887 1049 1983 1083
rect -1983 987 -1949 1049
rect 1949 987 1983 1049
rect -1803 911 -1787 945
rect -1419 911 -1403 945
rect -1345 911 -1329 945
rect -961 911 -945 945
rect -887 911 -871 945
rect -503 911 -487 945
rect -429 911 -413 945
rect -45 911 -29 945
rect 29 911 45 945
rect 413 911 429 945
rect 487 911 503 945
rect 871 911 887 945
rect 945 911 961 945
rect 1329 911 1345 945
rect 1403 911 1419 945
rect 1787 911 1803 945
rect -1849 852 -1815 868
rect -1849 60 -1815 76
rect -1391 852 -1357 868
rect -1391 60 -1357 76
rect -933 852 -899 868
rect -933 60 -899 76
rect -475 852 -441 868
rect -475 60 -441 76
rect -17 852 17 868
rect -17 60 17 76
rect 441 852 475 868
rect 441 60 475 76
rect 899 852 933 868
rect 899 60 933 76
rect 1357 852 1391 868
rect 1357 60 1391 76
rect 1815 852 1849 868
rect 1815 60 1849 76
rect -1803 -17 -1787 17
rect -1419 -17 -1403 17
rect -1345 -17 -1329 17
rect -961 -17 -945 17
rect -887 -17 -871 17
rect -503 -17 -487 17
rect -429 -17 -413 17
rect -45 -17 -29 17
rect 29 -17 45 17
rect 413 -17 429 17
rect 487 -17 503 17
rect 871 -17 887 17
rect 945 -17 961 17
rect 1329 -17 1345 17
rect 1403 -17 1419 17
rect 1787 -17 1803 17
rect -1849 -76 -1815 -60
rect -1849 -868 -1815 -852
rect -1391 -76 -1357 -60
rect -1391 -868 -1357 -852
rect -933 -76 -899 -60
rect -933 -868 -899 -852
rect -475 -76 -441 -60
rect -475 -868 -441 -852
rect -17 -76 17 -60
rect -17 -868 17 -852
rect 441 -76 475 -60
rect 441 -868 475 -852
rect 899 -76 933 -60
rect 899 -868 933 -852
rect 1357 -76 1391 -60
rect 1357 -868 1391 -852
rect 1815 -76 1849 -60
rect 1815 -868 1849 -852
rect -1803 -945 -1787 -911
rect -1419 -945 -1403 -911
rect -1345 -945 -1329 -911
rect -961 -945 -945 -911
rect -887 -945 -871 -911
rect -503 -945 -487 -911
rect -429 -945 -413 -911
rect -45 -945 -29 -911
rect 29 -945 45 -911
rect 413 -945 429 -911
rect 487 -945 503 -911
rect 871 -945 887 -911
rect 945 -945 961 -911
rect 1329 -945 1345 -911
rect 1403 -945 1419 -911
rect 1787 -945 1803 -911
rect -1983 -1049 -1949 -987
rect 1949 -1049 1983 -987
rect -1983 -1083 -1887 -1049
rect 1887 -1083 1983 -1049
<< viali >>
rect -1787 911 -1419 945
rect -1329 911 -961 945
rect -871 911 -503 945
rect -413 911 -45 945
rect 45 911 413 945
rect 503 911 871 945
rect 961 911 1329 945
rect 1419 911 1787 945
rect -1849 76 -1815 852
rect -1391 76 -1357 852
rect -933 76 -899 852
rect -475 76 -441 852
rect -17 76 17 852
rect 441 76 475 852
rect 899 76 933 852
rect 1357 76 1391 852
rect 1815 76 1849 852
rect -1787 -17 -1419 17
rect -1329 -17 -961 17
rect -871 -17 -503 17
rect -413 -17 -45 17
rect 45 -17 413 17
rect 503 -17 871 17
rect 961 -17 1329 17
rect 1419 -17 1787 17
rect -1849 -852 -1815 -76
rect -1391 -852 -1357 -76
rect -933 -852 -899 -76
rect -475 -852 -441 -76
rect -17 -852 17 -76
rect 441 -852 475 -76
rect 899 -852 933 -76
rect 1357 -852 1391 -76
rect 1815 -852 1849 -76
rect -1787 -945 -1419 -911
rect -1329 -945 -961 -911
rect -871 -945 -503 -911
rect -413 -945 -45 -911
rect 45 -945 413 -911
rect 503 -945 871 -911
rect 961 -945 1329 -911
rect 1419 -945 1787 -911
<< metal1 >>
rect -1799 945 -1407 951
rect -1799 911 -1787 945
rect -1419 911 -1407 945
rect -1799 905 -1407 911
rect -1341 945 -949 951
rect -1341 911 -1329 945
rect -961 911 -949 945
rect -1341 905 -949 911
rect -883 945 -491 951
rect -883 911 -871 945
rect -503 911 -491 945
rect -883 905 -491 911
rect -425 945 -33 951
rect -425 911 -413 945
rect -45 911 -33 945
rect -425 905 -33 911
rect 33 945 425 951
rect 33 911 45 945
rect 413 911 425 945
rect 33 905 425 911
rect 491 945 883 951
rect 491 911 503 945
rect 871 911 883 945
rect 491 905 883 911
rect 949 945 1341 951
rect 949 911 961 945
rect 1329 911 1341 945
rect 949 905 1341 911
rect 1407 945 1799 951
rect 1407 911 1419 945
rect 1787 911 1799 945
rect 1407 905 1799 911
rect -1855 852 -1809 864
rect -1855 76 -1849 852
rect -1815 76 -1809 852
rect -1855 64 -1809 76
rect -1397 852 -1351 864
rect -1397 76 -1391 852
rect -1357 76 -1351 852
rect -1397 64 -1351 76
rect -939 852 -893 864
rect -939 76 -933 852
rect -899 76 -893 852
rect -939 64 -893 76
rect -481 852 -435 864
rect -481 76 -475 852
rect -441 76 -435 852
rect -481 64 -435 76
rect -23 852 23 864
rect -23 76 -17 852
rect 17 76 23 852
rect -23 64 23 76
rect 435 852 481 864
rect 435 76 441 852
rect 475 76 481 852
rect 435 64 481 76
rect 893 852 939 864
rect 893 76 899 852
rect 933 76 939 852
rect 893 64 939 76
rect 1351 852 1397 864
rect 1351 76 1357 852
rect 1391 76 1397 852
rect 1351 64 1397 76
rect 1809 852 1855 864
rect 1809 76 1815 852
rect 1849 76 1855 852
rect 1809 64 1855 76
rect -1799 17 -1407 23
rect -1799 -17 -1787 17
rect -1419 -17 -1407 17
rect -1799 -23 -1407 -17
rect -1341 17 -949 23
rect -1341 -17 -1329 17
rect -961 -17 -949 17
rect -1341 -23 -949 -17
rect -883 17 -491 23
rect -883 -17 -871 17
rect -503 -17 -491 17
rect -883 -23 -491 -17
rect -425 17 -33 23
rect -425 -17 -413 17
rect -45 -17 -33 17
rect -425 -23 -33 -17
rect 33 17 425 23
rect 33 -17 45 17
rect 413 -17 425 17
rect 33 -23 425 -17
rect 491 17 883 23
rect 491 -17 503 17
rect 871 -17 883 17
rect 491 -23 883 -17
rect 949 17 1341 23
rect 949 -17 961 17
rect 1329 -17 1341 17
rect 949 -23 1341 -17
rect 1407 17 1799 23
rect 1407 -17 1419 17
rect 1787 -17 1799 17
rect 1407 -23 1799 -17
rect -1855 -76 -1809 -64
rect -1855 -852 -1849 -76
rect -1815 -852 -1809 -76
rect -1855 -864 -1809 -852
rect -1397 -76 -1351 -64
rect -1397 -852 -1391 -76
rect -1357 -852 -1351 -76
rect -1397 -864 -1351 -852
rect -939 -76 -893 -64
rect -939 -852 -933 -76
rect -899 -852 -893 -76
rect -939 -864 -893 -852
rect -481 -76 -435 -64
rect -481 -852 -475 -76
rect -441 -852 -435 -76
rect -481 -864 -435 -852
rect -23 -76 23 -64
rect -23 -852 -17 -76
rect 17 -852 23 -76
rect -23 -864 23 -852
rect 435 -76 481 -64
rect 435 -852 441 -76
rect 475 -852 481 -76
rect 435 -864 481 -852
rect 893 -76 939 -64
rect 893 -852 899 -76
rect 933 -852 939 -76
rect 893 -864 939 -852
rect 1351 -76 1397 -64
rect 1351 -852 1357 -76
rect 1391 -852 1397 -76
rect 1351 -864 1397 -852
rect 1809 -76 1855 -64
rect 1809 -852 1815 -76
rect 1849 -852 1855 -76
rect 1809 -864 1855 -852
rect -1799 -911 -1407 -905
rect -1799 -945 -1787 -911
rect -1419 -945 -1407 -911
rect -1799 -951 -1407 -945
rect -1341 -911 -949 -905
rect -1341 -945 -1329 -911
rect -961 -945 -949 -911
rect -1341 -951 -949 -945
rect -883 -911 -491 -905
rect -883 -945 -871 -911
rect -503 -945 -491 -911
rect -883 -951 -491 -945
rect -425 -911 -33 -905
rect -425 -945 -413 -911
rect -45 -945 -33 -911
rect -425 -951 -33 -945
rect 33 -911 425 -905
rect 33 -945 45 -911
rect 413 -945 425 -911
rect 33 -951 425 -945
rect 491 -911 883 -905
rect 491 -945 503 -911
rect 871 -945 883 -911
rect 491 -951 883 -945
rect 949 -911 1341 -905
rect 949 -945 961 -911
rect 1329 -945 1341 -911
rect 949 -951 1341 -945
rect 1407 -911 1799 -905
rect 1407 -945 1419 -911
rect 1787 -945 1799 -911
rect 1407 -951 1799 -945
<< properties >>
string FIXED_BBOX -1966 -1066 1966 1066
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 2.0 m 2 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
