magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< metal4 >>
rect -1349 5839 1349 5880
rect -1349 3761 1093 5839
rect 1329 3761 1349 5839
rect -1349 3720 1349 3761
rect -1349 3439 1349 3480
rect -1349 1361 1093 3439
rect 1329 1361 1349 3439
rect -1349 1320 1349 1361
rect -1349 1039 1349 1080
rect -1349 -1039 1093 1039
rect 1329 -1039 1349 1039
rect -1349 -1080 1349 -1039
rect -1349 -1361 1349 -1320
rect -1349 -3439 1093 -1361
rect 1329 -3439 1349 -1361
rect -1349 -3480 1349 -3439
rect -1349 -3761 1349 -3720
rect -1349 -5839 1093 -3761
rect 1329 -5839 1349 -3761
rect -1349 -5880 1349 -5839
<< via4 >>
rect 1093 3761 1329 5839
rect 1093 1361 1329 3439
rect 1093 -1039 1329 1039
rect 1093 -3439 1329 -1361
rect 1093 -5839 1329 -3761
<< mimcap2 >>
rect -1269 5760 731 5800
rect -1269 3840 -1229 5760
rect 691 3840 731 5760
rect -1269 3800 731 3840
rect -1269 3360 731 3400
rect -1269 1440 -1229 3360
rect 691 1440 731 3360
rect -1269 1400 731 1440
rect -1269 960 731 1000
rect -1269 -960 -1229 960
rect 691 -960 731 960
rect -1269 -1000 731 -960
rect -1269 -1440 731 -1400
rect -1269 -3360 -1229 -1440
rect 691 -3360 731 -1440
rect -1269 -3400 731 -3360
rect -1269 -3840 731 -3800
rect -1269 -5760 -1229 -3840
rect 691 -5760 731 -3840
rect -1269 -5800 731 -5760
<< mimcap2contact >>
rect -1229 3840 691 5760
rect -1229 1440 691 3360
rect -1229 -960 691 960
rect -1229 -3360 691 -1440
rect -1229 -5760 691 -3840
<< metal5 >>
rect -429 5784 -109 6000
rect 1051 5839 1371 6000
rect -1253 5760 715 5784
rect -1253 3840 -1229 5760
rect 691 3840 715 5760
rect -1253 3816 715 3840
rect -429 3384 -109 3816
rect 1051 3761 1093 5839
rect 1329 3761 1371 5839
rect 1051 3439 1371 3761
rect -1253 3360 715 3384
rect -1253 1440 -1229 3360
rect 691 1440 715 3360
rect -1253 1416 715 1440
rect -429 984 -109 1416
rect 1051 1361 1093 3439
rect 1329 1361 1371 3439
rect 1051 1039 1371 1361
rect -1253 960 715 984
rect -1253 -960 -1229 960
rect 691 -960 715 960
rect -1253 -984 715 -960
rect -429 -1416 -109 -984
rect 1051 -1039 1093 1039
rect 1329 -1039 1371 1039
rect 1051 -1361 1371 -1039
rect -1253 -1440 715 -1416
rect -1253 -3360 -1229 -1440
rect 691 -3360 715 -1440
rect -1253 -3384 715 -3360
rect -429 -3816 -109 -3384
rect 1051 -3439 1093 -1361
rect 1329 -3439 1371 -1361
rect 1051 -3761 1371 -3439
rect -1253 -3840 715 -3816
rect -1253 -5760 -1229 -3840
rect 691 -5760 715 -3840
rect -1253 -5784 715 -5760
rect -429 -6000 -109 -5784
rect 1051 -5839 1093 -3761
rect 1329 -5839 1371 -3761
rect 1051 -6000 1371 -5839
<< properties >>
string FIXED_BBOX -1349 3720 811 5880
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
