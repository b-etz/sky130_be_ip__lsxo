magic
tech sky130A
timestamp 1713220443
<< pwell >>
rect -1343 -150 1343 150
<< mvnmos >>
rect -1229 -21 -429 21
rect -400 -21 400 21
rect 429 -21 1229 21
<< mvndiff >>
rect -1258 15 -1229 21
rect -1258 -15 -1252 15
rect -1235 -15 -1229 15
rect -1258 -21 -1229 -15
rect -429 15 -400 21
rect -429 -15 -423 15
rect -406 -15 -400 15
rect -429 -21 -400 -15
rect 400 15 429 21
rect 400 -15 406 15
rect 423 -15 429 15
rect 400 -21 429 -15
rect 1229 15 1258 21
rect 1229 -15 1235 15
rect 1252 -15 1258 15
rect 1229 -21 1258 -15
<< mvndiffc >>
rect -1252 -15 -1235 15
rect -423 -15 -406 15
rect 406 -15 423 15
rect 1235 -15 1252 15
<< mvpsubdiff >>
rect -1325 126 1325 132
rect -1325 109 -1271 126
rect 1271 109 1325 126
rect -1325 103 1325 109
rect -1325 78 -1296 103
rect -1325 -78 -1319 78
rect -1302 -78 -1296 78
rect 1296 78 1325 103
rect -1325 -103 -1296 -78
rect 1296 -78 1302 78
rect 1319 -78 1325 78
rect 1296 -103 1325 -78
rect -1325 -109 1325 -103
rect -1325 -126 -1271 -109
rect 1271 -126 1325 -109
rect -1325 -132 1325 -126
<< mvpsubdiffcont >>
rect -1271 109 1271 126
rect -1319 -78 -1302 78
rect 1302 -78 1319 78
rect -1271 -126 1271 -109
<< poly >>
rect -1229 57 -429 65
rect -1229 40 -1221 57
rect -437 40 -429 57
rect -1229 21 -429 40
rect -400 57 400 65
rect -400 40 -392 57
rect 392 40 400 57
rect -400 21 400 40
rect 429 57 1229 65
rect 429 40 437 57
rect 1221 40 1229 57
rect 429 21 1229 40
rect -1229 -40 -429 -21
rect -1229 -57 -1221 -40
rect -437 -57 -429 -40
rect -1229 -65 -429 -57
rect -400 -40 400 -21
rect -400 -57 -392 -40
rect 392 -57 400 -40
rect -400 -65 400 -57
rect 429 -40 1229 -21
rect 429 -57 437 -40
rect 1221 -57 1229 -40
rect 429 -65 1229 -57
<< polycont >>
rect -1221 40 -437 57
rect -392 40 392 57
rect 437 40 1221 57
rect -1221 -57 -437 -40
rect -392 -57 392 -40
rect 437 -57 1221 -40
<< locali >>
rect -1319 109 -1271 126
rect 1271 109 1319 126
rect -1319 78 -1302 109
rect 1302 78 1319 109
rect -1229 40 -1221 57
rect -437 40 -429 57
rect -400 40 -392 57
rect 392 40 400 57
rect 429 40 437 57
rect 1221 40 1229 57
rect -1252 15 -1235 23
rect -1252 -23 -1235 -15
rect -423 15 -406 23
rect -423 -23 -406 -15
rect 406 15 423 23
rect 406 -23 423 -15
rect 1235 15 1252 23
rect 1235 -23 1252 -15
rect -1229 -57 -1221 -40
rect -437 -57 -429 -40
rect -400 -57 -392 -40
rect 392 -57 400 -40
rect 429 -57 437 -40
rect 1221 -57 1229 -40
rect -1319 -109 -1302 -78
rect 1302 -109 1319 -78
rect -1319 -126 -1271 -109
rect 1271 -126 1319 -109
<< viali >>
rect -1221 40 -437 57
rect -392 40 392 57
rect 437 40 1221 57
rect -1252 -15 -1235 15
rect -423 -15 -406 15
rect 406 -15 423 15
rect 1235 -15 1252 15
rect -1221 -57 -437 -40
rect -392 -57 392 -40
rect 437 -57 1221 -40
<< metal1 >>
rect -1227 57 -431 60
rect -1227 40 -1221 57
rect -437 40 -431 57
rect -1227 37 -431 40
rect -398 57 398 60
rect -398 40 -392 57
rect 392 40 398 57
rect -398 37 398 40
rect 431 57 1227 60
rect 431 40 437 57
rect 1221 40 1227 57
rect 431 37 1227 40
rect -1255 15 -1232 21
rect -1255 -15 -1252 15
rect -1235 -15 -1232 15
rect -1255 -21 -1232 -15
rect -426 15 -403 21
rect -426 -15 -423 15
rect -406 -15 -403 15
rect -426 -21 -403 -15
rect 403 15 426 21
rect 403 -15 406 15
rect 423 -15 426 15
rect 403 -21 426 -15
rect 1232 15 1255 21
rect 1232 -15 1235 15
rect 1252 -15 1255 15
rect 1232 -21 1255 -15
rect -1227 -40 -431 -37
rect -1227 -57 -1221 -40
rect -437 -57 -431 -40
rect -1227 -60 -431 -57
rect -398 -40 398 -37
rect -398 -57 -392 -40
rect 392 -57 398 -40
rect -398 -60 398 -57
rect 431 -40 1227 -37
rect 431 -57 437 -40
rect 1221 -57 1227 -40
rect 431 -60 1227 -57
<< properties >>
string FIXED_BBOX -1310 -117 1310 117
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.420 l 8 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
