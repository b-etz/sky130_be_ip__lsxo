magic
tech sky130A
magscale 1 2
timestamp 1712965163
<< viali >>
rect 2726 -412 3746 -378
rect 750 -512 1316 -478
rect 750 -902 784 -512
rect 1282 -636 1316 -512
rect 2726 -962 2760 -412
rect 3712 -962 3746 -412
rect 2726 -996 3746 -962
rect 2726 -1118 3746 -1084
rect 758 -1564 792 -1426
rect 1272 -1564 1306 -1162
rect 758 -1598 1306 -1564
rect 2726 -1668 2760 -1118
rect 3712 -1668 3746 -1118
rect 4020 -1586 4054 -460
rect 4592 -494 5262 -460
rect 4624 -1586 4658 -494
rect 4020 -1620 4698 -1586
rect 5228 -1620 5262 -494
rect 2726 -1702 3746 -1668
<< metal1 >>
rect 652 -478 1434 -128
rect 652 -902 750 -478
rect 784 -574 1282 -512
rect 784 -902 792 -574
rect 932 -626 1134 -574
rect 1274 -636 1282 -574
rect 1316 -636 1434 -478
rect 1274 -650 1434 -636
rect 2580 -378 3852 -128
rect 652 -914 792 -902
rect 820 -694 1472 -688
rect 820 -782 1180 -694
rect 1464 -782 1472 -694
rect 820 -788 1472 -782
rect 820 -972 900 -788
rect 652 -1288 900 -972
rect 982 -988 1082 -850
rect 982 -994 1948 -988
rect 982 -1082 1650 -994
rect 1942 -1082 1948 -994
rect 982 -1088 1948 -1082
rect 2580 -996 2726 -378
rect 2760 -422 3712 -412
rect 2760 -948 2772 -422
rect 2804 -458 2904 -452
rect 2804 -552 2810 -458
rect 2898 -552 2904 -458
rect 2936 -552 3536 -422
rect 3568 -458 3668 -452
rect 3568 -552 3574 -458
rect 3662 -552 3668 -458
rect 2804 -812 2904 -552
rect 2936 -594 3534 -586
rect 2936 -778 2944 -594
rect 3526 -778 3534 -594
rect 2936 -788 3534 -778
rect 3568 -812 3668 -552
rect 2936 -948 3536 -822
rect 3700 -948 3712 -422
rect 2760 -962 3712 -948
rect 3746 -996 3852 -378
rect 2580 -1084 3852 -996
rect 982 -1226 1082 -1088
rect 1258 -1162 1418 -1148
rect 652 -1356 1210 -1288
rect 820 -1388 1210 -1356
rect 652 -1426 812 -1416
rect 652 -1598 758 -1426
rect 792 -1502 812 -1426
rect 932 -1502 1132 -1448
rect 1258 -1502 1272 -1162
rect 792 -1564 1272 -1502
rect 1306 -1598 1418 -1162
rect 652 -1950 1418 -1598
rect 2580 -1702 2726 -1084
rect 2760 -1132 3712 -1118
rect 2760 -1658 2772 -1132
rect 2936 -1258 3536 -1132
rect 2804 -1528 2904 -1268
rect 2936 -1300 3534 -1292
rect 2936 -1484 2944 -1300
rect 3526 -1484 3534 -1300
rect 2936 -1494 3534 -1484
rect 2804 -1622 2810 -1528
rect 2898 -1622 2904 -1528
rect 2804 -1628 2904 -1622
rect 2936 -1658 3536 -1526
rect 3568 -1528 3668 -1268
rect 3568 -1622 3574 -1528
rect 3662 -1622 3668 -1528
rect 3568 -1628 3668 -1622
rect 3700 -1658 3712 -1132
rect 2760 -1668 3712 -1658
rect 3746 -1702 3852 -1084
rect 2580 -1950 3852 -1702
rect 3912 -400 5370 -128
rect 3912 -460 4092 -400
rect 3912 -1620 4020 -460
rect 4054 -1484 4092 -460
rect 4230 -448 4450 -438
rect 4230 -628 4240 -448
rect 4440 -628 4450 -448
rect 4230 -638 4450 -628
rect 4564 -460 5370 -400
rect 4564 -494 4592 -460
rect 4148 -850 4528 -786
rect 4148 -1230 4248 -850
rect 4428 -1230 4528 -850
rect 4148 -1286 4528 -1230
rect 4240 -1484 4440 -1446
rect 4564 -1484 4624 -494
rect 4054 -1586 4624 -1484
rect 4658 -596 5228 -494
rect 4658 -1586 4718 -596
rect 4842 -634 5042 -596
rect 4756 -848 5136 -788
rect 4756 -1228 4852 -848
rect 5032 -1228 5136 -848
rect 4756 -1288 5136 -1228
rect 4698 -1620 4718 -1586
rect 3912 -1680 4718 -1620
rect 4832 -1450 5052 -1440
rect 4832 -1630 4842 -1450
rect 5042 -1630 5052 -1450
rect 4832 -1640 5052 -1630
rect 5190 -1620 5228 -596
rect 5262 -1620 5370 -460
rect 5190 -1680 5370 -1620
rect 3912 -1950 5370 -1680
<< via1 >>
rect 1180 -782 1464 -694
rect 1650 -1082 1942 -994
rect 2810 -552 2898 -458
rect 3574 -552 3662 -458
rect 2944 -778 3526 -594
rect 2944 -1484 3526 -1300
rect 2810 -1622 2898 -1528
rect 3574 -1622 3662 -1528
rect 4240 -628 4440 -448
rect 4248 -1230 4428 -850
rect 4852 -1228 5032 -848
rect 4842 -1630 5042 -1450
<< metal2 >>
rect 3742 -448 5670 -438
rect 1854 -458 3668 -452
rect 1854 -552 2810 -458
rect 2898 -552 3574 -458
rect 3662 -552 3668 -458
rect 1854 -558 3668 -552
rect 1854 -688 1954 -558
rect 1166 -694 1954 -688
rect 1166 -782 1180 -694
rect 1464 -782 1954 -694
rect 1166 -788 1954 -782
rect 2936 -588 3534 -586
rect 3742 -588 4240 -448
rect 2936 -594 4240 -588
rect 2936 -778 2944 -594
rect 3526 -628 4240 -594
rect 4440 -628 5670 -448
rect 3526 -638 5670 -628
rect 3526 -778 3942 -638
rect 2936 -788 3942 -778
rect 4240 -850 4438 -840
rect 1644 -994 2074 -988
rect 1644 -1082 1650 -994
rect 1942 -1082 2074 -994
rect 1644 -1088 2074 -1082
rect 1822 -1522 2074 -1088
rect 4240 -1230 4248 -850
rect 4428 -1230 4438 -850
rect 2936 -1300 3942 -1292
rect 2936 -1484 2944 -1300
rect 3526 -1440 3942 -1300
rect 4240 -1440 4438 -1230
rect 4844 -848 5042 -638
rect 4844 -1228 4852 -848
rect 5032 -1228 5042 -848
rect 4844 -1238 5042 -1228
rect 3526 -1450 5670 -1440
rect 3526 -1484 4842 -1450
rect 2936 -1492 4842 -1484
rect 2936 -1494 3534 -1492
rect 1822 -1528 3668 -1522
rect 1822 -1622 2810 -1528
rect 2898 -1622 3574 -1528
rect 3662 -1622 3668 -1528
rect 1822 -1628 3668 -1622
rect 1822 -1950 2074 -1628
rect 3742 -1630 4842 -1492
rect 5042 -1630 5670 -1450
rect 3742 -1640 5670 -1630
use sky130_fd_pr__nfet_01v8_69TQ3K  XM1
timestamp 1712965163
transform 0 -1 1032 1 0 -1338
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_3HMWVM  XM2
timestamp 1712965163
transform 0 -1 1033 1 0 -738
box -296 -319 296 319
use sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B  XM3
timestamp 1712965163
transform 0 1 3236 -1 0 -687
box -357 -558 357 558
use sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B  XM4
timestamp 1712965163
transform 0 1 3236 -1 0 -1393
box -357 -558 357 558
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM5
timestamp 1712965163
transform 0 1 4339 -1 0 -1040
box -658 -397 658 397
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM6
timestamp 1712965163
transform 0 1 4943 -1 0 -1040
box -658 -397 658 397
<< labels >>
flabel metal1 2580 -1950 3852 -1702 0 FreeSans 800 0 0 0 avss
port 3 nsew
flabel metal1 3912 -400 5370 -128 0 FreeSans 800 0 0 0 avdd
port 2 nsew
flabel metal1 652 -1950 1418 -1598 0 FreeSans 800 0 0 0 dvss
port 11 nsew
flabel metal1 652 -478 1434 -128 0 FreeSans 800 0 0 0 dvdd
port 12 nsew
flabel metal1 652 -1356 900 -972 0 FreeSans 800 0 0 0 in
port 1 nsew
flabel metal2 1822 -1950 2072 -1700 0 FreeSans 800 0 0 0 in_b
port 6 nsew
flabel metal2 4440 -638 5670 -438 0 FreeSans 800 0 0 0 out_b
port 10 nsew
flabel metal2 5042 -1640 5670 -1440 0 FreeSans 800 0 0 0 out
port 9 nsew
<< end >>
