magic
tech sky130A
magscale 1 2
timestamp 1712074743
<< error_p >>
rect 56788 -21011 56830 -19617
rect 57188 -21032 57230 -19638
rect 27600 -21414 27638 -21155
rect 28376 -21462 28412 -21430
rect 30387 -22368 30402 -22337
rect 30381 -22402 30402 -22368
rect 30387 -22433 30402 -22402
rect 30415 -22365 30430 -22334
rect 32525 -22365 32531 -22334
rect 30415 -22399 30436 -22365
rect 32519 -22399 32531 -22365
rect 30415 -22430 30430 -22399
rect 32525 -22430 32531 -22399
rect 32553 -22365 32559 -22334
rect 32553 -22399 32565 -22365
rect 32553 -22430 32559 -22399
rect 30387 -22912 30402 -22881
rect 30381 -22946 30402 -22912
rect 30387 -22977 30402 -22946
rect 30415 -22909 30430 -22878
rect 32525 -22909 32531 -22878
rect 30415 -22943 30436 -22909
rect 32519 -22943 32531 -22909
rect 30415 -22974 30430 -22943
rect 32525 -22974 32531 -22943
rect 32553 -22909 32559 -22878
rect 32553 -22943 32565 -22909
rect 32553 -22974 32559 -22943
rect 31035 -23468 31050 -23437
rect 31029 -23502 31050 -23468
rect 31035 -23533 31050 -23502
rect 31063 -23465 31078 -23434
rect 33173 -23465 33179 -23434
rect 31063 -23499 31084 -23465
rect 33167 -23499 33179 -23465
rect 31063 -23530 31078 -23499
rect 33173 -23530 33179 -23499
rect 33201 -23465 33207 -23434
rect 33201 -23499 33213 -23465
rect 33201 -23530 33207 -23499
rect 31035 -24012 31050 -23981
rect 31029 -24046 31050 -24012
rect 31035 -24077 31050 -24046
rect 31063 -24009 31078 -23978
rect 33173 -24009 33179 -23978
rect 31063 -24043 31084 -24009
rect 33167 -24043 33179 -24009
rect 31063 -24074 31078 -24043
rect 33173 -24074 33179 -24043
rect 33201 -24009 33207 -23978
rect 33201 -24043 33213 -24009
rect 33201 -24074 33207 -24043
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use sky130_fd_pr__cap_mim_m3_1_4HHTN9  sky130_fd_pr__cap_mim_m3_1_4HHTN9_0
timestamp 1712073300
transform 1 0 21614 0 1 -17914
box -1186 -4640 1186 4640
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 2060 0 1 -1966
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x2
timestamp 1707688321
transform 1 0 2128 0 1 -6994
box -38 -48 314 592
use level_shift  x3
timestamp 1712071977
transform 1 0 3450 0 1 -836
box 0 -2800 3195 480
use level_shift  x4
timestamp 1712071977
transform 1 0 3306 0 1 -5912
box 0 -2800 3195 480
use bias_gen  x5
timestamp 1712073863
transform 1 0 35464 0 1 -13246
box 0 -3410 15466 14020
use dout_amp  x6
timestamp 1712071977
transform 1 0 49316 0 1 -16565
box 0 -18731 16839 3379
use ripl_dly_clk_buf  x7
timestamp 1712074743
transform 1 0 26499 0 1 -22222
box -53 -3176 8856 1139
use sky130_fd_pr__cap_mim_m3_1_KAF84V  XC1
timestamp 1712073300
transform 1 0 12864 0 1 -22240
box -886 -3440 886 3440
use sky130_fd_pr__cap_mim_m3_1_4RVTN9  XC2
timestamp 1712073300
transform 1 0 57742 0 1 -742
box -5104 -9280 5104 9280
use sky130_fd_pr__cap_mim_m3_1_4HHTN9  XC3
timestamp 1712073300
transform 1 0 9312 0 1 -26182
box -1186 -4640 1186 4640
use sky130_fd_pr__nfet_g5v0d10v5_LB4DGD  XM1
timestamp 1712071977
transform 1 0 20474 0 1 -65
box -278 -5239 278 5239
use sky130_fd_pr__pfet_g5v0d10v5_CLHFX9  XM2
timestamp 1712071977
transform 1 0 24424 0 1 345
box -458 -5359 458 5359
use sky130_fd_pr__nfet_01v8_AHZR5K  XM3
timestamp 1712071977
transform 1 0 35056 0 1 -18500
box -596 -260 596 260
use sky130_fd_pr__nfet_01v8_HZ6WG7  XM4
timestamp 1712071977
transform 1 0 64008 0 1 -7677
box -296 -285 296 285
use sky130_fd_pr__nfet_g5v0d10v5_9PDQJ3  XM5
timestamp 1712071977
transform 1 0 22432 0 1 -362
box -278 -2694 278 2694
use sky130_fd_pr__pfet_g5v0d10v5_E43JVH  XM6
timestamp 1712071977
transform 1 0 18040 0 1 -939
box -308 -2769 308 2769
use sky130_fd_pr__pfet_01v8_3H68VM  XM7
timestamp 1712071977
transform 1 0 64008 0 1 -6049
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_EDBGFV  XM8
timestamp 1712071977
transform 1 0 32622 0 1 2659
box -246 -5281 246 5281
use sky130_fd_pr__pfet_g5v0d10v5_KL3SY6  XM9
timestamp 1712071977
transform 1 0 34860 0 1 -2939
box -308 -697 308 697
use sky130_fd_pr__nfet_01v8_8WM5KZ  XM11
timestamp 1712071977
transform 1 0 27402 0 1 -41
box -246 -5191 246 5191
use sky130_fd_pr__res_xhigh_po_0p35_LKPHWV  XR2
timestamp 1712073300
transform 1 0 11706 0 1 -11556
box -4268 -5782 4268 5782
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 dvdd
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 dvss
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 ibias
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 ena
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 standby
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 dout
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 xin
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 xout
port 9 nsew
<< end >>
