magic
tech sky130A
magscale 1 2
timestamp 1713144909
<< pwell >>
rect -2193 -11582 2193 11582
<< psubdiff >>
rect -2157 11512 -2061 11546
rect 2061 11512 2157 11546
rect -2157 11450 -2123 11512
rect 2123 11450 2157 11512
rect -2157 -11512 -2123 -11450
rect 2123 -11512 2157 -11450
rect -2157 -11546 -2061 -11512
rect 2061 -11546 2157 -11512
<< psubdiffcont >>
rect -2061 11512 2061 11546
rect -2157 -11450 -2123 11450
rect 2123 -11450 2157 11450
rect -2061 -11546 2061 -11512
<< xpolycontact >>
rect -2027 10984 -1957 11416
rect -2027 -11416 -1957 -10984
rect -1861 10984 -1791 11416
rect -1861 -11416 -1791 -10984
rect -1695 10984 -1625 11416
rect -1695 -11416 -1625 -10984
rect -1529 10984 -1459 11416
rect -1529 -11416 -1459 -10984
rect -1363 10984 -1293 11416
rect -1363 -11416 -1293 -10984
rect -1197 10984 -1127 11416
rect -1197 -11416 -1127 -10984
rect -1031 10984 -961 11416
rect -1031 -11416 -961 -10984
rect -865 10984 -795 11416
rect -865 -11416 -795 -10984
rect -699 10984 -629 11416
rect -699 -11416 -629 -10984
rect -533 10984 -463 11416
rect -533 -11416 -463 -10984
rect -367 10984 -297 11416
rect -367 -11416 -297 -10984
rect -201 10984 -131 11416
rect -201 -11416 -131 -10984
rect -35 10984 35 11416
rect -35 -11416 35 -10984
rect 131 10984 201 11416
rect 131 -11416 201 -10984
rect 297 10984 367 11416
rect 297 -11416 367 -10984
rect 463 10984 533 11416
rect 463 -11416 533 -10984
rect 629 10984 699 11416
rect 629 -11416 699 -10984
rect 795 10984 865 11416
rect 795 -11416 865 -10984
rect 961 10984 1031 11416
rect 961 -11416 1031 -10984
rect 1127 10984 1197 11416
rect 1127 -11416 1197 -10984
rect 1293 10984 1363 11416
rect 1293 -11416 1363 -10984
rect 1459 10984 1529 11416
rect 1459 -11416 1529 -10984
rect 1625 10984 1695 11416
rect 1625 -11416 1695 -10984
rect 1791 10984 1861 11416
rect 1791 -11416 1861 -10984
rect 1957 10984 2027 11416
rect 1957 -11416 2027 -10984
<< xpolyres >>
rect -2027 -10984 -1957 10984
rect -1861 -10984 -1791 10984
rect -1695 -10984 -1625 10984
rect -1529 -10984 -1459 10984
rect -1363 -10984 -1293 10984
rect -1197 -10984 -1127 10984
rect -1031 -10984 -961 10984
rect -865 -10984 -795 10984
rect -699 -10984 -629 10984
rect -533 -10984 -463 10984
rect -367 -10984 -297 10984
rect -201 -10984 -131 10984
rect -35 -10984 35 10984
rect 131 -10984 201 10984
rect 297 -10984 367 10984
rect 463 -10984 533 10984
rect 629 -10984 699 10984
rect 795 -10984 865 10984
rect 961 -10984 1031 10984
rect 1127 -10984 1197 10984
rect 1293 -10984 1363 10984
rect 1459 -10984 1529 10984
rect 1625 -10984 1695 10984
rect 1791 -10984 1861 10984
rect 1957 -10984 2027 10984
<< locali >>
rect -2157 11512 -2061 11546
rect 2061 11512 2157 11546
rect -2157 11450 -2123 11512
rect 2123 11450 2157 11512
rect -2157 -11512 -2123 -11450
rect 2123 -11512 2157 -11450
rect -2157 -11546 -2061 -11512
rect 2061 -11546 2157 -11512
<< viali >>
rect -2011 11001 -1973 11398
rect -1845 11001 -1807 11398
rect -1679 11001 -1641 11398
rect -1513 11001 -1475 11398
rect -1347 11001 -1309 11398
rect -1181 11001 -1143 11398
rect -1015 11001 -977 11398
rect -849 11001 -811 11398
rect -683 11001 -645 11398
rect -517 11001 -479 11398
rect -351 11001 -313 11398
rect -185 11001 -147 11398
rect -19 11001 19 11398
rect 147 11001 185 11398
rect 313 11001 351 11398
rect 479 11001 517 11398
rect 645 11001 683 11398
rect 811 11001 849 11398
rect 977 11001 1015 11398
rect 1143 11001 1181 11398
rect 1309 11001 1347 11398
rect 1475 11001 1513 11398
rect 1641 11001 1679 11398
rect 1807 11001 1845 11398
rect 1973 11001 2011 11398
rect -2011 -11398 -1973 -11001
rect -1845 -11398 -1807 -11001
rect -1679 -11398 -1641 -11001
rect -1513 -11398 -1475 -11001
rect -1347 -11398 -1309 -11001
rect -1181 -11398 -1143 -11001
rect -1015 -11398 -977 -11001
rect -849 -11398 -811 -11001
rect -683 -11398 -645 -11001
rect -517 -11398 -479 -11001
rect -351 -11398 -313 -11001
rect -185 -11398 -147 -11001
rect -19 -11398 19 -11001
rect 147 -11398 185 -11001
rect 313 -11398 351 -11001
rect 479 -11398 517 -11001
rect 645 -11398 683 -11001
rect 811 -11398 849 -11001
rect 977 -11398 1015 -11001
rect 1143 -11398 1181 -11001
rect 1309 -11398 1347 -11001
rect 1475 -11398 1513 -11001
rect 1641 -11398 1679 -11001
rect 1807 -11398 1845 -11001
rect 1973 -11398 2011 -11001
<< metal1 >>
rect -2017 11398 -1967 11410
rect -2017 11001 -2011 11398
rect -1973 11001 -1967 11398
rect -2017 10989 -1967 11001
rect -1851 11398 -1801 11410
rect -1851 11001 -1845 11398
rect -1807 11001 -1801 11398
rect -1851 10989 -1801 11001
rect -1685 11398 -1635 11410
rect -1685 11001 -1679 11398
rect -1641 11001 -1635 11398
rect -1685 10989 -1635 11001
rect -1519 11398 -1469 11410
rect -1519 11001 -1513 11398
rect -1475 11001 -1469 11398
rect -1519 10989 -1469 11001
rect -1353 11398 -1303 11410
rect -1353 11001 -1347 11398
rect -1309 11001 -1303 11398
rect -1353 10989 -1303 11001
rect -1187 11398 -1137 11410
rect -1187 11001 -1181 11398
rect -1143 11001 -1137 11398
rect -1187 10989 -1137 11001
rect -1021 11398 -971 11410
rect -1021 11001 -1015 11398
rect -977 11001 -971 11398
rect -1021 10989 -971 11001
rect -855 11398 -805 11410
rect -855 11001 -849 11398
rect -811 11001 -805 11398
rect -855 10989 -805 11001
rect -689 11398 -639 11410
rect -689 11001 -683 11398
rect -645 11001 -639 11398
rect -689 10989 -639 11001
rect -523 11398 -473 11410
rect -523 11001 -517 11398
rect -479 11001 -473 11398
rect -523 10989 -473 11001
rect -357 11398 -307 11410
rect -357 11001 -351 11398
rect -313 11001 -307 11398
rect -357 10989 -307 11001
rect -191 11398 -141 11410
rect -191 11001 -185 11398
rect -147 11001 -141 11398
rect -191 10989 -141 11001
rect -25 11398 25 11410
rect -25 11001 -19 11398
rect 19 11001 25 11398
rect -25 10989 25 11001
rect 141 11398 191 11410
rect 141 11001 147 11398
rect 185 11001 191 11398
rect 141 10989 191 11001
rect 307 11398 357 11410
rect 307 11001 313 11398
rect 351 11001 357 11398
rect 307 10989 357 11001
rect 473 11398 523 11410
rect 473 11001 479 11398
rect 517 11001 523 11398
rect 473 10989 523 11001
rect 639 11398 689 11410
rect 639 11001 645 11398
rect 683 11001 689 11398
rect 639 10989 689 11001
rect 805 11398 855 11410
rect 805 11001 811 11398
rect 849 11001 855 11398
rect 805 10989 855 11001
rect 971 11398 1021 11410
rect 971 11001 977 11398
rect 1015 11001 1021 11398
rect 971 10989 1021 11001
rect 1137 11398 1187 11410
rect 1137 11001 1143 11398
rect 1181 11001 1187 11398
rect 1137 10989 1187 11001
rect 1303 11398 1353 11410
rect 1303 11001 1309 11398
rect 1347 11001 1353 11398
rect 1303 10989 1353 11001
rect 1469 11398 1519 11410
rect 1469 11001 1475 11398
rect 1513 11001 1519 11398
rect 1469 10989 1519 11001
rect 1635 11398 1685 11410
rect 1635 11001 1641 11398
rect 1679 11001 1685 11398
rect 1635 10989 1685 11001
rect 1801 11398 1851 11410
rect 1801 11001 1807 11398
rect 1845 11001 1851 11398
rect 1801 10989 1851 11001
rect 1967 11398 2017 11410
rect 1967 11001 1973 11398
rect 2011 11001 2017 11398
rect 1967 10989 2017 11001
rect -2017 -11001 -1967 -10989
rect -2017 -11398 -2011 -11001
rect -1973 -11398 -1967 -11001
rect -2017 -11410 -1967 -11398
rect -1851 -11001 -1801 -10989
rect -1851 -11398 -1845 -11001
rect -1807 -11398 -1801 -11001
rect -1851 -11410 -1801 -11398
rect -1685 -11001 -1635 -10989
rect -1685 -11398 -1679 -11001
rect -1641 -11398 -1635 -11001
rect -1685 -11410 -1635 -11398
rect -1519 -11001 -1469 -10989
rect -1519 -11398 -1513 -11001
rect -1475 -11398 -1469 -11001
rect -1519 -11410 -1469 -11398
rect -1353 -11001 -1303 -10989
rect -1353 -11398 -1347 -11001
rect -1309 -11398 -1303 -11001
rect -1353 -11410 -1303 -11398
rect -1187 -11001 -1137 -10989
rect -1187 -11398 -1181 -11001
rect -1143 -11398 -1137 -11001
rect -1187 -11410 -1137 -11398
rect -1021 -11001 -971 -10989
rect -1021 -11398 -1015 -11001
rect -977 -11398 -971 -11001
rect -1021 -11410 -971 -11398
rect -855 -11001 -805 -10989
rect -855 -11398 -849 -11001
rect -811 -11398 -805 -11001
rect -855 -11410 -805 -11398
rect -689 -11001 -639 -10989
rect -689 -11398 -683 -11001
rect -645 -11398 -639 -11001
rect -689 -11410 -639 -11398
rect -523 -11001 -473 -10989
rect -523 -11398 -517 -11001
rect -479 -11398 -473 -11001
rect -523 -11410 -473 -11398
rect -357 -11001 -307 -10989
rect -357 -11398 -351 -11001
rect -313 -11398 -307 -11001
rect -357 -11410 -307 -11398
rect -191 -11001 -141 -10989
rect -191 -11398 -185 -11001
rect -147 -11398 -141 -11001
rect -191 -11410 -141 -11398
rect -25 -11001 25 -10989
rect -25 -11398 -19 -11001
rect 19 -11398 25 -11001
rect -25 -11410 25 -11398
rect 141 -11001 191 -10989
rect 141 -11398 147 -11001
rect 185 -11398 191 -11001
rect 141 -11410 191 -11398
rect 307 -11001 357 -10989
rect 307 -11398 313 -11001
rect 351 -11398 357 -11001
rect 307 -11410 357 -11398
rect 473 -11001 523 -10989
rect 473 -11398 479 -11001
rect 517 -11398 523 -11001
rect 473 -11410 523 -11398
rect 639 -11001 689 -10989
rect 639 -11398 645 -11001
rect 683 -11398 689 -11001
rect 639 -11410 689 -11398
rect 805 -11001 855 -10989
rect 805 -11398 811 -11001
rect 849 -11398 855 -11001
rect 805 -11410 855 -11398
rect 971 -11001 1021 -10989
rect 971 -11398 977 -11001
rect 1015 -11398 1021 -11001
rect 971 -11410 1021 -11398
rect 1137 -11001 1187 -10989
rect 1137 -11398 1143 -11001
rect 1181 -11398 1187 -11001
rect 1137 -11410 1187 -11398
rect 1303 -11001 1353 -10989
rect 1303 -11398 1309 -11001
rect 1347 -11398 1353 -11001
rect 1303 -11410 1353 -11398
rect 1469 -11001 1519 -10989
rect 1469 -11398 1475 -11001
rect 1513 -11398 1519 -11001
rect 1469 -11410 1519 -11398
rect 1635 -11001 1685 -10989
rect 1635 -11398 1641 -11001
rect 1679 -11398 1685 -11001
rect 1635 -11410 1685 -11398
rect 1801 -11001 1851 -10989
rect 1801 -11398 1807 -11001
rect 1845 -11398 1851 -11001
rect 1801 -11410 1851 -11398
rect 1967 -11001 2017 -10989
rect 1967 -11398 1973 -11001
rect 2011 -11398 2017 -11001
rect 1967 -11410 2017 -11398
<< properties >>
string FIXED_BBOX -2140 -11529 2140 11529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 110 m 1 nx 25 wmin 0.350 lmin 0.50 rho 2000 val 629.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
