magic
tech sky130A
magscale 1 2
timestamp 1712853061
<< nwell >>
rect -1312 -683 1312 683
<< pmos >>
rect -1116 64 -716 464
rect -658 64 -258 464
rect -200 64 200 464
rect 258 64 658 464
rect 716 64 1116 464
rect -1116 -464 -716 -64
rect -658 -464 -258 -64
rect -200 -464 200 -64
rect 258 -464 658 -64
rect 716 -464 1116 -64
<< pdiff >>
rect -1174 452 -1116 464
rect -1174 76 -1162 452
rect -1128 76 -1116 452
rect -1174 64 -1116 76
rect -716 452 -658 464
rect -716 76 -704 452
rect -670 76 -658 452
rect -716 64 -658 76
rect -258 452 -200 464
rect -258 76 -246 452
rect -212 76 -200 452
rect -258 64 -200 76
rect 200 452 258 464
rect 200 76 212 452
rect 246 76 258 452
rect 200 64 258 76
rect 658 452 716 464
rect 658 76 670 452
rect 704 76 716 452
rect 658 64 716 76
rect 1116 452 1174 464
rect 1116 76 1128 452
rect 1162 76 1174 452
rect 1116 64 1174 76
rect -1174 -76 -1116 -64
rect -1174 -452 -1162 -76
rect -1128 -452 -1116 -76
rect -1174 -464 -1116 -452
rect -716 -76 -658 -64
rect -716 -452 -704 -76
rect -670 -452 -658 -76
rect -716 -464 -658 -452
rect -258 -76 -200 -64
rect -258 -452 -246 -76
rect -212 -452 -200 -76
rect -258 -464 -200 -452
rect 200 -76 258 -64
rect 200 -452 212 -76
rect 246 -452 258 -76
rect 200 -464 258 -452
rect 658 -76 716 -64
rect 658 -452 670 -76
rect 704 -452 716 -76
rect 658 -464 716 -452
rect 1116 -76 1174 -64
rect 1116 -452 1128 -76
rect 1162 -452 1174 -76
rect 1116 -464 1174 -452
<< pdiffc >>
rect -1162 76 -1128 452
rect -704 76 -670 452
rect -246 76 -212 452
rect 212 76 246 452
rect 670 76 704 452
rect 1128 76 1162 452
rect -1162 -452 -1128 -76
rect -704 -452 -670 -76
rect -246 -452 -212 -76
rect 212 -452 246 -76
rect 670 -452 704 -76
rect 1128 -452 1162 -76
<< nsubdiff >>
rect -1276 613 -1180 647
rect 1180 613 1276 647
rect -1276 551 -1242 613
rect 1242 551 1276 613
rect -1276 -613 -1242 -551
rect 1242 -613 1276 -551
rect -1276 -647 -1180 -613
rect 1180 -647 1276 -613
<< nsubdiffcont >>
rect -1180 613 1180 647
rect -1276 -551 -1242 551
rect 1242 -551 1276 551
rect -1180 -647 1180 -613
<< poly >>
rect -1116 545 -716 561
rect -1116 511 -1100 545
rect -732 511 -716 545
rect -1116 464 -716 511
rect -658 545 -258 561
rect -658 511 -642 545
rect -274 511 -258 545
rect -658 464 -258 511
rect -200 545 200 561
rect -200 511 -184 545
rect 184 511 200 545
rect -200 464 200 511
rect 258 545 658 561
rect 258 511 274 545
rect 642 511 658 545
rect 258 464 658 511
rect 716 545 1116 561
rect 716 511 732 545
rect 1100 511 1116 545
rect 716 464 1116 511
rect -1116 17 -716 64
rect -1116 -17 -1100 17
rect -732 -17 -716 17
rect -1116 -64 -716 -17
rect -658 17 -258 64
rect -658 -17 -642 17
rect -274 -17 -258 17
rect -658 -64 -258 -17
rect -200 17 200 64
rect -200 -17 -184 17
rect 184 -17 200 17
rect -200 -64 200 -17
rect 258 17 658 64
rect 258 -17 274 17
rect 642 -17 658 17
rect 258 -64 658 -17
rect 716 17 1116 64
rect 716 -17 732 17
rect 1100 -17 1116 17
rect 716 -64 1116 -17
rect -1116 -511 -716 -464
rect -1116 -545 -1100 -511
rect -732 -545 -716 -511
rect -1116 -561 -716 -545
rect -658 -511 -258 -464
rect -658 -545 -642 -511
rect -274 -545 -258 -511
rect -658 -561 -258 -545
rect -200 -511 200 -464
rect -200 -545 -184 -511
rect 184 -545 200 -511
rect -200 -561 200 -545
rect 258 -511 658 -464
rect 258 -545 274 -511
rect 642 -545 658 -511
rect 258 -561 658 -545
rect 716 -511 1116 -464
rect 716 -545 732 -511
rect 1100 -545 1116 -511
rect 716 -561 1116 -545
<< polycont >>
rect -1100 511 -732 545
rect -642 511 -274 545
rect -184 511 184 545
rect 274 511 642 545
rect 732 511 1100 545
rect -1100 -17 -732 17
rect -642 -17 -274 17
rect -184 -17 184 17
rect 274 -17 642 17
rect 732 -17 1100 17
rect -1100 -545 -732 -511
rect -642 -545 -274 -511
rect -184 -545 184 -511
rect 274 -545 642 -511
rect 732 -545 1100 -511
<< locali >>
rect -1276 613 -1180 647
rect 1180 613 1276 647
rect -1276 551 -1242 613
rect 1242 551 1276 613
rect -1116 511 -1100 545
rect -732 511 -716 545
rect -658 511 -642 545
rect -274 511 -258 545
rect -200 511 -184 545
rect 184 511 200 545
rect 258 511 274 545
rect 642 511 658 545
rect 716 511 732 545
rect 1100 511 1116 545
rect -1162 452 -1128 468
rect -1162 60 -1128 76
rect -704 452 -670 468
rect -704 60 -670 76
rect -246 452 -212 468
rect -246 60 -212 76
rect 212 452 246 468
rect 212 60 246 76
rect 670 452 704 468
rect 670 60 704 76
rect 1128 452 1162 468
rect 1128 60 1162 76
rect -1116 -17 -1100 17
rect -732 -17 -716 17
rect -658 -17 -642 17
rect -274 -17 -258 17
rect -200 -17 -184 17
rect 184 -17 200 17
rect 258 -17 274 17
rect 642 -17 658 17
rect 716 -17 732 17
rect 1100 -17 1116 17
rect -1162 -76 -1128 -60
rect -1162 -468 -1128 -452
rect -704 -76 -670 -60
rect -704 -468 -670 -452
rect -246 -76 -212 -60
rect -246 -468 -212 -452
rect 212 -76 246 -60
rect 212 -468 246 -452
rect 670 -76 704 -60
rect 670 -468 704 -452
rect 1128 -76 1162 -60
rect 1128 -468 1162 -452
rect -1116 -545 -1100 -511
rect -732 -545 -716 -511
rect -658 -545 -642 -511
rect -274 -545 -258 -511
rect -200 -545 -184 -511
rect 184 -545 200 -511
rect 258 -545 274 -511
rect 642 -545 658 -511
rect 716 -545 732 -511
rect 1100 -545 1116 -511
rect -1276 -613 -1242 -551
rect 1242 -613 1276 -551
rect -1276 -647 -1180 -613
rect 1180 -647 1276 -613
<< viali >>
rect -1100 511 -732 545
rect -642 511 -274 545
rect -184 511 184 545
rect 274 511 642 545
rect 732 511 1100 545
rect -1162 76 -1128 452
rect -704 76 -670 452
rect -246 76 -212 452
rect 212 76 246 452
rect 670 76 704 452
rect 1128 76 1162 452
rect -1100 -17 -732 17
rect -642 -17 -274 17
rect -184 -17 184 17
rect 274 -17 642 17
rect 732 -17 1100 17
rect -1162 -452 -1128 -76
rect -704 -452 -670 -76
rect -246 -452 -212 -76
rect 212 -452 246 -76
rect 670 -452 704 -76
rect 1128 -452 1162 -76
rect -1100 -545 -732 -511
rect -642 -545 -274 -511
rect -184 -545 184 -511
rect 274 -545 642 -511
rect 732 -545 1100 -511
<< metal1 >>
rect -1112 545 -720 551
rect -1112 511 -1100 545
rect -732 511 -720 545
rect -1112 505 -720 511
rect -654 545 -262 551
rect -654 511 -642 545
rect -274 511 -262 545
rect -654 505 -262 511
rect -196 545 196 551
rect -196 511 -184 545
rect 184 511 196 545
rect -196 505 196 511
rect 262 545 654 551
rect 262 511 274 545
rect 642 511 654 545
rect 262 505 654 511
rect 720 545 1112 551
rect 720 511 732 545
rect 1100 511 1112 545
rect 720 505 1112 511
rect -1168 452 -1122 464
rect -1168 76 -1162 452
rect -1128 76 -1122 452
rect -1168 64 -1122 76
rect -710 452 -664 464
rect -710 76 -704 452
rect -670 76 -664 452
rect -710 64 -664 76
rect -252 452 -206 464
rect -252 76 -246 452
rect -212 76 -206 452
rect -252 64 -206 76
rect 206 452 252 464
rect 206 76 212 452
rect 246 76 252 452
rect 206 64 252 76
rect 664 452 710 464
rect 664 76 670 452
rect 704 76 710 452
rect 664 64 710 76
rect 1122 452 1168 464
rect 1122 76 1128 452
rect 1162 76 1168 452
rect 1122 64 1168 76
rect -1112 17 -720 23
rect -1112 -17 -1100 17
rect -732 -17 -720 17
rect -1112 -23 -720 -17
rect -654 17 -262 23
rect -654 -17 -642 17
rect -274 -17 -262 17
rect -654 -23 -262 -17
rect -196 17 196 23
rect -196 -17 -184 17
rect 184 -17 196 17
rect -196 -23 196 -17
rect 262 17 654 23
rect 262 -17 274 17
rect 642 -17 654 17
rect 262 -23 654 -17
rect 720 17 1112 23
rect 720 -17 732 17
rect 1100 -17 1112 17
rect 720 -23 1112 -17
rect -1168 -76 -1122 -64
rect -1168 -452 -1162 -76
rect -1128 -452 -1122 -76
rect -1168 -464 -1122 -452
rect -710 -76 -664 -64
rect -710 -452 -704 -76
rect -670 -452 -664 -76
rect -710 -464 -664 -452
rect -252 -76 -206 -64
rect -252 -452 -246 -76
rect -212 -452 -206 -76
rect -252 -464 -206 -452
rect 206 -76 252 -64
rect 206 -452 212 -76
rect 246 -452 252 -76
rect 206 -464 252 -452
rect 664 -76 710 -64
rect 664 -452 670 -76
rect 704 -452 710 -76
rect 664 -464 710 -452
rect 1122 -76 1168 -64
rect 1122 -452 1128 -76
rect 1162 -452 1168 -76
rect 1122 -464 1168 -452
rect -1112 -511 -720 -505
rect -1112 -545 -1100 -511
rect -732 -545 -720 -511
rect -1112 -551 -720 -545
rect -654 -511 -262 -505
rect -654 -545 -642 -511
rect -274 -545 -262 -511
rect -654 -551 -262 -545
rect -196 -511 196 -505
rect -196 -545 -184 -511
rect 184 -545 196 -511
rect -196 -551 196 -545
rect 262 -511 654 -505
rect 262 -545 274 -511
rect 642 -545 654 -511
rect 262 -551 654 -545
rect 720 -511 1112 -505
rect 720 -545 732 -511
rect 1100 -545 1112 -511
rect 720 -551 1112 -545
<< properties >>
string FIXED_BBOX -1259 -630 1259 630
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 2.0 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
