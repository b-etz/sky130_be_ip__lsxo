magic
tech sky130A
magscale 1 2
timestamp 1713142410
<< pwell >>
rect -1363 -7182 1363 7182
<< psubdiff >>
rect -1327 7112 -1231 7146
rect 1231 7112 1327 7146
rect -1327 7050 -1293 7112
rect 1293 7050 1327 7112
rect -1327 -7112 -1293 -7050
rect 1293 -7112 1327 -7050
rect -1327 -7146 -1231 -7112
rect 1231 -7146 1327 -7112
<< psubdiffcont >>
rect -1231 7112 1231 7146
rect -1327 -7050 -1293 7050
rect 1293 -7050 1327 7050
rect -1231 -7146 1231 -7112
<< xpolycontact >>
rect -1197 6584 -1127 7016
rect -1197 -7016 -1127 -6584
rect -1031 6584 -961 7016
rect -1031 -7016 -961 -6584
rect -865 6584 -795 7016
rect -865 -7016 -795 -6584
rect -699 6584 -629 7016
rect -699 -7016 -629 -6584
rect -533 6584 -463 7016
rect -533 -7016 -463 -6584
rect -367 6584 -297 7016
rect -367 -7016 -297 -6584
rect -201 6584 -131 7016
rect -201 -7016 -131 -6584
rect -35 6584 35 7016
rect -35 -7016 35 -6584
rect 131 6584 201 7016
rect 131 -7016 201 -6584
rect 297 6584 367 7016
rect 297 -7016 367 -6584
rect 463 6584 533 7016
rect 463 -7016 533 -6584
rect 629 6584 699 7016
rect 629 -7016 699 -6584
rect 795 6584 865 7016
rect 795 -7016 865 -6584
rect 961 6584 1031 7016
rect 961 -7016 1031 -6584
rect 1127 6584 1197 7016
rect 1127 -7016 1197 -6584
<< xpolyres >>
rect -1197 -6584 -1127 6584
rect -1031 -6584 -961 6584
rect -865 -6584 -795 6584
rect -699 -6584 -629 6584
rect -533 -6584 -463 6584
rect -367 -6584 -297 6584
rect -201 -6584 -131 6584
rect -35 -6584 35 6584
rect 131 -6584 201 6584
rect 297 -6584 367 6584
rect 463 -6584 533 6584
rect 629 -6584 699 6584
rect 795 -6584 865 6584
rect 961 -6584 1031 6584
rect 1127 -6584 1197 6584
<< locali >>
rect -1327 7112 -1231 7146
rect 1231 7112 1327 7146
rect -1327 7050 -1293 7112
rect 1293 7050 1327 7112
rect -1327 -7112 -1293 -7050
rect 1293 -7112 1327 -7050
rect -1327 -7146 -1231 -7112
rect 1231 -7146 1327 -7112
<< viali >>
rect -1181 6601 -1143 6998
rect -1015 6601 -977 6998
rect -849 6601 -811 6998
rect -683 6601 -645 6998
rect -517 6601 -479 6998
rect -351 6601 -313 6998
rect -185 6601 -147 6998
rect -19 6601 19 6998
rect 147 6601 185 6998
rect 313 6601 351 6998
rect 479 6601 517 6998
rect 645 6601 683 6998
rect 811 6601 849 6998
rect 977 6601 1015 6998
rect 1143 6601 1181 6998
rect -1181 -6998 -1143 -6601
rect -1015 -6998 -977 -6601
rect -849 -6998 -811 -6601
rect -683 -6998 -645 -6601
rect -517 -6998 -479 -6601
rect -351 -6998 -313 -6601
rect -185 -6998 -147 -6601
rect -19 -6998 19 -6601
rect 147 -6998 185 -6601
rect 313 -6998 351 -6601
rect 479 -6998 517 -6601
rect 645 -6998 683 -6601
rect 811 -6998 849 -6601
rect 977 -6998 1015 -6601
rect 1143 -6998 1181 -6601
<< metal1 >>
rect -1187 6998 -1137 7010
rect -1187 6601 -1181 6998
rect -1143 6601 -1137 6998
rect -1187 6589 -1137 6601
rect -1021 6998 -971 7010
rect -1021 6601 -1015 6998
rect -977 6601 -971 6998
rect -1021 6589 -971 6601
rect -855 6998 -805 7010
rect -855 6601 -849 6998
rect -811 6601 -805 6998
rect -855 6589 -805 6601
rect -689 6998 -639 7010
rect -689 6601 -683 6998
rect -645 6601 -639 6998
rect -689 6589 -639 6601
rect -523 6998 -473 7010
rect -523 6601 -517 6998
rect -479 6601 -473 6998
rect -523 6589 -473 6601
rect -357 6998 -307 7010
rect -357 6601 -351 6998
rect -313 6601 -307 6998
rect -357 6589 -307 6601
rect -191 6998 -141 7010
rect -191 6601 -185 6998
rect -147 6601 -141 6998
rect -191 6589 -141 6601
rect -25 6998 25 7010
rect -25 6601 -19 6998
rect 19 6601 25 6998
rect -25 6589 25 6601
rect 141 6998 191 7010
rect 141 6601 147 6998
rect 185 6601 191 6998
rect 141 6589 191 6601
rect 307 6998 357 7010
rect 307 6601 313 6998
rect 351 6601 357 6998
rect 307 6589 357 6601
rect 473 6998 523 7010
rect 473 6601 479 6998
rect 517 6601 523 6998
rect 473 6589 523 6601
rect 639 6998 689 7010
rect 639 6601 645 6998
rect 683 6601 689 6998
rect 639 6589 689 6601
rect 805 6998 855 7010
rect 805 6601 811 6998
rect 849 6601 855 6998
rect 805 6589 855 6601
rect 971 6998 1021 7010
rect 971 6601 977 6998
rect 1015 6601 1021 6998
rect 971 6589 1021 6601
rect 1137 6998 1187 7010
rect 1137 6601 1143 6998
rect 1181 6601 1187 6998
rect 1137 6589 1187 6601
rect -1187 -6601 -1137 -6589
rect -1187 -6998 -1181 -6601
rect -1143 -6998 -1137 -6601
rect -1187 -7010 -1137 -6998
rect -1021 -6601 -971 -6589
rect -1021 -6998 -1015 -6601
rect -977 -6998 -971 -6601
rect -1021 -7010 -971 -6998
rect -855 -6601 -805 -6589
rect -855 -6998 -849 -6601
rect -811 -6998 -805 -6601
rect -855 -7010 -805 -6998
rect -689 -6601 -639 -6589
rect -689 -6998 -683 -6601
rect -645 -6998 -639 -6601
rect -689 -7010 -639 -6998
rect -523 -6601 -473 -6589
rect -523 -6998 -517 -6601
rect -479 -6998 -473 -6601
rect -523 -7010 -473 -6998
rect -357 -6601 -307 -6589
rect -357 -6998 -351 -6601
rect -313 -6998 -307 -6601
rect -357 -7010 -307 -6998
rect -191 -6601 -141 -6589
rect -191 -6998 -185 -6601
rect -147 -6998 -141 -6601
rect -191 -7010 -141 -6998
rect -25 -6601 25 -6589
rect -25 -6998 -19 -6601
rect 19 -6998 25 -6601
rect -25 -7010 25 -6998
rect 141 -6601 191 -6589
rect 141 -6998 147 -6601
rect 185 -6998 191 -6601
rect 141 -7010 191 -6998
rect 307 -6601 357 -6589
rect 307 -6998 313 -6601
rect 351 -6998 357 -6601
rect 307 -7010 357 -6998
rect 473 -6601 523 -6589
rect 473 -6998 479 -6601
rect 517 -6998 523 -6601
rect 473 -7010 523 -6998
rect 639 -6601 689 -6589
rect 639 -6998 645 -6601
rect 683 -6998 689 -6601
rect 639 -7010 689 -6998
rect 805 -6601 855 -6589
rect 805 -6998 811 -6601
rect 849 -6998 855 -6601
rect 805 -7010 855 -6998
rect 971 -6601 1021 -6589
rect 971 -6998 977 -6601
rect 1015 -6998 1021 -6601
rect 971 -7010 1021 -6998
rect 1137 -6601 1187 -6589
rect 1137 -6998 1143 -6601
rect 1181 -6998 1187 -6601
rect 1137 -7010 1187 -6998
<< properties >>
string FIXED_BBOX -1310 -7129 1310 7129
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 66 m 1 nx 15 wmin 0.350 lmin 0.50 rho 2000 val 378.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
