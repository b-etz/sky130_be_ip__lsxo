magic
tech sky130A
magscale 1 2
timestamp 1713220443
<< viali >>
rect 2726 -380 3744 -284
rect 750 -512 1316 -478
rect 750 -574 784 -512
rect 1282 -574 1316 -512
rect 4622 -536 5296 -416
rect 2726 -1088 3744 -992
rect 758 -1564 792 -1502
rect 1272 -1564 1306 -1502
rect 758 -1598 1306 -1564
rect 3984 -1664 4658 -1544
rect 2728 -1794 3746 -1698
<< metal1 >>
rect 652 -478 1434 -128
rect 652 -574 750 -478
rect 784 -526 1282 -512
rect 784 -574 796 -526
rect 652 -580 796 -574
rect 960 -586 1106 -526
rect 1270 -574 1282 -526
rect 1316 -574 1434 -478
rect 1270 -580 1434 -574
rect 2580 -284 3852 -128
rect 2580 -380 2726 -284
rect 3744 -380 3852 -284
rect 2580 -422 3852 -380
rect 932 -626 1134 -586
rect 820 -694 1472 -688
rect 820 -782 1180 -694
rect 1464 -782 1472 -694
rect 820 -788 1472 -782
rect 820 -972 900 -788
rect 652 -1288 900 -972
rect 982 -988 1082 -850
rect 2580 -948 2772 -422
rect 2838 -498 2904 -492
rect 2838 -552 2844 -498
rect 2898 -552 2904 -498
rect 3136 -502 3336 -422
rect 3568 -498 3634 -492
rect 2936 -552 3536 -502
rect 3568 -552 3574 -498
rect 3628 -552 3634 -498
rect 2838 -558 2904 -552
rect 2846 -812 2904 -558
rect 3568 -558 3634 -552
rect 2936 -594 3534 -586
rect 2936 -778 2944 -594
rect 3526 -778 3534 -594
rect 2936 -788 3534 -778
rect 3568 -812 3626 -558
rect 2936 -868 3536 -822
rect 3136 -948 3336 -868
rect 3700 -948 3852 -422
rect 982 -994 1472 -988
rect 982 -1082 1160 -994
rect 1466 -1082 1472 -994
rect 982 -1088 1472 -1082
rect 2580 -992 3852 -948
rect 2580 -1088 2726 -992
rect 3744 -1088 3852 -992
rect 982 -1226 1082 -1088
rect 2580 -1132 3852 -1088
rect 652 -1356 1210 -1288
rect 820 -1388 1210 -1356
rect 932 -1492 1132 -1448
rect 652 -1502 804 -1496
rect 652 -1598 758 -1502
rect 792 -1552 804 -1502
rect 958 -1552 1104 -1492
rect 1260 -1502 1418 -1496
rect 1260 -1552 1272 -1502
rect 792 -1564 1272 -1552
rect 1306 -1598 1418 -1502
rect 652 -1950 1418 -1598
rect 2580 -1658 2772 -1132
rect 3136 -1212 3336 -1132
rect 2936 -1258 3536 -1212
rect 2846 -1522 2904 -1268
rect 2936 -1300 3534 -1292
rect 2936 -1484 2944 -1300
rect 3526 -1484 3534 -1300
rect 2936 -1494 3534 -1484
rect 2838 -1528 2904 -1522
rect 3568 -1522 3626 -1268
rect 2838 -1582 2844 -1528
rect 2898 -1582 2904 -1528
rect 2936 -1578 3536 -1526
rect 3568 -1528 3634 -1522
rect 2838 -1588 2904 -1582
rect 3136 -1658 3336 -1578
rect 3568 -1582 3574 -1528
rect 3628 -1582 3634 -1528
rect 3568 -1588 3634 -1582
rect 3700 -1658 3852 -1132
rect 2580 -1698 3852 -1658
rect 2580 -1794 2728 -1698
rect 3746 -1794 3852 -1698
rect 2580 -1950 3852 -1794
rect 3912 -378 5370 -128
rect 3912 -1520 4086 -378
rect 4588 -416 5370 -378
rect 4230 -448 4450 -438
rect 4230 -628 4240 -448
rect 4440 -628 4450 -448
rect 4230 -638 4450 -628
rect 4588 -536 4622 -416
rect 5296 -536 5370 -416
rect 4588 -560 5370 -536
rect 4148 -850 4528 -786
rect 4148 -1230 4248 -850
rect 4428 -1230 4528 -850
rect 4148 -1286 4528 -1230
rect 4238 -1520 4440 -1446
rect 4588 -1520 4696 -560
rect 4842 -634 5044 -560
rect 4756 -848 5136 -788
rect 4756 -1228 4852 -848
rect 5032 -1228 5136 -848
rect 4756 -1288 5136 -1228
rect 3912 -1544 4696 -1520
rect 3912 -1664 3984 -1544
rect 4658 -1664 4696 -1544
rect 4832 -1450 5052 -1440
rect 4832 -1630 4842 -1450
rect 5042 -1630 5052 -1450
rect 4832 -1640 5052 -1630
rect 3912 -1700 4696 -1664
rect 5196 -1700 5370 -560
rect 3912 -1950 5370 -1700
<< via1 >>
rect 1180 -782 1464 -694
rect 2844 -552 2898 -498
rect 3574 -552 3628 -498
rect 2944 -778 3526 -594
rect 1160 -1082 1466 -994
rect 2944 -1484 3526 -1300
rect 2844 -1582 2898 -1528
rect 3574 -1582 3628 -1528
rect 4240 -628 4440 -448
rect 4248 -1230 4428 -850
rect 4852 -1228 5032 -848
rect 4842 -1630 5042 -1450
<< metal2 >>
rect 3742 -448 5670 -438
rect 1854 -498 3634 -452
rect 1854 -552 2844 -498
rect 2898 -552 3574 -498
rect 3628 -552 3634 -498
rect 1854 -558 3634 -552
rect 1854 -688 1954 -558
rect 1166 -694 1954 -688
rect 1166 -782 1180 -694
rect 1464 -782 1954 -694
rect 1166 -788 1954 -782
rect 2936 -588 3534 -586
rect 3742 -588 4240 -448
rect 2936 -594 4240 -588
rect 2936 -778 2944 -594
rect 3526 -628 4240 -594
rect 4440 -628 5670 -448
rect 3526 -638 5670 -628
rect 3526 -778 3942 -638
rect 2936 -788 3942 -778
rect 4240 -850 4438 -840
rect 1152 -994 2074 -988
rect 1152 -1082 1160 -994
rect 1466 -1082 2074 -994
rect 1152 -1088 2074 -1082
rect 1822 -1522 2074 -1088
rect 4240 -1230 4248 -850
rect 4428 -1230 4438 -850
rect 2936 -1300 3942 -1292
rect 2936 -1484 2944 -1300
rect 3526 -1440 3942 -1300
rect 4240 -1440 4438 -1230
rect 4844 -848 5042 -638
rect 4844 -1228 4852 -848
rect 5032 -1228 5042 -848
rect 4844 -1238 5042 -1228
rect 3526 -1450 5670 -1440
rect 3526 -1484 4842 -1450
rect 2936 -1492 4842 -1484
rect 2936 -1494 3534 -1492
rect 1822 -1528 3634 -1522
rect 1822 -1582 2844 -1528
rect 2898 -1582 3574 -1528
rect 3628 -1582 3634 -1528
rect 1822 -1628 3634 -1582
rect 3742 -1630 4842 -1492
rect 5042 -1630 5670 -1450
rect 3742 -1640 5670 -1630
use sky130_fd_pr__nfet_01v8_69TQ3K  XM1
timestamp 1713220443
transform 0 -1 1032 1 0 -1338
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_3HMWVM  XM2
timestamp 1713220443
transform 0 -1 1033 1 0 -738
box -296 -319 296 319
use sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B  XM3
timestamp 1713220443
transform 0 1 3236 -1 0 -687
box -357 -558 357 558
use sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B  XM4
timestamp 1713220443
transform 0 1 3236 -1 0 -1393
box -357 -558 357 558
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM5
timestamp 1713220443
transform 0 1 4339 -1 0 -1040
box -658 -397 658 397
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM6
timestamp 1713220443
transform 0 1 4943 -1 0 -1040
box -658 -397 658 397
<< labels >>
flabel metal1 652 -478 1434 -128 0 FreeSans 1600 0 0 0 dvdd
port 1 nsew
flabel metal1 652 -1950 1418 -1598 0 FreeSans 1600 0 0 0 dvss
port 2 nsew
flabel metal1 3912 -378 5370 -128 0 FreeSans 1600 0 0 0 avdd
port 3 nsew
flabel metal1 2580 -1950 3852 -1794 0 FreeSans 1200 0 0 0 avss
port 4 nsew
flabel metal1 652 -1356 900 -972 0 FreeSans 1200 0 0 0 in
port 5 nsew
flabel metal2 1822 -1628 2074 -988 0 FreeSans 800 0 0 0 in_b
port 6 nsew
flabel metal2 4440 -638 5670 -438 0 FreeSans 1200 0 0 0 out_b
port 7 nsew
flabel metal2 5042 -1640 5670 -1440 0 FreeSans 1200 0 0 0 out
port 8 nsew
<< end >>
