magic
tech sky130A
magscale 1 2
timestamp 1712073300
<< pwell >>
rect -4268 -260582 4268 260582
<< psubdiff >>
rect -4232 260512 -4136 260546
rect 4136 260512 4232 260546
rect -4232 260450 -4198 260512
rect 4198 260450 4232 260512
rect -4232 -260512 -4198 -260450
rect 4198 -260512 4232 -260450
rect -4232 -260546 -4136 -260512
rect 4136 -260546 4232 -260512
<< psubdiffcont >>
rect -4136 260512 4136 260546
rect -4232 -260450 -4198 260450
rect 4198 -260450 4232 260450
rect -4136 -260546 4136 -260512
<< xpolycontact >>
rect -4102 259984 -4032 260416
rect -4102 -260416 -4032 -259984
rect -3936 259984 -3866 260416
rect -3936 -260416 -3866 -259984
rect -3770 259984 -3700 260416
rect -3770 -260416 -3700 -259984
rect -3604 259984 -3534 260416
rect -3604 -260416 -3534 -259984
rect -3438 259984 -3368 260416
rect -3438 -260416 -3368 -259984
rect -3272 259984 -3202 260416
rect -3272 -260416 -3202 -259984
rect -3106 259984 -3036 260416
rect -3106 -260416 -3036 -259984
rect -2940 259984 -2870 260416
rect -2940 -260416 -2870 -259984
rect -2774 259984 -2704 260416
rect -2774 -260416 -2704 -259984
rect -2608 259984 -2538 260416
rect -2608 -260416 -2538 -259984
rect -2442 259984 -2372 260416
rect -2442 -260416 -2372 -259984
rect -2276 259984 -2206 260416
rect -2276 -260416 -2206 -259984
rect -2110 259984 -2040 260416
rect -2110 -260416 -2040 -259984
rect -1944 259984 -1874 260416
rect -1944 -260416 -1874 -259984
rect -1778 259984 -1708 260416
rect -1778 -260416 -1708 -259984
rect -1612 259984 -1542 260416
rect -1612 -260416 -1542 -259984
rect -1446 259984 -1376 260416
rect -1446 -260416 -1376 -259984
rect -1280 259984 -1210 260416
rect -1280 -260416 -1210 -259984
rect -1114 259984 -1044 260416
rect -1114 -260416 -1044 -259984
rect -948 259984 -878 260416
rect -948 -260416 -878 -259984
rect -782 259984 -712 260416
rect -782 -260416 -712 -259984
rect -616 259984 -546 260416
rect -616 -260416 -546 -259984
rect -450 259984 -380 260416
rect -450 -260416 -380 -259984
rect -284 259984 -214 260416
rect -284 -260416 -214 -259984
rect -118 259984 -48 260416
rect -118 -260416 -48 -259984
rect 48 259984 118 260416
rect 48 -260416 118 -259984
rect 214 259984 284 260416
rect 214 -260416 284 -259984
rect 380 259984 450 260416
rect 380 -260416 450 -259984
rect 546 259984 616 260416
rect 546 -260416 616 -259984
rect 712 259984 782 260416
rect 712 -260416 782 -259984
rect 878 259984 948 260416
rect 878 -260416 948 -259984
rect 1044 259984 1114 260416
rect 1044 -260416 1114 -259984
rect 1210 259984 1280 260416
rect 1210 -260416 1280 -259984
rect 1376 259984 1446 260416
rect 1376 -260416 1446 -259984
rect 1542 259984 1612 260416
rect 1542 -260416 1612 -259984
rect 1708 259984 1778 260416
rect 1708 -260416 1778 -259984
rect 1874 259984 1944 260416
rect 1874 -260416 1944 -259984
rect 2040 259984 2110 260416
rect 2040 -260416 2110 -259984
rect 2206 259984 2276 260416
rect 2206 -260416 2276 -259984
rect 2372 259984 2442 260416
rect 2372 -260416 2442 -259984
rect 2538 259984 2608 260416
rect 2538 -260416 2608 -259984
rect 2704 259984 2774 260416
rect 2704 -260416 2774 -259984
rect 2870 259984 2940 260416
rect 2870 -260416 2940 -259984
rect 3036 259984 3106 260416
rect 3036 -260416 3106 -259984
rect 3202 259984 3272 260416
rect 3202 -260416 3272 -259984
rect 3368 259984 3438 260416
rect 3368 -260416 3438 -259984
rect 3534 259984 3604 260416
rect 3534 -260416 3604 -259984
rect 3700 259984 3770 260416
rect 3700 -260416 3770 -259984
rect 3866 259984 3936 260416
rect 3866 -260416 3936 -259984
rect 4032 259984 4102 260416
rect 4032 -260416 4102 -259984
<< xpolyres >>
rect -4102 -259984 -4032 259984
rect -3936 -259984 -3866 259984
rect -3770 -259984 -3700 259984
rect -3604 -259984 -3534 259984
rect -3438 -259984 -3368 259984
rect -3272 -259984 -3202 259984
rect -3106 -259984 -3036 259984
rect -2940 -259984 -2870 259984
rect -2774 -259984 -2704 259984
rect -2608 -259984 -2538 259984
rect -2442 -259984 -2372 259984
rect -2276 -259984 -2206 259984
rect -2110 -259984 -2040 259984
rect -1944 -259984 -1874 259984
rect -1778 -259984 -1708 259984
rect -1612 -259984 -1542 259984
rect -1446 -259984 -1376 259984
rect -1280 -259984 -1210 259984
rect -1114 -259984 -1044 259984
rect -948 -259984 -878 259984
rect -782 -259984 -712 259984
rect -616 -259984 -546 259984
rect -450 -259984 -380 259984
rect -284 -259984 -214 259984
rect -118 -259984 -48 259984
rect 48 -259984 118 259984
rect 214 -259984 284 259984
rect 380 -259984 450 259984
rect 546 -259984 616 259984
rect 712 -259984 782 259984
rect 878 -259984 948 259984
rect 1044 -259984 1114 259984
rect 1210 -259984 1280 259984
rect 1376 -259984 1446 259984
rect 1542 -259984 1612 259984
rect 1708 -259984 1778 259984
rect 1874 -259984 1944 259984
rect 2040 -259984 2110 259984
rect 2206 -259984 2276 259984
rect 2372 -259984 2442 259984
rect 2538 -259984 2608 259984
rect 2704 -259984 2774 259984
rect 2870 -259984 2940 259984
rect 3036 -259984 3106 259984
rect 3202 -259984 3272 259984
rect 3368 -259984 3438 259984
rect 3534 -259984 3604 259984
rect 3700 -259984 3770 259984
rect 3866 -259984 3936 259984
rect 4032 -259984 4102 259984
<< locali >>
rect -4232 260512 -4136 260546
rect 4136 260512 4232 260546
rect -4232 260450 -4198 260512
rect 4198 260450 4232 260512
rect -4232 -260512 -4198 -260450
rect 4198 -260512 4232 -260450
rect -4232 -260546 -4136 -260512
rect 4136 -260546 4232 -260512
<< viali >>
rect -4086 260001 -4048 260398
rect -3920 260001 -3882 260398
rect -3754 260001 -3716 260398
rect -3588 260001 -3550 260398
rect -3422 260001 -3384 260398
rect -3256 260001 -3218 260398
rect -3090 260001 -3052 260398
rect -2924 260001 -2886 260398
rect -2758 260001 -2720 260398
rect -2592 260001 -2554 260398
rect -2426 260001 -2388 260398
rect -2260 260001 -2222 260398
rect -2094 260001 -2056 260398
rect -1928 260001 -1890 260398
rect -1762 260001 -1724 260398
rect -1596 260001 -1558 260398
rect -1430 260001 -1392 260398
rect -1264 260001 -1226 260398
rect -1098 260001 -1060 260398
rect -932 260001 -894 260398
rect -766 260001 -728 260398
rect -600 260001 -562 260398
rect -434 260001 -396 260398
rect -268 260001 -230 260398
rect -102 260001 -64 260398
rect 64 260001 102 260398
rect 230 260001 268 260398
rect 396 260001 434 260398
rect 562 260001 600 260398
rect 728 260001 766 260398
rect 894 260001 932 260398
rect 1060 260001 1098 260398
rect 1226 260001 1264 260398
rect 1392 260001 1430 260398
rect 1558 260001 1596 260398
rect 1724 260001 1762 260398
rect 1890 260001 1928 260398
rect 2056 260001 2094 260398
rect 2222 260001 2260 260398
rect 2388 260001 2426 260398
rect 2554 260001 2592 260398
rect 2720 260001 2758 260398
rect 2886 260001 2924 260398
rect 3052 260001 3090 260398
rect 3218 260001 3256 260398
rect 3384 260001 3422 260398
rect 3550 260001 3588 260398
rect 3716 260001 3754 260398
rect 3882 260001 3920 260398
rect 4048 260001 4086 260398
rect -4086 -260398 -4048 -260001
rect -3920 -260398 -3882 -260001
rect -3754 -260398 -3716 -260001
rect -3588 -260398 -3550 -260001
rect -3422 -260398 -3384 -260001
rect -3256 -260398 -3218 -260001
rect -3090 -260398 -3052 -260001
rect -2924 -260398 -2886 -260001
rect -2758 -260398 -2720 -260001
rect -2592 -260398 -2554 -260001
rect -2426 -260398 -2388 -260001
rect -2260 -260398 -2222 -260001
rect -2094 -260398 -2056 -260001
rect -1928 -260398 -1890 -260001
rect -1762 -260398 -1724 -260001
rect -1596 -260398 -1558 -260001
rect -1430 -260398 -1392 -260001
rect -1264 -260398 -1226 -260001
rect -1098 -260398 -1060 -260001
rect -932 -260398 -894 -260001
rect -766 -260398 -728 -260001
rect -600 -260398 -562 -260001
rect -434 -260398 -396 -260001
rect -268 -260398 -230 -260001
rect -102 -260398 -64 -260001
rect 64 -260398 102 -260001
rect 230 -260398 268 -260001
rect 396 -260398 434 -260001
rect 562 -260398 600 -260001
rect 728 -260398 766 -260001
rect 894 -260398 932 -260001
rect 1060 -260398 1098 -260001
rect 1226 -260398 1264 -260001
rect 1392 -260398 1430 -260001
rect 1558 -260398 1596 -260001
rect 1724 -260398 1762 -260001
rect 1890 -260398 1928 -260001
rect 2056 -260398 2094 -260001
rect 2222 -260398 2260 -260001
rect 2388 -260398 2426 -260001
rect 2554 -260398 2592 -260001
rect 2720 -260398 2758 -260001
rect 2886 -260398 2924 -260001
rect 3052 -260398 3090 -260001
rect 3218 -260398 3256 -260001
rect 3384 -260398 3422 -260001
rect 3550 -260398 3588 -260001
rect 3716 -260398 3754 -260001
rect 3882 -260398 3920 -260001
rect 4048 -260398 4086 -260001
<< metal1 >>
rect -4092 260398 -4042 260410
rect -4092 260001 -4086 260398
rect -4048 260001 -4042 260398
rect -4092 259989 -4042 260001
rect -3926 260398 -3876 260410
rect -3926 260001 -3920 260398
rect -3882 260001 -3876 260398
rect -3926 259989 -3876 260001
rect -3760 260398 -3710 260410
rect -3760 260001 -3754 260398
rect -3716 260001 -3710 260398
rect -3760 259989 -3710 260001
rect -3594 260398 -3544 260410
rect -3594 260001 -3588 260398
rect -3550 260001 -3544 260398
rect -3594 259989 -3544 260001
rect -3428 260398 -3378 260410
rect -3428 260001 -3422 260398
rect -3384 260001 -3378 260398
rect -3428 259989 -3378 260001
rect -3262 260398 -3212 260410
rect -3262 260001 -3256 260398
rect -3218 260001 -3212 260398
rect -3262 259989 -3212 260001
rect -3096 260398 -3046 260410
rect -3096 260001 -3090 260398
rect -3052 260001 -3046 260398
rect -3096 259989 -3046 260001
rect -2930 260398 -2880 260410
rect -2930 260001 -2924 260398
rect -2886 260001 -2880 260398
rect -2930 259989 -2880 260001
rect -2764 260398 -2714 260410
rect -2764 260001 -2758 260398
rect -2720 260001 -2714 260398
rect -2764 259989 -2714 260001
rect -2598 260398 -2548 260410
rect -2598 260001 -2592 260398
rect -2554 260001 -2548 260398
rect -2598 259989 -2548 260001
rect -2432 260398 -2382 260410
rect -2432 260001 -2426 260398
rect -2388 260001 -2382 260398
rect -2432 259989 -2382 260001
rect -2266 260398 -2216 260410
rect -2266 260001 -2260 260398
rect -2222 260001 -2216 260398
rect -2266 259989 -2216 260001
rect -2100 260398 -2050 260410
rect -2100 260001 -2094 260398
rect -2056 260001 -2050 260398
rect -2100 259989 -2050 260001
rect -1934 260398 -1884 260410
rect -1934 260001 -1928 260398
rect -1890 260001 -1884 260398
rect -1934 259989 -1884 260001
rect -1768 260398 -1718 260410
rect -1768 260001 -1762 260398
rect -1724 260001 -1718 260398
rect -1768 259989 -1718 260001
rect -1602 260398 -1552 260410
rect -1602 260001 -1596 260398
rect -1558 260001 -1552 260398
rect -1602 259989 -1552 260001
rect -1436 260398 -1386 260410
rect -1436 260001 -1430 260398
rect -1392 260001 -1386 260398
rect -1436 259989 -1386 260001
rect -1270 260398 -1220 260410
rect -1270 260001 -1264 260398
rect -1226 260001 -1220 260398
rect -1270 259989 -1220 260001
rect -1104 260398 -1054 260410
rect -1104 260001 -1098 260398
rect -1060 260001 -1054 260398
rect -1104 259989 -1054 260001
rect -938 260398 -888 260410
rect -938 260001 -932 260398
rect -894 260001 -888 260398
rect -938 259989 -888 260001
rect -772 260398 -722 260410
rect -772 260001 -766 260398
rect -728 260001 -722 260398
rect -772 259989 -722 260001
rect -606 260398 -556 260410
rect -606 260001 -600 260398
rect -562 260001 -556 260398
rect -606 259989 -556 260001
rect -440 260398 -390 260410
rect -440 260001 -434 260398
rect -396 260001 -390 260398
rect -440 259989 -390 260001
rect -274 260398 -224 260410
rect -274 260001 -268 260398
rect -230 260001 -224 260398
rect -274 259989 -224 260001
rect -108 260398 -58 260410
rect -108 260001 -102 260398
rect -64 260001 -58 260398
rect -108 259989 -58 260001
rect 58 260398 108 260410
rect 58 260001 64 260398
rect 102 260001 108 260398
rect 58 259989 108 260001
rect 224 260398 274 260410
rect 224 260001 230 260398
rect 268 260001 274 260398
rect 224 259989 274 260001
rect 390 260398 440 260410
rect 390 260001 396 260398
rect 434 260001 440 260398
rect 390 259989 440 260001
rect 556 260398 606 260410
rect 556 260001 562 260398
rect 600 260001 606 260398
rect 556 259989 606 260001
rect 722 260398 772 260410
rect 722 260001 728 260398
rect 766 260001 772 260398
rect 722 259989 772 260001
rect 888 260398 938 260410
rect 888 260001 894 260398
rect 932 260001 938 260398
rect 888 259989 938 260001
rect 1054 260398 1104 260410
rect 1054 260001 1060 260398
rect 1098 260001 1104 260398
rect 1054 259989 1104 260001
rect 1220 260398 1270 260410
rect 1220 260001 1226 260398
rect 1264 260001 1270 260398
rect 1220 259989 1270 260001
rect 1386 260398 1436 260410
rect 1386 260001 1392 260398
rect 1430 260001 1436 260398
rect 1386 259989 1436 260001
rect 1552 260398 1602 260410
rect 1552 260001 1558 260398
rect 1596 260001 1602 260398
rect 1552 259989 1602 260001
rect 1718 260398 1768 260410
rect 1718 260001 1724 260398
rect 1762 260001 1768 260398
rect 1718 259989 1768 260001
rect 1884 260398 1934 260410
rect 1884 260001 1890 260398
rect 1928 260001 1934 260398
rect 1884 259989 1934 260001
rect 2050 260398 2100 260410
rect 2050 260001 2056 260398
rect 2094 260001 2100 260398
rect 2050 259989 2100 260001
rect 2216 260398 2266 260410
rect 2216 260001 2222 260398
rect 2260 260001 2266 260398
rect 2216 259989 2266 260001
rect 2382 260398 2432 260410
rect 2382 260001 2388 260398
rect 2426 260001 2432 260398
rect 2382 259989 2432 260001
rect 2548 260398 2598 260410
rect 2548 260001 2554 260398
rect 2592 260001 2598 260398
rect 2548 259989 2598 260001
rect 2714 260398 2764 260410
rect 2714 260001 2720 260398
rect 2758 260001 2764 260398
rect 2714 259989 2764 260001
rect 2880 260398 2930 260410
rect 2880 260001 2886 260398
rect 2924 260001 2930 260398
rect 2880 259989 2930 260001
rect 3046 260398 3096 260410
rect 3046 260001 3052 260398
rect 3090 260001 3096 260398
rect 3046 259989 3096 260001
rect 3212 260398 3262 260410
rect 3212 260001 3218 260398
rect 3256 260001 3262 260398
rect 3212 259989 3262 260001
rect 3378 260398 3428 260410
rect 3378 260001 3384 260398
rect 3422 260001 3428 260398
rect 3378 259989 3428 260001
rect 3544 260398 3594 260410
rect 3544 260001 3550 260398
rect 3588 260001 3594 260398
rect 3544 259989 3594 260001
rect 3710 260398 3760 260410
rect 3710 260001 3716 260398
rect 3754 260001 3760 260398
rect 3710 259989 3760 260001
rect 3876 260398 3926 260410
rect 3876 260001 3882 260398
rect 3920 260001 3926 260398
rect 3876 259989 3926 260001
rect 4042 260398 4092 260410
rect 4042 260001 4048 260398
rect 4086 260001 4092 260398
rect 4042 259989 4092 260001
rect -4092 -260001 -4042 -259989
rect -4092 -260398 -4086 -260001
rect -4048 -260398 -4042 -260001
rect -4092 -260410 -4042 -260398
rect -3926 -260001 -3876 -259989
rect -3926 -260398 -3920 -260001
rect -3882 -260398 -3876 -260001
rect -3926 -260410 -3876 -260398
rect -3760 -260001 -3710 -259989
rect -3760 -260398 -3754 -260001
rect -3716 -260398 -3710 -260001
rect -3760 -260410 -3710 -260398
rect -3594 -260001 -3544 -259989
rect -3594 -260398 -3588 -260001
rect -3550 -260398 -3544 -260001
rect -3594 -260410 -3544 -260398
rect -3428 -260001 -3378 -259989
rect -3428 -260398 -3422 -260001
rect -3384 -260398 -3378 -260001
rect -3428 -260410 -3378 -260398
rect -3262 -260001 -3212 -259989
rect -3262 -260398 -3256 -260001
rect -3218 -260398 -3212 -260001
rect -3262 -260410 -3212 -260398
rect -3096 -260001 -3046 -259989
rect -3096 -260398 -3090 -260001
rect -3052 -260398 -3046 -260001
rect -3096 -260410 -3046 -260398
rect -2930 -260001 -2880 -259989
rect -2930 -260398 -2924 -260001
rect -2886 -260398 -2880 -260001
rect -2930 -260410 -2880 -260398
rect -2764 -260001 -2714 -259989
rect -2764 -260398 -2758 -260001
rect -2720 -260398 -2714 -260001
rect -2764 -260410 -2714 -260398
rect -2598 -260001 -2548 -259989
rect -2598 -260398 -2592 -260001
rect -2554 -260398 -2548 -260001
rect -2598 -260410 -2548 -260398
rect -2432 -260001 -2382 -259989
rect -2432 -260398 -2426 -260001
rect -2388 -260398 -2382 -260001
rect -2432 -260410 -2382 -260398
rect -2266 -260001 -2216 -259989
rect -2266 -260398 -2260 -260001
rect -2222 -260398 -2216 -260001
rect -2266 -260410 -2216 -260398
rect -2100 -260001 -2050 -259989
rect -2100 -260398 -2094 -260001
rect -2056 -260398 -2050 -260001
rect -2100 -260410 -2050 -260398
rect -1934 -260001 -1884 -259989
rect -1934 -260398 -1928 -260001
rect -1890 -260398 -1884 -260001
rect -1934 -260410 -1884 -260398
rect -1768 -260001 -1718 -259989
rect -1768 -260398 -1762 -260001
rect -1724 -260398 -1718 -260001
rect -1768 -260410 -1718 -260398
rect -1602 -260001 -1552 -259989
rect -1602 -260398 -1596 -260001
rect -1558 -260398 -1552 -260001
rect -1602 -260410 -1552 -260398
rect -1436 -260001 -1386 -259989
rect -1436 -260398 -1430 -260001
rect -1392 -260398 -1386 -260001
rect -1436 -260410 -1386 -260398
rect -1270 -260001 -1220 -259989
rect -1270 -260398 -1264 -260001
rect -1226 -260398 -1220 -260001
rect -1270 -260410 -1220 -260398
rect -1104 -260001 -1054 -259989
rect -1104 -260398 -1098 -260001
rect -1060 -260398 -1054 -260001
rect -1104 -260410 -1054 -260398
rect -938 -260001 -888 -259989
rect -938 -260398 -932 -260001
rect -894 -260398 -888 -260001
rect -938 -260410 -888 -260398
rect -772 -260001 -722 -259989
rect -772 -260398 -766 -260001
rect -728 -260398 -722 -260001
rect -772 -260410 -722 -260398
rect -606 -260001 -556 -259989
rect -606 -260398 -600 -260001
rect -562 -260398 -556 -260001
rect -606 -260410 -556 -260398
rect -440 -260001 -390 -259989
rect -440 -260398 -434 -260001
rect -396 -260398 -390 -260001
rect -440 -260410 -390 -260398
rect -274 -260001 -224 -259989
rect -274 -260398 -268 -260001
rect -230 -260398 -224 -260001
rect -274 -260410 -224 -260398
rect -108 -260001 -58 -259989
rect -108 -260398 -102 -260001
rect -64 -260398 -58 -260001
rect -108 -260410 -58 -260398
rect 58 -260001 108 -259989
rect 58 -260398 64 -260001
rect 102 -260398 108 -260001
rect 58 -260410 108 -260398
rect 224 -260001 274 -259989
rect 224 -260398 230 -260001
rect 268 -260398 274 -260001
rect 224 -260410 274 -260398
rect 390 -260001 440 -259989
rect 390 -260398 396 -260001
rect 434 -260398 440 -260001
rect 390 -260410 440 -260398
rect 556 -260001 606 -259989
rect 556 -260398 562 -260001
rect 600 -260398 606 -260001
rect 556 -260410 606 -260398
rect 722 -260001 772 -259989
rect 722 -260398 728 -260001
rect 766 -260398 772 -260001
rect 722 -260410 772 -260398
rect 888 -260001 938 -259989
rect 888 -260398 894 -260001
rect 932 -260398 938 -260001
rect 888 -260410 938 -260398
rect 1054 -260001 1104 -259989
rect 1054 -260398 1060 -260001
rect 1098 -260398 1104 -260001
rect 1054 -260410 1104 -260398
rect 1220 -260001 1270 -259989
rect 1220 -260398 1226 -260001
rect 1264 -260398 1270 -260001
rect 1220 -260410 1270 -260398
rect 1386 -260001 1436 -259989
rect 1386 -260398 1392 -260001
rect 1430 -260398 1436 -260001
rect 1386 -260410 1436 -260398
rect 1552 -260001 1602 -259989
rect 1552 -260398 1558 -260001
rect 1596 -260398 1602 -260001
rect 1552 -260410 1602 -260398
rect 1718 -260001 1768 -259989
rect 1718 -260398 1724 -260001
rect 1762 -260398 1768 -260001
rect 1718 -260410 1768 -260398
rect 1884 -260001 1934 -259989
rect 1884 -260398 1890 -260001
rect 1928 -260398 1934 -260001
rect 1884 -260410 1934 -260398
rect 2050 -260001 2100 -259989
rect 2050 -260398 2056 -260001
rect 2094 -260398 2100 -260001
rect 2050 -260410 2100 -260398
rect 2216 -260001 2266 -259989
rect 2216 -260398 2222 -260001
rect 2260 -260398 2266 -260001
rect 2216 -260410 2266 -260398
rect 2382 -260001 2432 -259989
rect 2382 -260398 2388 -260001
rect 2426 -260398 2432 -260001
rect 2382 -260410 2432 -260398
rect 2548 -260001 2598 -259989
rect 2548 -260398 2554 -260001
rect 2592 -260398 2598 -260001
rect 2548 -260410 2598 -260398
rect 2714 -260001 2764 -259989
rect 2714 -260398 2720 -260001
rect 2758 -260398 2764 -260001
rect 2714 -260410 2764 -260398
rect 2880 -260001 2930 -259989
rect 2880 -260398 2886 -260001
rect 2924 -260398 2930 -260001
rect 2880 -260410 2930 -260398
rect 3046 -260001 3096 -259989
rect 3046 -260398 3052 -260001
rect 3090 -260398 3096 -260001
rect 3046 -260410 3096 -260398
rect 3212 -260001 3262 -259989
rect 3212 -260398 3218 -260001
rect 3256 -260398 3262 -260001
rect 3212 -260410 3262 -260398
rect 3378 -260001 3428 -259989
rect 3378 -260398 3384 -260001
rect 3422 -260398 3428 -260001
rect 3378 -260410 3428 -260398
rect 3544 -260001 3594 -259989
rect 3544 -260398 3550 -260001
rect 3588 -260398 3594 -260001
rect 3544 -260410 3594 -260398
rect 3710 -260001 3760 -259989
rect 3710 -260398 3716 -260001
rect 3754 -260398 3760 -260001
rect 3710 -260410 3760 -260398
rect 3876 -260001 3926 -259989
rect 3876 -260398 3882 -260001
rect 3920 -260398 3926 -260001
rect 3876 -260410 3926 -260398
rect 4042 -260001 4092 -259989
rect 4042 -260398 4048 -260001
rect 4086 -260398 4092 -260001
rect 4042 -260410 4092 -260398
<< properties >>
string FIXED_BBOX -4215 -260529 4215 260529
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 2600.0 m 1 nx 50 wmin 0.350 lmin 0.50 rho 2000 val 14.858meg dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
