magic
tech sky130A
magscale 1 2
timestamp 1712250795
<< nwell >>
rect -2519 -697 2519 697
<< mvpmos >>
rect -2261 -400 -1861 400
rect -1803 -400 -1403 400
rect -1345 -400 -945 400
rect -887 -400 -487 400
rect -429 -400 -29 400
rect 29 -400 429 400
rect 487 -400 887 400
rect 945 -400 1345 400
rect 1403 -400 1803 400
rect 1861 -400 2261 400
<< mvpdiff >>
rect -2319 388 -2261 400
rect -2319 -388 -2307 388
rect -2273 -388 -2261 388
rect -2319 -400 -2261 -388
rect -1861 388 -1803 400
rect -1861 -388 -1849 388
rect -1815 -388 -1803 388
rect -1861 -400 -1803 -388
rect -1403 388 -1345 400
rect -1403 -388 -1391 388
rect -1357 -388 -1345 388
rect -1403 -400 -1345 -388
rect -945 388 -887 400
rect -945 -388 -933 388
rect -899 -388 -887 388
rect -945 -400 -887 -388
rect -487 388 -429 400
rect -487 -388 -475 388
rect -441 -388 -429 388
rect -487 -400 -429 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 429 388 487 400
rect 429 -388 441 388
rect 475 -388 487 388
rect 429 -400 487 -388
rect 887 388 945 400
rect 887 -388 899 388
rect 933 -388 945 388
rect 887 -400 945 -388
rect 1345 388 1403 400
rect 1345 -388 1357 388
rect 1391 -388 1403 388
rect 1345 -400 1403 -388
rect 1803 388 1861 400
rect 1803 -388 1815 388
rect 1849 -388 1861 388
rect 1803 -400 1861 -388
rect 2261 388 2319 400
rect 2261 -388 2273 388
rect 2307 -388 2319 388
rect 2261 -400 2319 -388
<< mvpdiffc >>
rect -2307 -388 -2273 388
rect -1849 -388 -1815 388
rect -1391 -388 -1357 388
rect -933 -388 -899 388
rect -475 -388 -441 388
rect -17 -388 17 388
rect 441 -388 475 388
rect 899 -388 933 388
rect 1357 -388 1391 388
rect 1815 -388 1849 388
rect 2273 -388 2307 388
<< mvnsubdiff >>
rect -2453 619 2453 631
rect -2453 585 -2345 619
rect 2345 585 2453 619
rect -2453 573 2453 585
rect -2453 523 -2395 573
rect -2453 -523 -2441 523
rect -2407 -523 -2395 523
rect 2395 523 2453 573
rect -2453 -573 -2395 -523
rect 2395 -523 2407 523
rect 2441 -523 2453 523
rect 2395 -573 2453 -523
rect -2453 -585 2453 -573
rect -2453 -619 -2345 -585
rect 2345 -619 2453 -585
rect -2453 -631 2453 -619
<< mvnsubdiffcont >>
rect -2345 585 2345 619
rect -2441 -523 -2407 523
rect 2407 -523 2441 523
rect -2345 -619 2345 -585
<< poly >>
rect -2261 481 -1861 497
rect -2261 447 -2245 481
rect -1877 447 -1861 481
rect -2261 400 -1861 447
rect -1803 481 -1403 497
rect -1803 447 -1787 481
rect -1419 447 -1403 481
rect -1803 400 -1403 447
rect -1345 481 -945 497
rect -1345 447 -1329 481
rect -961 447 -945 481
rect -1345 400 -945 447
rect -887 481 -487 497
rect -887 447 -871 481
rect -503 447 -487 481
rect -887 400 -487 447
rect -429 481 -29 497
rect -429 447 -413 481
rect -45 447 -29 481
rect -429 400 -29 447
rect 29 481 429 497
rect 29 447 45 481
rect 413 447 429 481
rect 29 400 429 447
rect 487 481 887 497
rect 487 447 503 481
rect 871 447 887 481
rect 487 400 887 447
rect 945 481 1345 497
rect 945 447 961 481
rect 1329 447 1345 481
rect 945 400 1345 447
rect 1403 481 1803 497
rect 1403 447 1419 481
rect 1787 447 1803 481
rect 1403 400 1803 447
rect 1861 481 2261 497
rect 1861 447 1877 481
rect 2245 447 2261 481
rect 1861 400 2261 447
rect -2261 -447 -1861 -400
rect -2261 -481 -2245 -447
rect -1877 -481 -1861 -447
rect -2261 -497 -1861 -481
rect -1803 -447 -1403 -400
rect -1803 -481 -1787 -447
rect -1419 -481 -1403 -447
rect -1803 -497 -1403 -481
rect -1345 -447 -945 -400
rect -1345 -481 -1329 -447
rect -961 -481 -945 -447
rect -1345 -497 -945 -481
rect -887 -447 -487 -400
rect -887 -481 -871 -447
rect -503 -481 -487 -447
rect -887 -497 -487 -481
rect -429 -447 -29 -400
rect -429 -481 -413 -447
rect -45 -481 -29 -447
rect -429 -497 -29 -481
rect 29 -447 429 -400
rect 29 -481 45 -447
rect 413 -481 429 -447
rect 29 -497 429 -481
rect 487 -447 887 -400
rect 487 -481 503 -447
rect 871 -481 887 -447
rect 487 -497 887 -481
rect 945 -447 1345 -400
rect 945 -481 961 -447
rect 1329 -481 1345 -447
rect 945 -497 1345 -481
rect 1403 -447 1803 -400
rect 1403 -481 1419 -447
rect 1787 -481 1803 -447
rect 1403 -497 1803 -481
rect 1861 -447 2261 -400
rect 1861 -481 1877 -447
rect 2245 -481 2261 -447
rect 1861 -497 2261 -481
<< polycont >>
rect -2245 447 -1877 481
rect -1787 447 -1419 481
rect -1329 447 -961 481
rect -871 447 -503 481
rect -413 447 -45 481
rect 45 447 413 481
rect 503 447 871 481
rect 961 447 1329 481
rect 1419 447 1787 481
rect 1877 447 2245 481
rect -2245 -481 -1877 -447
rect -1787 -481 -1419 -447
rect -1329 -481 -961 -447
rect -871 -481 -503 -447
rect -413 -481 -45 -447
rect 45 -481 413 -447
rect 503 -481 871 -447
rect 961 -481 1329 -447
rect 1419 -481 1787 -447
rect 1877 -481 2245 -447
<< locali >>
rect -2441 585 -2345 619
rect 2345 585 2441 619
rect -2441 523 -2407 585
rect 2407 523 2441 585
rect -2261 447 -2245 481
rect -1877 447 -1861 481
rect -1803 447 -1787 481
rect -1419 447 -1403 481
rect -1345 447 -1329 481
rect -961 447 -945 481
rect -887 447 -871 481
rect -503 447 -487 481
rect -429 447 -413 481
rect -45 447 -29 481
rect 29 447 45 481
rect 413 447 429 481
rect 487 447 503 481
rect 871 447 887 481
rect 945 447 961 481
rect 1329 447 1345 481
rect 1403 447 1419 481
rect 1787 447 1803 481
rect 1861 447 1877 481
rect 2245 447 2261 481
rect -2307 388 -2273 404
rect -2307 -404 -2273 -388
rect -1849 388 -1815 404
rect -1849 -404 -1815 -388
rect -1391 388 -1357 404
rect -1391 -404 -1357 -388
rect -933 388 -899 404
rect -933 -404 -899 -388
rect -475 388 -441 404
rect -475 -404 -441 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 441 388 475 404
rect 441 -404 475 -388
rect 899 388 933 404
rect 899 -404 933 -388
rect 1357 388 1391 404
rect 1357 -404 1391 -388
rect 1815 388 1849 404
rect 1815 -404 1849 -388
rect 2273 388 2307 404
rect 2273 -404 2307 -388
rect -2261 -481 -2245 -447
rect -1877 -481 -1861 -447
rect -1803 -481 -1787 -447
rect -1419 -481 -1403 -447
rect -1345 -481 -1329 -447
rect -961 -481 -945 -447
rect -887 -481 -871 -447
rect -503 -481 -487 -447
rect -429 -481 -413 -447
rect -45 -481 -29 -447
rect 29 -481 45 -447
rect 413 -481 429 -447
rect 487 -481 503 -447
rect 871 -481 887 -447
rect 945 -481 961 -447
rect 1329 -481 1345 -447
rect 1403 -481 1419 -447
rect 1787 -481 1803 -447
rect 1861 -481 1877 -447
rect 2245 -481 2261 -447
rect -2441 -585 -2407 -523
rect 2407 -585 2441 -523
rect -2441 -619 -2345 -585
rect 2345 -619 2441 -585
<< viali >>
rect -2245 447 -1877 481
rect -1787 447 -1419 481
rect -1329 447 -961 481
rect -871 447 -503 481
rect -413 447 -45 481
rect 45 447 413 481
rect 503 447 871 481
rect 961 447 1329 481
rect 1419 447 1787 481
rect 1877 447 2245 481
rect -2307 -388 -2273 388
rect -1849 -388 -1815 388
rect -1391 -388 -1357 388
rect -933 -388 -899 388
rect -475 -388 -441 388
rect -17 -388 17 388
rect 441 -388 475 388
rect 899 -388 933 388
rect 1357 -388 1391 388
rect 1815 -388 1849 388
rect 2273 -388 2307 388
rect -2245 -481 -1877 -447
rect -1787 -481 -1419 -447
rect -1329 -481 -961 -447
rect -871 -481 -503 -447
rect -413 -481 -45 -447
rect 45 -481 413 -447
rect 503 -481 871 -447
rect 961 -481 1329 -447
rect 1419 -481 1787 -447
rect 1877 -481 2245 -447
<< metal1 >>
rect -2257 481 -1865 487
rect -2257 447 -2245 481
rect -1877 447 -1865 481
rect -2257 441 -1865 447
rect -1799 481 -1407 487
rect -1799 447 -1787 481
rect -1419 447 -1407 481
rect -1799 441 -1407 447
rect -1341 481 -949 487
rect -1341 447 -1329 481
rect -961 447 -949 481
rect -1341 441 -949 447
rect -883 481 -491 487
rect -883 447 -871 481
rect -503 447 -491 481
rect -883 441 -491 447
rect -425 481 -33 487
rect -425 447 -413 481
rect -45 447 -33 481
rect -425 441 -33 447
rect 33 481 425 487
rect 33 447 45 481
rect 413 447 425 481
rect 33 441 425 447
rect 491 481 883 487
rect 491 447 503 481
rect 871 447 883 481
rect 491 441 883 447
rect 949 481 1341 487
rect 949 447 961 481
rect 1329 447 1341 481
rect 949 441 1341 447
rect 1407 481 1799 487
rect 1407 447 1419 481
rect 1787 447 1799 481
rect 1407 441 1799 447
rect 1865 481 2257 487
rect 1865 447 1877 481
rect 2245 447 2257 481
rect 1865 441 2257 447
rect -2313 388 -2267 400
rect -2313 -388 -2307 388
rect -2273 -388 -2267 388
rect -2313 -400 -2267 -388
rect -1855 388 -1809 400
rect -1855 -388 -1849 388
rect -1815 -388 -1809 388
rect -1855 -400 -1809 -388
rect -1397 388 -1351 400
rect -1397 -388 -1391 388
rect -1357 -388 -1351 388
rect -1397 -400 -1351 -388
rect -939 388 -893 400
rect -939 -388 -933 388
rect -899 -388 -893 388
rect -939 -400 -893 -388
rect -481 388 -435 400
rect -481 -388 -475 388
rect -441 -388 -435 388
rect -481 -400 -435 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 435 388 481 400
rect 435 -388 441 388
rect 475 -388 481 388
rect 435 -400 481 -388
rect 893 388 939 400
rect 893 -388 899 388
rect 933 -388 939 388
rect 893 -400 939 -388
rect 1351 388 1397 400
rect 1351 -388 1357 388
rect 1391 -388 1397 388
rect 1351 -400 1397 -388
rect 1809 388 1855 400
rect 1809 -388 1815 388
rect 1849 -388 1855 388
rect 1809 -400 1855 -388
rect 2267 388 2313 400
rect 2267 -388 2273 388
rect 2307 -388 2313 388
rect 2267 -400 2313 -388
rect -2257 -447 -1865 -441
rect -2257 -481 -2245 -447
rect -1877 -481 -1865 -447
rect -2257 -487 -1865 -481
rect -1799 -447 -1407 -441
rect -1799 -481 -1787 -447
rect -1419 -481 -1407 -447
rect -1799 -487 -1407 -481
rect -1341 -447 -949 -441
rect -1341 -481 -1329 -447
rect -961 -481 -949 -447
rect -1341 -487 -949 -481
rect -883 -447 -491 -441
rect -883 -481 -871 -447
rect -503 -481 -491 -447
rect -883 -487 -491 -481
rect -425 -447 -33 -441
rect -425 -481 -413 -447
rect -45 -481 -33 -447
rect -425 -487 -33 -481
rect 33 -447 425 -441
rect 33 -481 45 -447
rect 413 -481 425 -447
rect 33 -487 425 -481
rect 491 -447 883 -441
rect 491 -481 503 -447
rect 871 -481 883 -447
rect 491 -487 883 -481
rect 949 -447 1341 -441
rect 949 -481 961 -447
rect 1329 -481 1341 -447
rect 949 -487 1341 -481
rect 1407 -447 1799 -441
rect 1407 -481 1419 -447
rect 1787 -481 1799 -447
rect 1407 -487 1799 -481
rect 1865 -447 2257 -441
rect 1865 -481 1877 -447
rect 2245 -481 2257 -447
rect 1865 -487 2257 -481
<< properties >>
string FIXED_BBOX -2424 -602 2424 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 2.0 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
