magic
tech sky130A
magscale 1 2
timestamp 1712071977
<< metal3 >>
rect -2686 13152 2686 13180
rect -2686 8128 2602 13152
rect 2666 8128 2686 13152
rect -2686 8100 2686 8128
rect -2686 7832 2686 7860
rect -2686 2808 2602 7832
rect 2666 2808 2686 7832
rect -2686 2780 2686 2808
rect -2686 2512 2686 2540
rect -2686 -2512 2602 2512
rect 2666 -2512 2686 2512
rect -2686 -2540 2686 -2512
rect -2686 -2808 2686 -2780
rect -2686 -7832 2602 -2808
rect 2666 -7832 2686 -2808
rect -2686 -7860 2686 -7832
rect -2686 -8128 2686 -8100
rect -2686 -13152 2602 -8128
rect 2666 -13152 2686 -8128
rect -2686 -13180 2686 -13152
<< via3 >>
rect 2602 8128 2666 13152
rect 2602 2808 2666 7832
rect 2602 -2512 2666 2512
rect 2602 -7832 2666 -2808
rect 2602 -13152 2666 -8128
<< mimcap >>
rect -2646 13100 2354 13140
rect -2646 8180 -2606 13100
rect 2314 8180 2354 13100
rect -2646 8140 2354 8180
rect -2646 7780 2354 7820
rect -2646 2860 -2606 7780
rect 2314 2860 2354 7780
rect -2646 2820 2354 2860
rect -2646 2460 2354 2500
rect -2646 -2460 -2606 2460
rect 2314 -2460 2354 2460
rect -2646 -2500 2354 -2460
rect -2646 -2860 2354 -2820
rect -2646 -7780 -2606 -2860
rect 2314 -7780 2354 -2860
rect -2646 -7820 2354 -7780
rect -2646 -8180 2354 -8140
rect -2646 -13100 -2606 -8180
rect 2314 -13100 2354 -8180
rect -2646 -13140 2354 -13100
<< mimcapcontact >>
rect -2606 8180 2314 13100
rect -2606 2860 2314 7780
rect -2606 -2460 2314 2460
rect -2606 -7780 2314 -2860
rect -2606 -13100 2314 -8180
<< metal4 >>
rect -198 13101 -94 13300
rect 2582 13152 2686 13300
rect -2607 13100 2315 13101
rect -2607 8180 -2606 13100
rect 2314 8180 2315 13100
rect -2607 8179 2315 8180
rect -198 7781 -94 8179
rect 2582 8128 2602 13152
rect 2666 8128 2686 13152
rect 2582 7832 2686 8128
rect -2607 7780 2315 7781
rect -2607 2860 -2606 7780
rect 2314 2860 2315 7780
rect -2607 2859 2315 2860
rect -198 2461 -94 2859
rect 2582 2808 2602 7832
rect 2666 2808 2686 7832
rect 2582 2512 2686 2808
rect -2607 2460 2315 2461
rect -2607 -2460 -2606 2460
rect 2314 -2460 2315 2460
rect -2607 -2461 2315 -2460
rect -198 -2859 -94 -2461
rect 2582 -2512 2602 2512
rect 2666 -2512 2686 2512
rect 2582 -2808 2686 -2512
rect -2607 -2860 2315 -2859
rect -2607 -7780 -2606 -2860
rect 2314 -7780 2315 -2860
rect -2607 -7781 2315 -7780
rect -198 -8179 -94 -7781
rect 2582 -7832 2602 -2808
rect 2666 -7832 2686 -2808
rect 2582 -8128 2686 -7832
rect -2607 -8180 2315 -8179
rect -2607 -13100 -2606 -8180
rect 2314 -13100 2315 -8180
rect -2607 -13101 2315 -13100
rect -198 -13300 -94 -13101
rect 2582 -13152 2602 -8128
rect 2666 -13152 2686 -8128
rect 2582 -13300 2686 -13152
<< properties >>
string FIXED_BBOX -2686 8100 2394 13180
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25.0 l 25.0 val 1.269k carea 2.00 cperi 0.19 nx 1 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
