magic
tech sky130A
magscale 1 2
timestamp 1713210209
<< metal3 >>
rect -1186 2440 890 4520
rect -400 2200 90 2440
rect -1186 120 890 2200
rect -400 -120 90 120
rect -1186 -2200 890 -120
rect -400 -2440 90 -2200
rect -1186 -4520 890 -2440
<< mimcap >>
rect -1146 4440 854 4480
rect -1146 2520 -1106 4440
rect 814 2520 854 4440
rect -1146 2480 854 2520
rect -1146 2120 854 2160
rect -1146 200 -1106 2120
rect 814 200 854 2120
rect -1146 160 854 200
rect -1146 -200 854 -160
rect -1146 -2120 -1106 -200
rect 814 -2120 854 -200
rect -1146 -2160 854 -2120
rect -1146 -2520 854 -2480
rect -1146 -4440 -1106 -2520
rect 814 -4440 854 -2520
rect -1146 -4480 854 -4440
<< mimcapcontact >>
rect -1106 2520 814 4440
rect -1106 200 814 2120
rect -1106 -2120 814 -200
rect -1106 -4440 814 -2520
<< metal4 >>
rect -198 4441 -94 4640
rect -1107 4440 815 4441
rect -1107 2520 -1106 4440
rect 814 2520 815 4440
rect -1107 2519 815 2520
rect -400 2121 90 2519
rect -1107 2120 815 2121
rect -1107 200 -1106 2120
rect 814 200 815 2120
rect -1107 199 815 200
rect -400 -199 90 199
rect -1107 -200 815 -199
rect -1107 -2120 -1106 -200
rect 814 -2120 815 -200
rect -1107 -2121 815 -2120
rect -400 -2519 90 -2121
rect -1107 -2520 815 -2519
rect -1107 -4440 -1106 -2520
rect 814 -4440 815 -2520
rect -1107 -4441 815 -4440
rect -198 -4640 -94 -4441
<< properties >>
string FIXED_BBOX -1186 2440 894 4520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
